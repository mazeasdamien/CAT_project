��   �c�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����DCSS_C�PC_T 4 �$COMMEN�T $EN�ABLE  �$MODJGRP�_NUMKL\�  $UFR�M\] _VTX �M �   $�Y�Z1K $Z�2�STOP_T�YPKDSBIO�IDXKENBL_CALMD��USE_PRED�IC? �ELAY�_TIMJSPEED_CTRLKOVR_LIM? *p D� �L�0�UT�OOi��O���&S. ǰ 8J\TC �u
!���\�� jY0 � � �CHG�_SIZ�$A�P!�E�DIS"�]$!�C_+{#�s%O#J�p 	]$J d#� �&s"�"{#�)�$��'�_SEEX�PAN#N�iG�STAT/ D�FP_BASE_ $0K$4�!� .6_V7>H�73hJ- � q}�\AXS\3UP�LW�7����a7r � < w?�?�?��?�?�x//	7ELEM/ T �&B.2�NO�G]@%CNHA��DF#� $DAT�A)he0  �PJ�@ 2� 
&P5 �� 1U*n   �_VSiSZbRj0jR(��VyT(�R%S{TR/OBOT�X�SAR�o�U�V$CUR�_��RjSETU~4"	 $d �P_MGN�INP_ASSe#�P B!� `CiH�77`e��.fXc1�CONF�IG_CHK`E_�PO* }dSHRS�T�gM^#/eOTH�ERRBT�j_G]�R�dTv �ku�dVALD_7h�e�4,��&T1r
0R HpLHt� 0  lt<8NerRFYhH~tD�5�1� ��W��_A$R��UPH/ (G%Q��Q�Q3?wBOX/ 8�@F!�F!�G �r��zTUI}Ri@  ,��F�pER%@2 {$�p l��_Sf�B�ZN>/ 0 IF1(@�p��Z_�0��_�0?wu0  @��QWyv	*��~����$$CL`  O���!���Q���Q�VERSIO�N�  �XK2�IRTU�AL�0�' 2 �?�Q  ((�����&@^���ʐ����ϟ��������d<�9�Cz  P�8���a��� ������ׯ���� �.�@�R�d�f����� �������Կ	��*� <�N�`�r����ϫϺ� ̿����߮�8�J� \�n�)ߒϧ߶��ς� �����%�4�F�X�~� |ߎߣ�.��������� �!�0�B�T�f�x�� ������������ />�P�b���v��� �������+: L^p����� �� /'/9/HZ l/�/��/��� �//#?5?D/V/h/z/ �/�?�/�?�/�/�?
? O1OCOR?d?v?�?�O �?�O�?�?O	_�O-_ ?_NO`OrO�O�O�O�_ �_�O�Oo_)o;o�_ \_n_�_�_Mo�_�o�_ �_�oo7IXojo |o�o�o�o�R�o�o �3�E�Tfx� ����Տ��ݏ� �A�S�b�t������� ��џ�����(�=� O�^�p���������ʟ ߯� ��$�9�K�]� l�~���6���Ưۿ� ���#�2�G�Y�h�z� ��������Կ����
� �.�C�U�g�vψϚ� �Ϯ��������<�-� �Q�c�r߄ߖߨߺ� ��������)�8�M� _�������q��� �������4�&[m |������������v 3BWix� ������ />?/e/w/��� ��/��///(/=? L/a?s?�/�/�/�/�/ �?�/O?$?9OH?]O oO�O�?�?�?ZO�O�? �OO O2OG_VOk_}_ �O�O�O�O�O�_�Oo _._CoR_goyo�o�_ �_�_�_�o�_	o*o `oQ@u��o�o�o �o�o�o��&8M� \q�������� ����"�4��X�J� �������ď������$DCSS_C?SC 25���Q  P�;���Z���~�A� ����w�د������ � �D�V��z�=���a� ¿��濩����߿@� �d�'ψ�KϬϾρ� �ϥ����*���N�� r߄�Gߨ�k��ߏ��� ���&���J��n�1� ��U��y������~�GRP 2�' ����	�s� ^��������������� '��7]H�l ������� 5 2kV�z� �����/
/// U/@/y/d/�/�/�/�/ �/�/	?�/-??*?c? N?�?r?�?�?�?�?�? �?OO'OMO8OqO\O �O�O�O�O�O�O_�O %__"_[_F__�_�_ n_�_�_�_�_o�_o�Eo0oio�_GST�AT 2�E�ߜ< 6�4���Z�a?�  5O+�ӿ�`�`S�d�Ҵ��aD/ ����D1	��X`<�e�a��e����dZ����o
s)���}uu9i�PqD1��d�`"ouW�a|q�`]Pb�8r�wuD 9ͺp�e�r�u�q�`��`���o�o �g��\�n��P��� ����Џ����o��� ��� �N�4�F�h��� |���̟��ԟ���� �J�ďz�������¯ ������
� �N�4�b� ,�j�P�b��������� �ο����8�f� h����گ�������� �&� �2�\��Dߒ� ��>����ߴ����"� ��F�X�2�|��h�z� ����������0�B� �.�x����߮���Z� ��������,>b tN������ �(4^8J ������v�/ $/�H/Z/4/f/�/j/ |/�/�/�/�/?�/? D??0?z?�?f?�?�? �?�?�?��?.O@O�? dOvOPObO�O�O�O�O �O�O_*___`_r_ L_�_�_�_�_�_�_�_ o&oOJo\o�_ho�o lo~o�o�o�o�o�o F 2|�h� ������0�B� 8oJ�x��d������� ���Џ�,���b� t�N������������� ̟�(��L�^�8�j� ��N�|�ʯܯv� �� ���H�Z�4�~���j� ��ƿ��������2� D��h�z�T�fϰ��� �����ϒ��.��� d�v�Pߚ߬߆߸��� �����*��N�`�:� l��p���������� ��� �J�\�6����� l������������� 4F R|Vh� �����0�� fx���� ���/,//P/b/ </N/�/�/�/�/�/�/ ??�/?L?^?T�? �?.?�?�?�?�? OO �?6OHO"OTO~OXOjO �O�O�O�O�O�O_2_ __h_z_p?�_�_J_ �_�_�_�_o.oo:o do>oPo�o�o�o�o�o �o�o�oN`: ��p���_�� ��8�J�$�6����� l���ȏ�����؏� 4�F� �j�|�V����� ���������0�ʟ <�f�@�R�������ү 䯾������P�b� <�����r���ο���� ����L��8ς� ��nϸ��Ϥ��� ��� ��6�H�"�l�~�Xߊ� �ߎߠ������� �2� �>�h�"�P���J� ���������.��R� d�>�����t������� ����<N(: �����f� ��8J$n�Z �������"/ 4//@/j/D/V/�/�/ ��/�/�/�/?0?
? T?f?@?r?�?v?�?�? �?�?OO�?&OPO*O <O�O�OrO�O�O�O�O _�/�O:_L_�Op_�_ \_n_�_�_�_�_ o�_ $o6oo"olo~oXo�o �o�o�o�o�o�o 2 (_Vht�x� ���
���(�R� ,�>�����t���Џ�� ܏����<�N�DV� ���p���̟���� ܟ�8��$�n���Z� ������¯�Ưد"��4��X�j�`��$D�CSS_JPC �2`�Q ( DQ�����ʴԿذ����ʿܿ 1� ��$�y�Hχ�l� �ϐ��ϴ�	�����,� Q� �2߇�V�h�z��� ���������;�
�_� .�@��d�v����� ����%���I��m�<� N��������������� ��3W&{J� n������� AO4�X�| ����/��O/ /0/B/�/f/�/�/�/ �/?�/'?�/?]?,? >?P?�?t?�?�?�?�? O�?5OOOXO}OLO ^O�O�O�O�O�O�O_ �OC__g_6_�_Z_l_ �_�_�_�_	o�_o4c*��S����Louo&o�o�`ddo�o�o�o �o	�o-�oQu <�`r���� ��;��_�&���J� ��n�ˏ��ُ���ڏ ����m�4���X��� |�ٟ����ğ!��E� ��0�y���f�ï�� 篮��ү/���S�� w�>���b��������� ����=��a�(υ� Lϩ�p��ϔ��ϸ��� ��%�K��o�6ߓ�Z� ��~��ߢ�����#��� 1��k�2�D�V�h��� ��������1���U� �y�@���d�v����� ������?c* �N�r���� ��q8� \����/�%/��FdMODEL ;2Skx�o(�
 <o$c (  o&�(�/�/ �/�/�/�/�/�/?? d?;?M?�?q?�?�?�? �?�?O�?ONO%O7O IO[OmOO�_�Oy/�O �O&_�O_\_3_E_W_ �_{_�_�_�_�_o�_ �_oXo/oAo�oeowo �o�o�o�o�o�o�O �O�O/��� ������P�'� 9�K�]�o���Ώ���� �ۏ����#�5��� Y�k���Se����� ������1�C���g� y�Ư������ӯ��� D��-�z�Q�c�u��� ������Ͽ�.�ɟ۟ 	�ψ��qσ��ϧ� �������<��%�7� ��[�mߺߑߣ����� ����8��!�n�E�W� ��?�Q�cϑ��y��� ��F��/�|�S�e�w� ������������0 +=Oa��� ������>�� �]o���� ����/#/p/G/ Y/�/}/�/�/�/�/�/ $?�/?Z?1?C?U?+ �?O}?�?�?�?�?2O 	OOhO?OQOcO�O�O �O�O�O�O_�O__ d_;_M_�_q_�_�_�_ �_�_�?*o�?�_oro Io[o�oo�o�o�o�o �o&�o\3EW i{������ ���/�A�o��;o i�{�菿�я���� �+�=�O���s���ҟ ����͟ߟ��P�'� 9���]�o��������� �����߯�^�5�G� ��k�}���ܿ��ſ� ���H��1�Cϐ�g� y��ϝϯ��������� D��-���'�U�g� ��O߽��������R� )�;��_�q���� �������<��%�7� I�[�m����������� ������J��3EW i{������ �/|Se� ������0// /f/A/S/�/;/ �/�/?�/�/>??'? t?K?]?o?�?�?�?�? �?�?(O�?O#OpOGO YO�O}O�O�Ow/�/�/ �O�O�O_1_~_U_g_ �_�_�_�_�_�_�_2o 	ooho?oQocouo�o �o�o�o�o�o �Ov_?Q'�� ���*���%�7� I�[������ޏ��Ǐ ُ����\�3�E����i�{���Җ�$DC�SS_PSTAT �����Q    ��� � A(&�K�2�o���� ������$�˟į֯���� ������'��SETUP ;	�Bȶ���X�r�������িۿ�g��T1SOC 2
K���鱃Cz�#�5�G� �CoP R�D$�Dl�Ϥ�^������ ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ������������,� >�P�b�t��������� ������(:L ^p����~�� ����-�Qc u������� //)/;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�__/_BS_ e_w_F_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1� _ U�g�y��_�������� ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{�J��߱�ğ ���������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ������/1/C/ /g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_�!o3o EoX/io{o�o\o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� ����ɟ۟����#� 5�G�ok�}��o^��� ů�������1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� �ߧ߹���������%�7�I�[�m�����$DCSS_TC�PMAP  ������Q_ @ ������������������	��
������������W�  �����������J����⡋���U��������U�� ��!��"��U#��$��%��&��U'��(��)��*��U+��,��-��.��U/��0��1��2��U3��4��5��6��U7��8��9��:��U;��<��=��>���?��@��UIROw 2�����������0B Tfx�����@��,1�� U��y����� ��	//-/?/Q/c/ u/�/�/�/6�/Z�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7O�/[O�/O�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_�NO�_��UIZN �2��	 ��� ��(o:oLoR�%ozo�o �oao�o�o�o�o
 .�oRdvE�� ������*�<� N�`�#�����e���̏ ޏ�����&�8��\� n���C�����ȟ��� ���ӟ4�F�X�'�|� ����c�u�֯请����0��_��UFRM; R������� w���������ѿ��� ��+�=�O�a�sυ� �ϩϻ���������`'�9�K�\�r��\� �ߖ�qߺ��ߧ���� ��&�8��\�n�I�� ������������� 4�F�]�o�|���-��� ����������0 TfA��w�� ���>Pg� t�%����� �/(//L/^/9/o/ �/�/�/�/�/�/ ?? �/6?H?_l?~??�? �?�?�?�?�?�? O2O OVOhOCO�O�OyO�O �O�O�O
_�O._@_W? d_v__�_�_�_�_�_ �_�_o*ooNo`o;o �o�oqo�o�o�o�o �o&8O_!n� �������"� �F�X�3�|���i��� ď�����Տ�0�B� Yf�x��������ҟ 䟿�����>�P�+� t���a�����ί��� �߯(�:�@�