��   v��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@���&�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	>4SUSRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  wXKaIRTs1�	o`'2 L1���L2�R�	 %,��?���b1`�c�c~a��a��� � � �d�o��
 ��a�o�o1CU �oz���� �c�
��.�@�R� �v���������Џ� q���*�<�N�`�� ��������̟ޟm�� �&�8�J�\�n����� ����ȯگ�{��"� 4�F�X�j����������Ŀֿ���`/TPTX������/�` sȄ��$/softpa�rt/genli�nk?help=�/md/tpmenu.dg���Ϩ� ���υ�����&�8� J���n߀ߒߤ߶��� W������"�4�F�X� ��|�����������a�`��oC ($p�-����T�?�x���a�a��c��H�c����l��k
��T�a���dh��at2�h�	f�����������`������h��_ep)��h#h�F�bc� Xc�B 1)hR_ \ _�� REG �VED]���w�holemod.�htm�	sing}l	doub �trip8?browsQ� ����u����//@/���d/ev.sl�/3� 1�,	t�/_�/ ;/i/??/?�/S?e?pw?�?�?�?� � �?�?OO%O7OIO[OmOO�E @�?�O�O �O�O�O_�F�	�?�? ;_M___q_�_�_�_�_ �_�_�_oo%o7oIo [omooM'�o�o�o�o �o�o+=Oa s������� ��?>�P�b�t����� ����Ώ���O��� ��L�^�_'_����� ��ş�����6�1� C�U�~�y�����Ư�� ӯ�o���-�?�Q� c�u���������Ͽ� ���)�;�M�_�-� �ϬϾ��������� *�<�7�`�r�A�Sߨ� ��q���i�����!� J�E�W�i����� ��������"��/��� O�I�w����������� ����+=Oa s������� ,>Pbt�� �߼���//�� ���^/Y/k/}/�/�/ �/�/�/�/�/?6?1? C?U?~?y?�?Y��?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__�R_d_v_�_ �_�_�_�_�_�_�o�*o�_o`oro�j�$�UI_TOPME?NU 1K`�a�R 
�d�a*Q)*de�fault5_]�*level0{ * [	 �o��0�o'rtp�io[23]�8?tpst[1[x)�w9�o	�=h5�8E01_l.p�ng��6mencu5�y�p�13�z���z	�4���q��]���������̏ޏ )Rr���+�=�O�a�~��prim=��page,1422,1h�����şן ����1�C�U�g����|�class,5p�����ɯۯ�����13��*�<��N�`�r���|�53�������ҿ�����|�8��1�C�U�g�y� ���ϯ���������"Y�`�a�o/��m!ηq0�Y�w�avtyl}T�fqmf[0nl�	>��c[164[w��59[x�qG���/��29��o�%�1���{ ��m��!�����0� B���f�x��������� O�����,>����2P����� \��'9K� �����������1��/$/6/H/Z/���|�ainedi'ߑ/�/�/�/�/���config=single&|�wintp���/$? 6?H?Z?	�ߐ??ٷ�gl[�<��?���08��
A���?,OH2��DO�?cO�O�z �6� �4s�x�O �O�$��Ol�E_W_i_ {_�_�_���_�_�_�_ oo/o�_Soeowo�o�o�o�$;�$dou�b5o��13��&odual�i38��C,4�o&�o9�o �n�o�a8���Ao ����&�8��\� n���������m��� ��
��.�@�K�d�v� ��������Z{?�;�M�sc�_;���s ��X�}���e�u��0� ���O_ �J�p�^�6e�u7������ ��Ͽ���P�)�;� M�_�qσ�ϧϹ��Ϡ�������"�1 �M�_�q߃ߕߠϹ� ���������7�I� [�m���������@�����!�����6(��]�o��������$��74������)�C��ߟT�	TPT�X[20�=Aw2A4#GJ���Bw1H ������8�"H����A#��[�tv�`�R��@2�K0F�11���5S:�$�treeview�3�f3��o}381,26M/_/q/0� �/�/�/�/�/�/~/? %?7?I?[?m?�o/܈5�o5%���?�?�?
? #O5OGOYOkO}O�?�? "2�?8"2K��O�O_�O��1�?�E�f_�x_�_ �6_ڀedit�a>_P_�_�_ oˉ/���_�Cooo �o�oB�o�o��oA �o�+=Oa s��o����� ��(�9���Q�x��� ������ҏO���� ,�>�P�ߏt������� ��Ο]�����(�:� L�^�ퟂ�������ʯ ܯk� ��$�6�H�Z� �l�������ƿؿ� y�� �2�D�V�h��� �Ϟϰ������ϕo�o ��o@ߧE�c�u߇� �߽߬�����O���� )�<�M�_�q���W� ��������&�8��� \�n���������E��� ����"4��Xj |����S�� 0B�fx� ���O��// ,/>/P/�t/�/�/�/ �/�/]/�/??(?:? L?��߂?1ߦ?�� �?�?�?�?O$O5OGO �?SO}O�O�O�O�O�O �O�O��2_D_V_h_z_ �_�_�/�_�_�_�_
o o�_@oRodovo�o�o )o�o�o�o�o* �oN`r���7 �����&��J� \�n���������E�ڏ ����"�4�ÏX�j� |�������a?s?蟗? �sO_/�A�S�e�w� ������������� �,�=�O�a�#_���� ��ο��=��(�:� L�^�pς�Ϧϸ��� ���� ߏ�$�6�H�Z� l�~�ߐߴ������� ����2�D�V�h�z� ������������
� ���@�R�d�v����� )���������ƚ�Ԕ*defau�lt%��*level8�ٯw����? tpsOt[1]�	�y��tpio[23���u���J�\menu7__l.png_|13��5�{�y4�u6���/ /'/9/K/]/���/�/ �/�/�/�/j/�/?#?�5?G?Y?k?�"pr�im=|page,74,1p?�?�?��?�?�?�"�6cl?ass,13�?*O@<ONO`OrOOB5xO@�O�O�O�O�O�#L �O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo]ooo��o`�$UI_U�SERVIEW �1֑֑R 
���o��o�o[m�o' 9K] ���� �l���#�5��o B�T�f������ŏ׏ 鏌���1�C�U�g� 
���������ӟ~��� ��v�?�Q�c�u��� *�����ϯ�󯖯� )�;�M�_�
��~��� ���ݿ���%�ȿ I�[�m�ϑ�4ϵ��� �����Ϩ�
��.ߠ� i�{ߍߟ߱�T����� ����/���S�e�w� ���Fߨ����>�� �+�=�O���s����� ����^�����' ����FX��|�� ����#5G Y�}����p ���h1/C/U/g/ y//�/�/�/�/�/�/ �/?-???Q?c?/p? �?�??�?�?�?OO �?;OMO_OqO�O&O�O �O�O�O�O�?�O_ _ �OD_m__�_�_�_X_ �_�_�_o!o�_EoWo io{o�o0h