��   ��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ������CCFR_�LTST_T � x$TP�_PROG �%$DATEJ �$TIMR2SU�F_NUM  w$TlSCHm��CHSoER�Rm  $APPL_TYPR ��ENS�� I�NI_POS� � �FRC�F;IN�MAX�	��DF�F� EMyPq V_LEN,GORI� I .I� �6DUM_R��UL� _FOR�CE_OK�MO�MENTsEND_AVE_F_���OSC_GDW��� _OFST ��/COM9�  $TOT�AL�5 2 o ��/AL� ? x AS ew������ �+=Oas@���1M!: � //&/8/J/\/n/�/ �/�/�/�/�/�/�/?�"?4?F?X?�D9� 8 $� �2 �1P 9(Q4IDX�2�1�X���$$C�LASS  ����FQ��'��'�;PVERSION�CX  {XKWQIRTU�`D_VP��dX'��%  ����_�_�_�_�� |�S��  o ��:oLoyopo�o�o�o�o�o�o���o �o 0Vh�om���_ �o���!o3o� ?�Q�~�u��������� ���? �2��V�h� ߏ�������� ���+�����d�[�m� ��������ǯ��7�� *�	�N�`�r��w��� ��̿�ݿ�׿#�5� Jϡ�S�l�wωϛϭ� ������A�"�4��X� j��ώ߁߲������ �����-�?ϙ�K�]� ������������ K�,�>��b�t���� �����������%� 7����pgy�� ��� C�6 Zl~������ ���/AV/� _/x/�/�/�/�/�/�/ 
?M.?@??d?v?�/ �?�?�?��?/�?O *O9/K/�?WOiO�O�O �O�O�O�O__W?8_ J_)_n_�_�O�_�_�? �_O�_�_o1OCO�_ �_|oso�o�o�o�o�o �oO_B!fx ����_�o� ��;oMob��k��� ������ŏ���Y :�L�+�p��������� ʟ��%����6�E� W���c�u�������د ϯ�� �c�D�V�5��z��������љ�$�CCFR_D �����'� ݟ �)��1�V�I�[��� �ϕ��Ϲ�������� .�@�g�d�v�Uߚ߬� #�����џ�=��)� ;�]�o����ߨ��� ������ ��8�{�H� n�M�������-����� ��G�!3g�y� ��������� B��fxW� �%���/Q +/=/b/q���/�/ �/�/�/?�/?:?L? �p?�?a?�?�?/?�? �?�OI/O5OGOi/ {/�?�?�O�O�O�O�O �O__D_�?T_z_Y_ �_�_�_9_�_�_Oo SO-o?o'osO�O�o�_ �o�o�o�o�o�o*! N�_r�c��1 ���o&�]o7�I� n�}o�o�����ڏя ����F�X��|� ��m���ğ;��۟	� �U��A�S�u����� �����ɯ������ #�P���`���e����� οE�ӿ��(�_�9� K�3������������ ������	�6�-�Zߝ� ~ߐ�oߴ���=����� ��2�i�C�U�z�� ���ߧ��������� �%�R�d��߈���y� ����G������*a� 'M_���	��� ���$/\ ��l�q���Q ��4/kE/W/?/ ���/	/�/�/�/�/ ??B?9?f?��?�? {?�?�?I?�?�?O)/ >Ou/OOaO�O�/�/O �O�O�O�O�O(__1_ ^_p_�?�_�_�_�_�_ S_ o�_!O6omO3oYo ko�O�Ooo�o�o�o 0;h�_x �}���]�� +o@�woQ�c�K��o�o ���Ǐ������!� N�E�r��������̟ ޟU����&�5�J��� [�m����������ѯ �����4�+�=�j�|� ��������ֿ�_�� ��-�B�y�?�e�wϙ� ��!���������� #�<�G�t߷��ߪ߉� ������i����7�L� ��]�o�W�ϵ���!� ������	��-�Z�Q� ~��ߢ���������a� 2A�V��gy ������
 @7Iv���� ����k//9 N/�K/q/�/��-/ #/�/�/�/&??/?H? S?�?��?�?�?�?�?��?u?O OB$( I/bO�/sO�O�O�/�/ !O�O�O___L_C_ U_�_�_�?�_�_�_�_  ow_$oo=/Zo�OWo }o�o�O�O9o/o�o�o 2);T_��_ �����
��� ,�Ood��ou���o��o �o�9����!�3� E�r�i������̟�� ��y�&��J�Y�n� �������ŏ׏1�� ��"��+�X�O�a��� ���Ŀֿ����σ� 0�#�Q�fϝ�cωϛ� ��ϯE�;�����>� 5�G�`�kߘ�ۿ���� ��������8�[� p�ρ��{������� E�����-�?�Q�~� u������������� ��2%Ve�z�� ������=�. %7d[m���� ���//�</// ]r/�o/�/�/�� Q/G/???J?A?S? l?w?�?��?�?�?�? O"O�?'ODOg/|O�/ �O�O�O�/�/�OQO_ _'_9_K_]_�_�_�_ �?�_�_�_oo�_>o 1oboqO�o�O�o�o�o �O�OIo�o:1C pgy���_�� ��$��H�;�io~� �o{������o�o]�S�  ��)�V�M�_�x��� ������ş
��.� ��3�P�s��������� ��ߏ��]��(�3� E�W�i���������޿ �Ͽ�&ϝ�J�=�n� }���ɯ�ϵ������ U���F�=�O�|�s� �߲����������� 0��T�G�uϊ��χ� �������i�_�,�#� 5�b�Y�k��������� ������(:��? \������� ��i4?Qc u���	���  /2/�V/I/z/��/ ��/�/�/�a/? %?R?I?[?�??�?�? �?/�?O�?*O<O�? `OSO�/�O�/�O�O�O �/�/uOkO8_/_A_n_ e_w_�_�_�_O�_�_ �_"o4oFo�_Koho�O �o�O�o�o�o�O	_ uo'@K]o�� ��o���,�>� �b�U����o���o�� ͏�m��1�^� U�g�������ʟܟ�  ���6�H���l�_� ����ُ��ůׯ��� ��w�D�;�M�z�q��� ����Կ��
��.� @�R�ɿW�tϗ���� ���Ϸ���*߁�3� L�W�i�{ߍߺ߱��� !�����8�J���n� a��϶��������� ��y�+�=�j�a�s� ����������+� ��BT��xk�� �������� PGY�}��� �#�/�:/L/^/ �c/�/��/��/�/ �/!6?�/??X?c? u?�?�?�?�?�?-/O  O�?DOVO�?zOmO�O �/�O�/�O�O
_?+? �O7_I_v_m__�_�_ �_�_�_7Oo*o	oNo `o�_�owo�O�o�O�o �o�o_#_�o�o\S e������/o �"��F�X�j��o� ���oď�oՏ�Ϗ -B���K�d�o����� ��ҟɟ��9��,�� P�b�ٟ��y�����ί �߯��%�7���C� U���y����������  �C�$�6��Z�l�� �σϱ����������� �/��ϛ�h�_�qߞ� �ߧ�������;��.� �R�d�v���{��� ���������'�9�N� ��W�p�{��������� ��E�&8\n ���������� �"1�C��Oa� ������/O 0/B/!/f/x/��/�/ ��/	�/�/?); �/�/t?k?}?�?�?�? �?�?OG/O:OO^O pO�O�?�O�O�/�O? �O�O�O3?E?Z_�Oc_ |_�_�_�_�_�_�_o QO2oDo#ohozo�_�o �o�o�O�o_�o	. =_O_�o[m��� �����[o<�N� -�r���������oޏ ۏ��5G���� ��w���������؟� �S� �F�%�j�|��� �����ӏ����� �?�Q�f���o����� ����ɿ����]�>� P�/�tφ����ϝ��� ݯ��)���:�I�[� ��g�yߦߝ߯����� ���$�g�H�Z�9�~� ���������!��� ��A�S������� ������������_� ,R1v��� ����+��K� ]�r�{���� �/�&/iJ/\/;/ �/�/	/�/�/�/��/ 5?!?F?Ug�/s? �?�?�?�?�?�?�?O 0Os/TOfOEO�O�OO�O�O�O  