��   K�A��*SYST�EM*��V9.4�0107 7/�23/2021 A 	  ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_���$$�CLASS  O�����D���DVERSIO�N  �XK/IRTU�AL-9LOO�R G��DD<x$?�������k,  1 <DwX< y�����Cu����	/��Z�Zm//�/�_/�/�/�/$ ��/�/	?';�$MNeU>A\"�  <�?/o?'_?�?�? �?�?�?�?�?OOO QO7OIOkO�OO�O�O �O�O_�O�O_M_�~;5NUM  ������92TOOLC?\ 
Y?[_�_ 3_�_o�_�_;o!o3o Uo�oio�o�o�o�o�o �o�o	7?mS e�����oZ�Q �Vy�Wy