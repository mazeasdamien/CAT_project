��   �A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG����DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !�� FT� @�� LOG_8	,C�MO>$DNL�D_FILTER��SUBDIRC�APC��8 .� 4� H{AD_DRTYP�H �NGTH�����z +LSq �D $ROBO�TIG �PEER��� MASK�M�RU~OMGDE�V��PINFO�.   $�$$TI ���RCM+T A$( /�QSIZ�!S� �TATUS_%$�MAILSERV~ $PLAN� �<$LIN<�$CLU��<${TO�P$CC�&sFR�&YJEC|!}Z%ENB � �ALAR:!B�TQP,�#,V8 S��_$VAR�)M��ON�&���&APPL�&PA� �%��''POR�Y#_�!�"�ALERT�&i2U�RL }Z3A�TTAC��0ER�R_THROU3UaS�9H!�8� CH- �c%�4MAX?WS�_|1��1MO	D��1I�  �1o �(�1PWD  Ɵ LA��0�ND��1TRYFDEL�A-C�0G'AERS�I��1Q'ROBIC�LK_HM 0Q'� X�ML+ 3SGFReMU3T� !OUU3f G_�-COP1�F33�AQ'C[2�%�B_AU�� 9 R�!�UPDb&PCO�U{!�CFO 3 
$V*W�@�c%ACC_HYQSN}A�UMMY1oW�2"$DM* �$DIS��SN,,	3 �	o!��"%"_WI�CT?Z_INDE�3�PgOFF� ~UR�Y�D�  �T�  �
 t Z!R%T�0N�(cD�)bHOUU#E%A/fVax>fVaMfLOCA� �#$NS0H_H-E���@I�/ w d�PARPH&��_IPF�W_�* O�F�PQFApsD90�VHO_� �5R42PS�a?�T;EL� P��r�90WORA5XQE� LVO#t�FS1�ICE��[p�$�c  O���zq��
���
op�PS�Axw  XK�qIz0ALw�q'0 V�x
���F������p�r�u�$� 2�{���r#� ��� �}��!�qi�����$� _FLT�R  �y�p *��������}��$�}2}��bSHA�R� 1�y Pe���t
�G�6�k� .���R���v������ �П1���U��y�<� ��`�r�ӯ������� ޯ?���u�8���\� ����ῤ�ڿ��;� ��_�"σ�FϏ�jϸ� �Ϡ����%���I�� m�0�Bߣ�f��ߊ��� �������E��i�,� ��P��t����������/���z _LUA1}��x!1.j�08���i�1z����255.��q���	��uh�2o��������������3����^  1C��4_��@� ������5����N�!3��6 O���u�������QJ�MA���MA�P��(�� Q�	 '��<a/�/�/{/��/�/�/�/?&?��P ?V?h?z?9?�?�?�?@�?�?�?
OO��?����ufOQL
ZD�T Status��?uO�O�O�O��}�iRConnec�t: irc�D/?/alert�N&_ 8_J_\_�G�O�_�_�_P�_�_�_���sP 2�q���_o1oCoUo goyo�o�o�o�o�o�o��o�s$$c962�b37a-1ac�0-eb2a-f�1c7-8c6e�b56401a8  (y_J�On�H�����ـP(!�X"�rZJ�p [D�r2cE\!)�,$e"� ـ[��M�4�q�X�~� ����ˏ�����%� �I�0�B��f���������w�W�8 D�M_=!W�G�S�NTP�	�%���-�������x�����4#��US?TOM 
�F���W  �3$T�CPIP���XHO%S"��ELO��W�T!�E�H!T�b���rj3/_tpdQO \��?!KCL��������v!CRT�Y�G���O"(�!OCONS�� ��ib_smon����