��  	vy�A��*SYST�EM*��V9.4�0107 7/�23/2021 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP�fBI�IZ@����ALRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� �� $ENABL�@C#� P dC#U5K�!MA�B �"�
� OG�f 0�CURR_D1P $�Q3LIN@S1I4$�C$AUSO4i O�D�"$SEV_A�ND_NOA�#PPINFOEQ/ �L �0?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� ���!PCOUPLE�,   $�!P=PV1CES0�24G�  C> �1�	 � $SO{FT�T_ID�2�TOTAL_EQ2� Q1}@NO�BU ?SPI_IN�0^��EX�3CREENu_�43BSIG@�3OEKw@PK_�FI0	$T�HKY�GPANE��D � DUMM�Y1dT�!#U4� Q�!RG1R�
 � $TIT1d ��� WTdWT� �WT7PWT5UV6UV7*UV8UV9UW0UW^W@QWUrW6QWU�W1�WU1�W1�W1�W2�R~�!SBN_CF�![�0$!J� �; 
2�1_CMNT��$FLAGS�]�CHE"$nb_OPTB� � �ELLSETUP�  `�0HO�@ PRZ1%�cM�ACRO�bREP	R�hD0D+�@��bl{�eHM MN�yB
1� UTOB �U�0 �9DEVICTST	I�0�� p@13�rpBqdf"VAL�#ISP_UNI��Cp_DO2v7iyFR_F�@K%D13�x[A�c�C_WA_t��a�zOFF_#@N.�DEL�xLF03q8�1�q%r?-q�pF�C?�>`�A�E�C#L�s�ATB�t�cW{�4c� $DB<0�"� S�("{&?��� \� VERq$F�!��d��_����dTMP1k_F��2��1_Rs���RrSAMO� �sE � [A��q�����REV�BI�L�!XI� �R�  � OD��`(�O2`M@��� �6�/�"�3�� A�l���@D�4d p E R�D_E �7�$F�SSB�&w`KBD�_S��VqAG� G
�2 "_��2ϑ� V�t:5?`��qC� �a�_EDu � �S C2��`S�p��4%$l �t$O�P�@qB�q7�_OqK���0, P_C� �7��d&�U �`LACI�!�a{�Ɛ� fqrX�M�  @$Dw�����@�p�_+R� BIGALLOW�G (KD2�2�@VAR�d!�AB ��BL{@S � ,�M�kp�h`S�pz@M�_O]8���C�F4d X�0GR�$@��M1�NFL�I�n�[@UIRE��84U�IT=$/0_�N�`S�"CFd0M�t� �#PEED��!ʹE`j��pS`JStVҒ`�\�3Np��`
ʗELBOF � �+ŷ+�p/0̲�3Pϲ� F�2f����1r�r@1J1E_y_T>!���`���g���G� �>A0WARNM�p�dp��E`ѳv`NST� �COR-$rFL{TR��TRAT �T�`� $ACC�%q�� �r��IX�.&��RT��S��� CHGV0I��.�Ti�pA�I9�T�!���� ��0�"`a���HDR�2��2�2J; �C�Ѫ��3��4��5��6*��7��8��9�!�`xD��@�2 @� TRQt�$Efl����C�N�_U��Y� �R�COC� <�� b�t���3Bq�L�LEC��MULTIV4�"��A
2>/�CHILD���c�� DET_Qb w 4� STY2�b�=��)2��8����C�  |A06$\����i`�d��C1TO���Ep�EXT���U��2��2G2�0��t�!/@AV�Qb.'������	� "�"	�/%�a�}����_sJ���# �W�[A��U�M�� N��" ��NP�$ L�0� �z�pA��$JOB ����b���IG�% d������-'p0|�����{�?q�s_M�r& t��3FL���BNG�A��BAi ���ߑ�/1�����0m��R0�P�Op�F��'��@:�$�bq��
2J�S_Rҳ�C,J�T(8,J��D/5CX)@�͑���@\�Q�P��(�`˻M?P~�ʂ��FACހ��SLEWL! % Y��!�:��R4d)�ː��ȓ�qG���@NHwANC��$LG����aRq��x���ī�A�p����aR�­�n4`6���o3P�m5RA�co3AZ�@�8찔����`FCT��S�_F����`�SM0�1I K�AE�0��0�Ұ D�����U��!����MP�B�a@Ж�H�KwAES�@NGT�1BWK�N�S �XYZW�`�2l���F}�Cg�C�*  ^0I\��B��}+.�STD_C�tt�A#�UST���U��,��PU�%V�IO�"�P�_up4�q��-|�$��SQOR�shR2p����`YOf0ʢSYېGP �q�Uupx�h`�ff����DBPXWOR�K��.�$SKcP_�paqO�DB0��TR�p / ����`��e��0+� D�q� _C�[bc,@gPLZc�a�t��"�"D��DgաcR "dE�С9ʨ� ���DB�1��0�RPQP�Rz�
 c�����1� �3�A�O�R�%L�i2�o[����� )3�o�dCF�4�o�����<�E�� 15�c�`RE���b6H $CE�o1$Lhs2$�c8���0y{INEҖ�Qs_D;A��ROS�� rֿ���q�s� �P�v�PAU�'�RETUsRN�rsBMMR��U���CR�pEWyMIP��SIGN��� ��LAL�(�@�3$P��4$�P�0+ 5<���PCW�+[�D#`ސ���t~qY�ҖGO_A�W� ��܀HP��rA�
�DCS"���C%Y�7�!�15ÁT3�̄2Ɗ2ԆNݐ�;��&KS��DEVI>�p 8 P� @�SRBѓճIԇP)�;�I_BYe�C�R�yTga�HNDG�b9 H��A.�۰��$DSBLR���Ն�P?��L��:0�P���FB✤�FE�q���Մ��v�
±;� '��A�ö�MCS<�А�TP����BH�0W��%�E����@�?��SLA�"�� <  p�IN�P�R������I�=/` ,��S0 P�6�J��x�FI0R�x��\%WQ�rWQW*�NTV�3r�V<��SKI�3TEL�v��j��ӄA�J�CjC_p��SA�F�¤�_SV�EOXCLU��}�� %D�PL��ϳY&������HI_V:@�BPPLY<`����}�����_ML+ }�$�VRFY_c��M�d�IOC��C_�&@��\���O7� �LQS�@}Bvd4\a��Ճk��PP�U�·�6S�AU��NF{F���Յ����+dQCHD`Q��D᮳`�AFSCP���T_�V�_B_VALi2 _�8͢'@ߑ ><p�PqTP��@|P �Ar͡N���� ?��j Tp��1 ���;��SGNԡ@�
$ ��"��q�@������ �R�دR��ANNUNp����Յ�$~P/�����&@
�&�ɢEF�PIqA @��F��.T�OT%�9�vd_�vd��؎�sa�PEM��NIB�bB���y'��A���DAYmSLOA�D8�kd��wc5b�EFF_AXIђ%C<paaCO���!���`_RTRQ�ԡD D��Yp� Q
�B(�E��1��� �C�@;?@�.� �A� �ԡEp���0�p�t�jDU%�j]��RCABԡFP�f2pNS��IDB�W�#l��1� V-�Vq_l�� � �DI�~�DG� 1$1��+T"�(!� w�0"
_��!E_����VE @SW�Y�! ��{�N�D���OH-���PPLY ��IRIQ�B�P ����q'��A ��C��0�0�-���N�F��@� RQDWf�MS�@AX�<G��LIFE`(�F}aRNY�b�W�� ��Cr@���NT�Y0PtAF3LAY4�OV;@n�HE��2SUPPIO�P|AR`_��Ց_XhC����Z�W�rA� Cጬ"�BXZ�0�a3Y2U(C�pT�P�p!QNG��JA ��_�0�B��10�DH{ `�CACH��)ѽ#SIZ��ٲ|-��@SUFFI��`đkd��wc�6sa��M�@�$I �8�KEYIMAG�sTM|q�3;1��66���Q9�OCVIIEc �aJ�B�0LK����?��@NP'@�$�K$�j�STw�!�2_��4\`�4��4|��0EMAIL����p5���FAULb�bL�B�s�SAX��9UP^2�DTWpԡ?M< $C=��Sl���IT��BU�F�'��'�<P2P�BBD=�C���BIS$@SAV�EOB8 @t"B�m �G�P�P�D=�Zpd��_B@sE-�F�HOT�r{���P:�0d`ZW�WAXmSC�bE�XB@���C_GY΢aYN_���N E<��D8�)`���UM���T��F�P�$�p��DI(��!E`WpX��aO���	GcA^�&�Ӕq�Q����G�F�� P (>pSV��r�kdw��p�ɡ�Q��aQ�0dp�Q
C�CC_�p�pAK�t:`��5d��R3184e�8�QDSPK6bPC{kIM�Crc�a	��Q UOg��u*��0IPL�c�� qdCTHs  �eb��T�q�rcHS�STcBSCY�� ��Vޠ"z p9SX(tn��NVԱGQs�(ts ofB@FY1�d0Tc�P7Q�qSC.��*cMER���aFBgCMP��`ET��� R)2FU�D�U6@��J"�CD hi�`P�3�PO��3!S$�� qgQ� u-�MS���z��-�������AK�T�� "��O2�T$CZO�P ����Ud�Ė�P=���CN�𢐚�����GROUȆ�����S� �MN ����������/�,����HR�b�{��0�PCYC���}����s�±��DE��_D�"��RO���Ԝ� #���|�i����d��� ��E�r��.��3M!�0&8�ALV K�U��Qj��P�pB���0�ER�TL �"V �,�P�.gQL0r1�U\P`Rg�����W��0$Ǥ��Ǥ��Pf�ɢC9�֥j�1���1ģP��XH *֡L��3y�� �v$���w�I�'�G����G���G���G�1G�7
D�8D�9D�YF�P�U1]�1j�1w�1��U1��1��1��1���2ƺ2P�]�2j�2�w�2��2��2��2���2��3ƺ3P�3T]�j�3w�3��3��U3��3��3��4ƲNAEXT��YlR �8qP��qP�u|P��U��AFDRZT"@VE��Q\��, r\RE��F\�2�OVMKc��A��T7ROV��DT�@�MX.�IN�ٚ�N��IND=�?�
i��PZPoPGBQ�(����bHD,�(�RIVx�p�2GEARKaKIO?K�҄�N�P���F�=�W0��2Z�_MCMM \�-F�UR�r[��ՠ�eA? ���?�;�X?;�E<��C�����OA�pR��\0P*Q �RI�5�OCETUP2_ ] w�FNCTD�` LET��S����^�OBBAC�fR^ T�0OB�T)��Z%�p+bl�=�I+FI{�l M0��p���PTe� �FL{UI�4_ �͑y7@UR�xA��Bp�Q pE@M�EMP���XR$wS+ ?x� J���@�CVRT|s��0x$SHOx9L>3�ASSp
Q8��`��BG_P������j��w����F�ORC B 4f�-`�2FU&�1�R)�2�R05s Aa �|y�NAVt���w ����S�2��$VISI���RSCTSEa�� Ps�5VӐO|�$w���,�w�$��I���@�FMR2��b ����� ���P���������樑����_����L�IMIT_���tC�_LM�����DGgCLFt��DY�(LDS��5����`��5c�B)� T�FS�@�d� P��2�SZP$GEX_158116P�np�q13W;5W6�9G<q��e �y��r�SWvEON9P%�E�BUG��1��GR��|`U�sBK��O�1� 1 PO@& �9�0�p�5�0M��YO%���SM��E�B���[���_E f� �p~� �TER�M'Eg0F�PORId�Q,@h0EaSM2�	O��,@i0E��h�oH�j0F_�UP� �k� -ZᎂQfw >C�@g�G�J� ELTOL���PWpFI?��Q&�13�|UD�Dh$UFR��$ʠ�AP�u] OT&WWpT���8SwNST��PAT�a=LTPTHJ�q�p�E���Sv��AART�~ �E� ~ FR�BREyL�Z��SHFT�b(�ATQ�X_� R�p�sJmF x@$�G�Pj}! �� �����PI�Pz$�U�r �pPAYLyO�`��DYN_8 �d�TQIޥ�`ERVO�am�Xs�4W����RP� ze�� RC�c�ޥASYMFL3TRޥ�AWJ�Gsтo�Es�~Q�im�qU��d��/a�U� nf�UP�[p9c[q�VOR��ML�P�GRA��l$@�2�6SPP���H���m �:R���OC�A�1���$OP��1�����Ѱ �RE�pR`�C��.�t�TSe] �RRU�u�x�Q��e$�PWR��,��R`R�_�swTy2��CUDps�i@lqR n���$H��!a�AD+DR��HAGVRz��o�h�A��R���o; H��SSC�P�����ç�j���w�SE�1�N�SCD_MN<p��p��8���pAaHOLL���p�p�Մ֣�CROH<�A\ND_C�ɢ�Na-�#pGROUP�[3`r_H�Y�0aq1 C���}�Q���P����р��j���w�����A����k2SAVEDȂ����� ���q3 $c��p_Dx��0���PZ�Y�H�TTP_ɠH��r; (ԠOBJ�h�6��$s�LEESO�|I�#�s � �הf ��_j�TC��S�`pcGKRL�HITCOU���1�L��p���s��p��pSSn���JQ�UERY_FLA�=��`_WEBSOC��HW���A�1�t��4�INCP	Uk2yOZ���.�3�s���r�˄r�� ��IOLN��u 8��R��@$SL�6r$INPUTM_A$�p��P�7 ��SL���1v���������c˵�b ��(�F_AuS2w��$L� o����Q�)��AP 0���0��!`HY��x��Q�,�UOP5x `=���s�M�h�M�o����pPc�p�����o�����y�?�I�P_ME�=y �X=�IPo�k2�_!NW�l2+�y1�r��7֞��SP��A�
F� BGk1�|M|a�=z lO0cTA47bv�AnpTI���e�� & �՞PPS��BU& ID0Ѣnp����p��M�p���FP{D���Ԗ�ɰN��& ��IRCA_�CN-� | �ڍ���CY��EA `�W�\��ct�r�;��b��qDAY_<����NTVAL�����rU�Ӹ�SCA�1`��CL�!�ѹ��ҏ=}���sR)�3�N_�pC5�����y�~�v�h����j�����,��� 2} o���=����j���LABpFQ��& ��UNI9��X@ITY��qьs�hAIR�@� 3�|��T R_URL[7�$A�EN�0��y:�=�T,�T_U>rABKY_�R�DIS��� ��iJY���$l�eJ	 Y�R�ō d �A�4�J��F�L@0I ��
��#
��UJR�� ���FH0�W� W�] f�J7a�tJ8!7u0��(7��	y8?APHI� �Q\D20J7�J8�buL_KE~��  �K���LM� � <��XR0�g�O�WA?TCH_VA�q<`<f�FIEL'�e�1yᰑ5� Y <Q1V)��`�CT �~1���LG��� $I�LG_SIZ���0>%�� =&4�=&FDH(I <(S(�1J&;()@U'G( : �sC#�&� �&4��&�j �&)@�&�a�5�@_0P_CM*S1G0:�1F�a 7:4: �t(9!�RE!_6R  _64�_6j k7I^8u8��0_6)@w7i8: RS�cP  Y3ZIPsDU��P�LNjFr���ӠDE%1�E��[*0�A`pL�CBDAU-EEA`8����tCB9@GH�r�l�@�BOO����� CW��IT0�wDs�S�REwЎHGSCRG0��X�D�|��o�MARGI�� T��LضKât�Bڤ@�	S{�?�W�D@�DK��JGM"WMNCHL;@�FN�%VKKW�9 IYUFWX�PWXF�WDWXHL�YSTPWZVWX��WX~@WX�RS�YHps[H�C�(t�S�bK���G"iU /�kT�G�3U `�^RG;YV�PObg�Z�E`�S2ATc�YYEXG�TUIIUI� N�S���!{��cS�cGP��@�^5��Fp�AN(��=�ANA@q��A�I@.���DCS��௃]s��]rOcxO"owSI�rzxS�x�HIGNS ��e#HQ �w�ftDEV gLLF�eA��yЈ���Ta2$I'��b��M��� �RAW�����m��V:�S1U�2U�3U�p4�b^pyЊ ���R�8tʵ�E˴���`�}`�F(��ST���RD@Y	�� �$E�C�.�����d%!� L T�f�� {�<�߃��[��.�8�u�i R�C_ � "�_ >��㼫@����MC�2�� �� CLDP|��TRQLI���יŔFLh��������D���E�LD8�����ORG��Q��8RESERV u�X���X���
���?� � 	��U�Ԕ��� PTא�	�<�����RCLMCȤX�j�ک�������MU /� ��$�DEBUGMASPiâ���2U�DTCp��E)+� �M�FRQ��� �� .)HRS_R%U��m�j�Ax�/e�FREQ%0�A$<P<'OVER��e#�2Џ��P`QEFI���%R�k�+����d���� \w ��(�$U��h�?L����PST�� 	��ACL@ɣ��%�ڣU �0�?( 	�1MwISC�� dA֕�RQ�	U�TB��@�� ���a��A�X��ǵ�EXC#ES.l�o�Mv��  ��X �n�SC�� � 	He��_���ȋ�!ۼ�����MK����@1�B_ F�LICM�B�@QU�IREcMO�OX����4�MLo�M� ���A��"m�Ȣ��NDA��e�!�B]/(�D*3[�INAUT�A[R#SM] %�pN��!�!c��S���PSTL�� 4�LOCf��RI��EX���ANG9r9���OD-Ah��|���� �MF"q%ʶ��n���`x����0/�SUP�t����FX� IG}G�A � ��� n��!Q�n�fn��� �@��P��_�@�c;��%�TI�N��r� M� �� t��+MD��IMA)��cp���ߡ��H����D#IAD�� W�A���;��a��DKC)b�O��� eМ ��C�US V ��9��Or�A_��� �� 0��������u ��P��P� P�KqEb�T3-$BF0zH�ND2ᢹ��2_TXw�XTR�Acs����LO�E@eО������2�N91�R�R2sŠ 1�))AA�� d$OCALI���%GQq�u2�� �Q�RINQ1y<$R�SW0���wABC��D_J� ��ѩ���_J3�
��1SP��) ��P��-3-SD���B@%J�P%y��!O�qyI�Y�CSKP暐$&0Js$J6X�Q�,�%�%�%�'��_A1Z��L!�!EL�qK"�OCMP��Y���@RTP�3+1�M ��1�/8p=:Z;4SMG�P���;JG��SCL����SPH_�pX��0�3� ���RTER$�y!pv_Pp�����A�@ڃX��4D�I�!n223U�"D�F��1LW�8VELבIN���`
@_BLcp9�D����DG0G(E� �N E�CH��TSA_<���IN�0��BeСN�E�B���A:A�__� ��E�B�5-��Dң�I�6���DH��g�D��$V�$�|3q$�Z0�����$�Q�RAeХH �$BEL� x��1�_ACCEA xPX�_PIRC_�0�h�K�NT��$PS��ʒL� ���Tߓ�@uW��RpvV �UY�WkS�W3�R_���_R�R�Pa��C�nUQ_MG��DDa�2��FW����[S;e�kSVR0hDEYkPP�ABN�WRO�0EEbV��oא�!V����VQ{A$USE_t�sP/�CTRt�Y{`1P�� G�YN�r�A� �fo ���aME�YHr`O@�QtINC3��Xb?d�¸8w���ENC�0L���9QVR�ďPIN�ʂI�Ru��l4NT|C)ENT23_�2��sLO�0���p��I�Љ��v�0��/��0�s�du.�C�@�vMOSI$aG�f a��X�PERCH  �s���2 ,���7�w��r �w�7 2�e�P`m#	A�R��L�dm#B�l'��u��zˆ�vTRK�5]�AY-����� �R
�����6!�Fr�MOM5���N�S ��Wcu��S�b_�DU��RS_BC?KLSH_C�R�� E�����c8ì�_r��| q�%CLALM�tpK�<��@�CHK� |���GLRTY{� �t��@���_�� �'_UM>�;�C>�-a�w1S���LMT _ALP�#l���w�Eq� ����p��U���X" D����Ӥp�PC=�p�Hp��#e;�CMC	\-`1gCN_�NL2�X#SFCQa�V�b���uw�1��Rv��CATB�SH��1d gv,�v�vv*�Q*00f `PAB�6r_PA�%�_� w0� ��!�$��JG������0�OG%��2TORQU�`%�s�g`p���1g`��_WT���91@ Q��S��S��I��I��ISF����W"X��f!)`VCUP0>�U��1#�!`7��!)ևJRK#�h�[�G D�Bu0MG M"�_sDLQ��GRV��`��S��S��H_08���P��COS��0��LNj��&��P �Z0���C�1�����1Z ����MY�������ۢ�THET=0�uNK23S��lS�CB��CBSC�AS�������S���SBS"���'GTS�!�aC!���37�C7X�@�$DU���}�E��(EeQl�_磿�NE�$�QK"�9�8�@��A������������LCPH����u��S&� >1�>@���O�hR
o���VVP'UV6
VCVQV_UVmV{V�	H@(.&��ECHQUH_HmH{H�	�O OO�%O�6
OCOQO_O*mO{Oo�F�����M)1�R$SPBA?LANCE_��}#�LE9�H_��SP��A"�"1�"@�PFULC�(�"�'�"@���J1�!1UTO_<��T1T29QR2N��\R�p14j15��� ��RLSP�T��O��0^Q��INSEG\R�qREVV6�p�qgDIF具I1��76�21��pOB�1ؑ���b�2s��p����L�CHWAR{bRA	B��d�bC�p��qdEV�X�P��'F���B0� 
(B��JQnwuROB �CR��XjE����CHQ_��T � x ?$WEIGHpր#$ �C'�Iq�psIF�a9`LAG�b�բS�b�0�bBIL��EOD>��p�BSTDbP�BP�1ؐ�@�/P(���A�@��@
[pHR<�a�  2��t�F/DEBU�CL�PR=|�MMY9�U�0qN޳kTր$D�Q�G�$UP"���  �DO_�PA�A� <�@%V0H���a��B�B�@N�sR�X_�p�`RO� �� %Z�T~p�qY�T�1MT�P�TICK�C�0T1"�P%c��&`N � 0�S �R���a�28e�2|De�PPROMPs�E�� $IR�i��a�b���bMA�I��@�r�e_�@��c�0�	pR��C�OD*SFU�`�FI�D_?��e0yb� G�_SUFF�� ��C�a�a3bDO`;gv0<e�@;fGR�C �2tYc$t�2/u�2;uP��t�T4P��@H�0�_FI)Q9�sO�RD�A �@]R3�6���r�a�P$Z�DT�e�AP�U��4 *�1L_NA��Q&`�r8eDEF_I�x�r^f�De�B7f�T7f0�De>�^fIS���j��Q��7dw�Dc��}�[T4;�͢RDP0����*SDf�O� >�RLOCKEޱs�8oJo\gy�rpUM u�rt0�t>�t�� $r�#u�$tN�$rV y�y�/s�0�/u�r/u@0�/s����x�PP�0 g��Ps����PW����6���pTE㑠T߫( �ALO�MB_�-�0�BV�IS��ITY�BA�"�O�CA_FRI3U��0SIs�W��!R#`~�.`~�3CS�B�WZ�Wf���\�l�_ɩ9qEAS�C9r3��T�ð���b�4|�5�|�6�CORMUL�A_Iޱ�TH]R�B��G�w��@���S\8cUCOEFF_O
am0��
aA��G���CS�@|RCA� �_�S$���C�Q�GR�� � �G $�D2�RX�PTM����b����SER�0T؄�t4P7�  �"LL:t��S��_SV��f�C���4P�u�U�4P� ��SETUs�MEA�`�`л@Q�r>�@� � ̰[@ eP>�������ǁD���r&`ǁ�Ą�����Dr�da�������ۢ��0�`R�EC�q��QSKy_� �� P�A?1_USER-1�2�l��0q�l�-1VEL@�l��0�҈��1I�p�0�MT�QCFG>bѰ  (`�0=OBNORE�@�P�����0��� 4� ��G�BAXYAZ�s1>0HS@���o_ERR�A� � 8��Q�`��/�0QX�����PBUFIN�DX��?*�MO�Rള H�@CU /��QA}�a�q�Ӑ2��q$J@���M�҄A>0��GⲴ � $SI9�0���`y1p�VO���t@OBJE� ��A�DJU�R����AYh�?E��D�OU�pp�}��a�r=|��T_0L���K��RDI�RP�X�0� x2g@D#YN��rB��T0���R\��P�@���OP�WORKbѵ,>�PSYSBU� чSOP��R�B���U����0P�PA`o���	B�OP-pU�1���1'RdQ8�/IMAGB��@D fRIM��^INɠ�/]RGOVRD����p�:P< \g@��0�����BL�B�,��0��PMC_E(�pR�YQN�M�dQ�]R1bR���S�L� cж � _$OVSL�6S�GDEX��L�2Be0��_� 6_p� 6@_p@UP]RuCX@��p�5�R� _ZE�R����$G�A:���bѷ �@�С1EO�`RI��B@
��`�!��Q��1��LbѸx�T<@
PATUS��sQGC_Tta�>#B�� H&1!�ĝ�cQ#�pcЇ� D�Q8 �<!L���0B<!�q]BѳX�EB �Ŗ"�"u$����@A UPԏ�m�CPX�`h&5[T3�^q"��PG�ջ��$SUB0!1E[��0!#JMPWAIqT� EH5LOW�<a�RCVF�a)`�BK1Ri���$CCC�R��b�7IGN�R_PL#DBTeB
PPq�ABW�`d�4��U�P�5IGzh`ICTNLN�6"�2R��肰�Nh`�PEED� 'HA�DOW
P�����E�&<D51�SPD.bѼ L�@AE �\@�jCUN�@;h@2�!R� �LY�p�0�:!T�PH_PK��ս��RETRI�E#��<��@�`FI�Ҿ ��p�@�D� 2���DBG�LV�3LOGSIYZ�㩁KTh1U^�2!TD'C�0_T����M9�CA�GP0]R�AS���CHECK��0�	�P��_A�26��It�LE�!��PAրT�B�"��PP�2_A� h $ARR�b� �s�K���O<p�7�ATT���2K�VGP�¥���S�CUX���P9L�`��� $���?SWITCHC2��-W��AS!RBCb�LLB_A�� /$BAI�D��чBAM�y�i!F�`J5�Ѷb6�f>ka_KNOW�S�b��U�AD�h��g@�Do��iPAYLOA����s_b�w��*wZsL[�A��<��LCL_�� !���Vr�a��ct�
qvF{yC:�Qz��Tt
i�IQxR<�QwN�mt�Bꠝ�J�q_Jt[q����ANDM��(��t[roq�աPL~z`AL_ �O`�g@��a�:�C�D:sE��J3�"��� T�PPDCK�� ���CO��_AgLPH2�x�BE��&�2�D�����1� � � �@D�_1z2DtD��A�R�!������TWIA4 �5 �6�MOM��,�L�9�L�4F���B_0AD,�p��9�p�F�PUB��R Q���9���F��!��"�|��`@�  �P9M>r� 2Ca�_��� e$PI�Aуx�w�~T9y�I!�I/�I=�@ݔ&n��!n�	1���n���u�� CHIG ^c C`5YD��YD`5�0 i��ƨ�1թ�1`5SAMP� ��)���p*�`5�`�s $� X���&��g�� q�Y@ 　�����)�o�d�h�H�0q�IN�� ����ۻ��`2���xش�!�GAMM��1SD!�ET��^�D����
$%�I�BR�!BI�$H�I�_yb����EĤ��A������LW ��������ֱƻ���t�0$�C�5CHK� �� g�I_ �����Ј���k��d��䎖j�"� {�$T� 1ĵ�}I RCH_D�1��0RNF'C��L�Eh���ػ����>@MSWFL�4̑wSCR�(100NPg�3(RL掷��,����`�Y@o�PI3A>�METHO����5��AX#� X8#@��BERI��)�%3U�R|@�u	͡���FF�*�n�
�}�����L��*�,�OO�Pn���B�}���AP	P�F� �PF�g�LR���RT��!�O��Y@՘�"�ޔ�1���ޔ~��=���R�A�PMGAsfS�V���P*PCU9R2�GRO&@�S_SA�a�$�#NO��C��"��$  t�Ϗ%7C��
�i���bq���DOXAA q�SQh�b꛵���Q����Q�"�Zs ��B`M��� � �p�YL��q�����S�r%�(Rt:����q�Ӏ�q_��C��є!M_WS �2���.�M�0�vp�!�m4;�CA:��"r�M��� ��A�l��!W4 �$��L"aGq4 ��2"��@2"��2"F��0��N�`Pv�Uc���X�@O����Z�%�j0��� ���M��ifx ���#����ѻP�:��_Ib� |e��( $ L�~69�~6F�$ %�`�7�6?�dan� sc�b2����@Hpb4P��Q�PMON_Q}U.� � 8�P�QCOU���PQT�HN HOm)@HY�S`ES�b)@UE�@�POGd�  ��@P ��ERUNW_TO�u`O��N��� PprEC��{Q INDE��R�OGRA�9`�2>2�NE_NO�DrE�IT��@V@INFO�A� Qa�J�A���OI�B�{ (��SLEQ��PQ��P�F V@SD���T� 4�PEN�AB`"p@PTIOyN�S�0ERVEv�pmW���AFRGCFNQ� @@J��zB+�z�R�Xn_�W|�pCQ_EDIT�A'� �A � Kϑ��5��E��NU�W�X�AUT@�UCOPAYϑ��l��L M���N#`'k<�PRUT�� *bN�POUCκ�$GwB�d���PRGADJn�A� he�X_�AI�ӷ �f� �fW�h�P�h�f���`��N^	�_CYC`"R/RGNSJU�b,��LGOIӔ�NYQ__FREQ��Wǰ���?qSIZ]TJ�L�A��6q�aG�ǰ��CcRE����J�IF/���CNA2�%}t_}G��STATUe0<��hGMAIL0�t�x�q��$DLAST�q�s�tELEMNQ�� �K XXFEASI[Q"]�V�I��r�� -(��⤰��I�@~��6r��,A�0��]�AB$DA��E�@ĠV�qu��BAS��v��µ�U8⠤�9 $����RMҐRW�����Ń`�#᠑��q�� 0 �r���m0	4� 2� 糝$մ ����� �����8E����DOU�C�Ԥa�tP����RG�RID�ADCBAR�S��TY\S푣�O\�0�A� cA_�t�!�`����O� KT�� � �@�0PO�R�C铚��SRV��p)	��DIB T_w�#�5���?���?�U4=�5=�6=�7=�I8!���FQ�NQ�a@?$VALU����Y1�@FJU��C !WUM!�Aӓ�q��ANǢ�q���Cr�TOTAL_X�t[�%�PW,sI��>:�REGEN8�M��3X���C,��1�@cTR���r8�_S ��M���V�a�T���Rv�E�s��.A�rB`n�V_H��DA3����S_YH�"Pv�S' AR02� }zbIG_SE%CȦ���u_v@ڴC_���$CM\�U%f�D�EW .�t�IL�Z�e�?�>TFT HAN�CA�m0
WW8�rSs��INT ��a��FlC�!MASK�㧀OVR��@��p+0�q�ѝ�OVCir�z�����SR��9�v�>���PSLG7�ա� \  QuI�""��pS��tx�UH�hG��γ��I�3U^0r�TE� ��� (u���JxQ�@`sIL_M_tb�Vc����0TQ@H���A��C�6�V=�CK�P_�9 U�M�l�V1k�V1y�2���2y�3��3y�4��4y�F�� +�����IN�VIAB E�2�9�25�U2A�35�3A�45�4A��@T�a2P� V���c���"��PLδpTOR@�IN����p�$�@�d��MC_F2@G �L	���Mb� I��%a� o0�2x��KEEP__HNADD!`$z�j	C�!������ЁOA_-`pŰ��ǁREM����q㒽��U��te�HPWD w `SBM��~ڐCOLLAB$�蠃���rPIT�p� 8bNO1FCsALW#�DON
s��$� ,�FL|] ��$SYN ��M�0CR����U_P_DLY�A��DELA��q�rY��0AD1$TA�BTP_R����QSKIP6%� 	���t@O� ��F��P_t@�B'�@�"�` ,'�Q:)�Q:)V�9*c� 9*p�9*}�9*��9*��z9*9�a�J2R�`*�@�SSX��T9s�! �A��!�`\�!�A\?i:�RDC����� ��PR�S��R�rq��,B���RGEp�PF���j�FLG	A�+��SWjY�SP9C�C�aUM_� ��_2TH2Nd��0��  1� ��� ��JR � �D�@��t9~�2_P�C�c�2S��ف@pL/10_C^rnп5�� �`��9��  N5�F�&�.A,4�`�Q)�=��1��eC�@�K�~��п5���0�� P�0DESIG\B9�VL1�91�6�C�G10� _DS`�Fἑ߰2`11Q� lQ ��ҍ XSDAT� �do�Bw*RIND���!Q2`��x!Q�R��HOMEKRW C�D2�B�_�_%_7_I_[_u�C3�B�~_�_�_�_�_�_W �D4�B��_@oo1oCoUo�W5�B��xo�o�o�o�o�o +�D6�B��o�+=Ogg7�B��r����� ��D8�B�����%�7�I� 0�@S|$�A�  Ѡ�Cb�p0�3� E��� T�0���IIO��!�I��G�O`_OP-�E��o1@��$��ASSp0����r�o0o0 �g��SI-�p��}�XK��I�RTUALo���A�AVM_WRK �2 ��� 0  �5�y����� �	7�(�K�o0B���9�v�]�{�'� ����6���������sBS�P1 1��� <ϯ @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ��������������0�B�T��C�AXkLM_�W��$�7  di�INr���h�PRE�0E������_UP<B��������IOCNV_��0�� Ȁ�P��U�S�� �
�IO�Vw 1̛P $����a�L��I��?� W�w�l~���� ��� 2DV hz������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯ԯ毀��
��.�@�R�i�L�ARMRECOV� ��{��%L�MDG 5�@ Z�LM_IF 5��W����#� 5�C��f�xϊϜϭ�?, 
 ���πQ�]��� �2�C�$ ��g�Nߋ�Jϯ����������¿NGTOL�  �� 	 �A   5�G�i�P�PINFO �� ��z����{�  �²�� ��	���-��)�c�M� ��q����������� ��1CUgy�����ǺPPL�ICATION �?$�����Hand�lingTool�  
V9.?40P/17F��
88340�$F0J7549�$+7DF�5�None��FRA� �6g�_ACoTIVE_�  ��.�  �UTOMOD���,���CHGAPONL�/ /#OUPL�ED 1ܹ� �l p/�/�/�CU�REQ 1	ܻ � T�)�,�,	��/ 5� 4����"��$�H�%o"�*HTTHKY?���/�/�/ ?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�׏����ŏ�� ����1�C�U�g�y� ӟ������ߟ���	� �-�?�Q�c�u�ϯ�� ����ۯ����)� ;�M�_�q�˿������ ׿ݿ���%�7�I� [�m��ϑϣϵ����ό<�%TO��#DO_CLEAN</|�s�NM  $� �/���������	�.DSPDRY�Rz��HI ��@ ��u�������������)�;�M��MAX� Z��1K'k��XZ�jg"j�PL�UGGZ [�g#%P�RC,�B�����d�V���O��5�G�SEGF3 K#. �߭�u������(LAPR�e'3 #5GYk}������.#TOT�AL����.#USE+NUR _+ @�D/�2� RGDISPWMMC1 ��C9&}�@@G�_$OP�r��=[#_STRI�NG 1
++
��M$ S��
�!_ITEM1�&  n��/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O�<OI/O S�IGNAL�%�Tryout M�ode�%Inp�|@Simulat{ed�!Out�LOVERRO� = 100�"In cycl�E��!Prog A�bor�C�!xDS�tatus�#	H�eartbeat��'MH FauylWSAlerY OO=_O_a_s_�_�_�_8�_�_�_ V��+ V��/�_0oBoTofoxo �o�o�o�o�o�o�o�,>Pbt�_WOR1 �+�q o�� ��
��.�@�R�d� v���������Џ��8��*�PO�+ Q P��{9�s��������� ͟ߟ���'�9�K� ]�o���������ɯK�DEVS���g��� -�?�Q�c�u������� ��Ͽ����)�;��M�_�q�PALT m���r��������� ��,�>�P�b�t߆� �ߪ߼���������GRIp��+<��� d�v��������� ����*�<�N�`�r� ������*�" Rm�� T��,>Pb t��������(:L��PREG�΅��^�� ���//*/</N/ `/r/�/�/�/�/�/�/��/RM�$ARG_��pD ?	����31� � 	$RF	+[G8]G7�RGh9�&0SBN_CONGFIGa@3;�A�B��1�1CII_S?AVE  RD�1��3&0TCELLSETUP 3:�%  OME_I�ORMRL%MOV�_H�0 OOREP���QO:UTOBA�CK�139�2�FRA:\r �\Or�0'`�@�r�H� �K�0� 25/1�2/01 20:_21:02ri8�r_$_Q_H_�L�� q_�_�_�_�_�_�_r��_ o2oDoVohozo o�o�o�o�o�o�o
 �o.@Rdv� ���������ׁ  �A_tC_\�ATBCKCTL.TM?�W�i�{���\��fKINI���E��5�1q@MESSA�G�0Ɓ�1;0ыODGE_D�0�6�5���O���nCPAUS�d� !�3; ,,		�i035h� v�\������������ ڟ����J�4�n�X��j�����;�E�TSK  K��O��q@�UPDT��ćd���XWZD_E�NBĄ�:�STA�Å31�%1WSM_�CFG 35��57b�GRP �2l� F2B��  A�9XIS~�0UNT 235:�1�0� 	ۯ�� M1�"��F�1�j�U����yϞ���ǴMET&��2ֹ��P���x��,߿�SCRDf�+1l��@��5�2!߅ߗߩ߻������OrQ�9r�/�A�S� e�w���߭������ ����+�����7tA�GRϰ	�)�j�:�N5A@2;	tDg��_ED1l�
� �%-@�ED�T-X�.J����L�4@-tC��r�i2g_F���  ��t2}-K[� .�&�Xj �v3I����r@�$6�Zv4/ �b/��>/�/�/�/&/v5�/Q/.?u/ �
?u?�/�/d?�/v6�??�?A?��?AO �?�?0O�?v7yO�? �OO��O_TOfO�O��Ov8E_���_P �n_�_ _2_�_V_v!9o�_^o�_S�:o��o�_�_�o"ovCR |�O);�Mo�o��o^�oj��NO_�DELv�h�GE_�UNUSEt�f�I�GALLOW 1���   (�*SYSTEM�*�	$SER�V���)�E�REG�2�$T��)�NU�MW�|�j�PMU|�p�LAY����PMPA�LJ���CYC10Ķ~Ɏ�����UL�SU��k�˂à3��L�>�BOXOR=I[�CUR_+�j��PMCNV���+�10ߎ��T4�DLI)�$�F�	*�PROGRA1�?PG_MI���F�AL�� ����B�)�$FLU?I_RESUχW�a�{���MR@�O��|�0�ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9� K�]�oρϓϥϷ���������rLAL_OUT �S��WD_ABORЀ��K�ITR_RT/N  rd���N�?NONSTO��y�� �CE_RIgA_I�py��������FCFG �����rn��_L�IM@�2�� �  N 	P�D1�}b<L�N����`�  ����rha
p���\���PA8��GP 1�����o�8�J�\��CO  C2���>��aH��������Cf��Uz��������x����\�������CU������m�rg?���HE�p�ONFI��X�.G�_Pq�1� �u�x��������.KPAU�SH�1���  ߂�>�,jPz �������
/ 0//T/f/L/�/ P��A�y�ի�Mn�NFoO 1	��� ���/}b�/%?�~b D��}bD��4  � 7?I;��O����rgJ��COLLECT_���	�B��ך7EN���y�`Ҷ2s1NDE��3 	���r�1234567890
G}bC���OF����~a)UOzOC| TOfO�OD{�O�O_�O �O�OK__(_:_�_^_ p_�_�_�_�_�_#o�_  ooko6oHoZo�o~o@�o�o�o�o�6�!�;� �=�2IO ##�9�1,7x�}����KwTR �2%$/}(��fy
�o�~�9 %Z}�z>Dy_WMOR�&� �� $t�1t���z������ԏM����'[�,�>?'']0)���KT1���*P��(/}�����>��_�=L����R���)}?������K1A�j,:Ⱦ�x��A]02��Bː��B����@������:�d�<� <#�
�1�$�����I�3*��@�N�+�[�k��d��T_D�EFPROG ����%���~�SpN�USE��/��KEY_TBL  �����"�	
��� !"#$%�&'()*+,-�./G:;<=>�?@ABC��GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~��������������������������������������������������������������������������������͓���������������������������������耇����������������������q��LCKpϬ�م�ϠSTAU�z~�X�1_ALM6��]��_AUTO_�DO����j�IN�D�48Ι1R_T1t�f�T2�ϧՔӚ���TRL��LET�Ew���_SCR�EEN �_kcsc��U���MMENU 1,~�  <�� ����,5gߑ���~#�� �������8��!�n� E�W�}�������� ��"����1�j�A�S� ��w����������� ��T+=�as ������> 'M�]o�� ����/://#/ p/G/Y/�/}/�/�/�/ �/�/$?�/?Z?1?C? i?�?y?�?�?�?�?O �?�?OVO-O?O�O|�J�_MANUAL�Ϫ�DB�����DBG_ERRL捠-V�pq ЕO!_3_E^�ANU�MJ��~���?�D�BPXWORK 1.V�_�_�_�_��_�_�DBTB_�� /�M��;qꚔqDR�WAYz�CpqGCP ��C=�>�AdS��J_�B�Y��Փ��H_�@ +10�{�
�_�o�5��o�of_M��I�S5�Nk@*�sON�TIM����ɼ5v�i
ޥ�cMO�TNENDӯ�dR�ECORD 26�V� ���G�O��q���Nb�	� �-��x5�\����� ����ȏ_�u���m�"� ��F�X�j�|����� ğ3��������B� ��f�՟��������/� �S��w�,�>�P�b� ѯ�������ο�� �s�(ϗ�!ϻ�pς� �Ϧ���ϵ��� �o� p�8�J߹�n�Y�g���o�MEN������@]�����H�o��E u�����,���P� ��)�;���_��������������L�wTOLERENCLdsBȕbZ`L���@�CSS_CNST_CY 27�Y��@	���b�M[m ������� %3EWm{���(DEVICE 288'f�// (/:/L/^/p/�/�/�/ �/�/�/�/ ??$?6?�H?Z?l?~?�?w+HNDGD 98�,`Cz�:�q+LSw 2:8 �? OO,O>OPObOtO�?�*PARAM �;�i|bpe�D�5�5SLAVE <�=��7_CFG =��O�CdMC:�\* L%04d.'CSV�OePc-_�b6��A ZSCHbP�1A�o�Nm_�_�G��F�R�Q�_�_�_�H�`�JP�c�^�a��$m�DRC_OUT >�=7a�O�_NOCOD�@?��g�MSGN �@�u�r�01�-DEC-25 20:22]P�o�c�� [�����i�a�N�`���s��M��Þ��,�\�EVE�RSION ��jV4.5.�2��EFLOGI�C 1A� 	h��ya�}sr�PROG_ENB�  �U�6�sULGSE E d�Esr_ACCLIM�v���C� �W?RSTJNT�w�a�csqMO�|�Q�BA�INIT B��e� ?�OPT��@ ?	~�W�
 	R575�CV��74��6��7��50Ո1Ոft�y��|mw��TO  ���	T�nvVe�DEX��wd�b�l�PA�TH v�bA�\Z���˟��HCP�_CLNTID y?Qv�C !k����IAG_G�RP 2G�I ��� 	 �E7� E?h �D�� C� �C ��B���@!�U���!�}�� �����C��C�m�B�N�Bz�oOB�)�B�k�!�f38�3 678901�2345��P�T���  A���A���A��A�O�A���A{+As��Aj�RAbJ�AY%!��3a@ŠZTpZPY� A�  ]PB4!���0!���3a
��������Q�A����A���A����A�����hA�x~�Ao�7A�f9X~�Q�>��mX�j�~���z�����_�AY�;�AS�TAM�^�AGdZA@��A:bA3%�A+�-A$J�z�Q���ϖ�@��;d�ƀ��@{��@u�-@o��@i�7@c�C�@\�j@Vs{`�n��5?t���Ϝ�"�@_��@�Z^5@T��@�O�@IG�@�C33@<��@�6�+@/N�(�`\�n�ߒ�0߶�s��nE�@h��@b�!@\��V�ff@P��Ihs�@B��@;� t߆ߘߪ߼ߞ�H�p� ��`���B���� � ���6������~��� n�����P�����U�,����E���]���p�>8�Q�0��R?��  <p�7�Ŭ�X'Ŭ5AF<dp�@�p���У@�� � }@m�A�hZP�U�=+�<��
=T���=�O�=���=�<���<�� ���^ ��?� �C�  �<(�U�R 4r|�V�)���4!�A@2b?x���j ��x��|�!�����/�@/R/��?�#�
t"�\>x� �%p���G��/G�p�8`�! �]T\Q�p�8���!���$����CnB�L�o�q��A?/<�M'�uv?�4�?�v�D�  D� � CΟ?0<�?�? <`�?O-O�V��?ZO�?~O1;�H �HE��OgO�O�O__ 	_B_-_f_Q_7�`/Z_��_0�CT_CON?FIG H�o/c�eg�u2�STBF_TTS�w�
�ycHp�U�f�}`MAU'���RM_SW_CF�PI?��  q�8zOCVI�EW/`[�we{���	O�o�o�o�o	 ��oDVhz�� -����
��� @�R�d�v�������;� Џ����*���N� `�r�������7�̟ޟ ���&�8�ǟ\�n� ��������E�گ�����"�4��\RChcK��<b!ЯB�l������ſ���ؿ�!dSB�L_FAULT �L_��h'�GPM�SKg:��PTDI�AG M�Y{a�D3�!aUD�1: 6789012345���R���WB�P�_������	� �-�?�Q�c�u߇ߙ� �߽�������R6��B��M
��;��VTRECPpς�
�Ă�� C��Ͼ��������� *�<�N�`�r������� ��������)�&�g�UMP_OPTIcON`3�@TRhbtc7�aPMEe�TY_TEMP � È�3B��"`� �A� �UN�IM`e�\fYN_?BRK N�o�f?EDITORFL�_X�ENT �1O_�  ,&��V/D��Up �����/�+/ /O/a/H/�/l/�/�/ �/�/�/?�/�/9? ? ]?D?l?�?z?�?�?�? �?�?O�?5OGO.OkO�RO�OvOMGDI_STA��Q���NC_INFO �1Pok�����P`�OW�C�B1Qok ���I_<_/
/d�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o n4FXjxy �Qx������ 
��.�@�R�d�v��� ������Џ����z -7�I�[�m������ ��ǟٟ����!�3� E�W�i�{�������ï կ����%�/�A�S� e����������ѿ� ����+�=�O�a�s� �ϗϩϻ�������� ��9�K�]�w�mߓ� �߷����������#� 5�G�Y�k�}���� ���������'�1�C� U���ߋ��������� ����	-?Qc u������� ��);M_y�� ������// %/7/I/[/m//�/�/ �/�/�/�/�/!?3? E?W?q{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �O?_+_=_O_i?[_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�o�o�o�o_�o# 5Ga_s_}��� ������1�C� U�g�y���������ӏ ��o�-�?�Q�k u���������ϟ�� ��)�;�M�_�q��� ������˯ݯW�	�� %�7�I�c�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� �������/�A�[� e�w߉ߛ߭߿����� ����+�=�O�a�s� ������������� �'�9�S�I�o����� ������������# 5GYk}��� �����1� ]�gy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�� ??)?;?U_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�/�O_!_3_ M?W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�O �o+E_7as �������� �'�9�K�]�o����� ����ɏ�oՏ���#� =OY�k�}������� şן�����1�C� U�g�y���������ۏ ���	��-�G�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ�3������ %�?�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������7�A�S� e�w������������� ��+=Oas �������� /�%K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ ���/�/?�/9C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�/�/�O�O __1?;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�O�o�o�o)_3 EWi{���� �����/�A�S� e�w��������oя� ���!�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ������ۯ����+� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϷ�ɯ�� ����	�#�-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������� %�7�I�[�m������ ����������!3 EWi{����� ����/AS ew������ �//+/=/O/a/s/ �/�/��/�/�/�/ ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O�5OGOYOkO}O�O�/ ��$ENETMO�DE 1R5�  � �� �%�O�K�@O�ATCFG S^5�AT��BC�UDATAW 1T�I!P��A*W_*�Hu_�_��_�_�[d�_�[1 �&�_	oo-o?oQoco uo�_o�o�o�o�o�o o,�oM_q� ��!3���� %�7�I�������� ��ǏُS� �w�!�3� E�W�i�{������ß�՟������@RP�OST_LOPV@[��
%V_�q�������ARROR_PR;�%�J%��ׯ���TABLE  ��K?�,�>�'�R�SEV_NUM ��B  ���An�1�_AUTO_ENB  �E��C��_NO�� �W�K�Am�  �*�ư�ư�ư�ưy�+Ű߿�ϟ��FLTR����HI�Sj����@��_AL�M 1X�K �2��Ƽ� +ϟ�@�����������_c�.��  �Kı�B�>ڸ@TCP_VE/R !�J!Ư	��$EXT:�_RE�Q?�薹��SI�Z�ߋ�STK�������TOL � ��DzG��{A ��_BWD�`��#���B�DI� YWJ��A��$�STEP5�G�@a��OP_DO�߶AF�ACTORY_T�UN?�d��DR_?GRP 1Z�I)��d 	9����@���x����� �n��So �k� ���+���=�N�8� q�\������������������7"
@R��Z@���?Ơ�s?*�>
 E����[>�H�8ө��E7� E??p D��� �D��Й  Cμ�	B�  ��  A@C@U�UU7UUC�>�]�>П��| EͰF@ F�5U�OL����M��Jk��K�v�H�,_�Hk�O?} ��%9tQv�8���6h�%%�O(/}�FEATU�RE [5���AHand�lingTool� v%��Eng�lish Dictionary|'�4D Stk ar�dv&~%Analo�g I/O�'�'g�le Shift��/uto Sof�tware Up�date�)mat�ic Backu�pz)1groun?d Edito |'�Camera� F��/CnrRndI�m!3X<ommon� calib U�IS3{6n:1�0Mo�nitor�;tr~t Reliab� �{(DHCPo9�:a�ta Acqui�s�3�9iagno�s1�!�;ispl�ay=1Licen�s�1�5ocume�nt Viewe��2�7ual Ch�eck Safe�ty�1&hanc�ed�6{*�EsS@F�rK0}'xt. D7IO �0fiD�Gwend�@Err�0QLB�M�Gs�Ir� �@ �y*FCTN_ Menul@v�3�WTP InPf�ac3U~%GigE�E^WU30p Mas_k Exc�@g�G�HTCPProxy� SvTD�Vigh�-Spe�@Ski�n4�U@�@mmun�ic0ons�Xu�r*PP�?�!FRconnect 2�X�ncrEPstruH�"�Z#`eJAd@JE�$KAREL C�md. L�Pua��XZcRun-TiΫ@EnvPhPel� +0s0S/W�|'5EgBSL�@Boo�k(System�)y*MACROs�,�R/Offse�� �eH�@0�?�`M�R�0�2NMech/Stop�Qt`�2"�ei�B�+Ovx�@� �0~od� wit#ch}#sA.v�{�Optm�#s�Pf�ilSL"wg�W�eulti-T�P=3z)PCM fun-g�+�o�4gB$�K�Re�gi�`r�P.�ri�L@F;���� Num� SelGu���@ Adju�P��Ɓ�*׍tatu��NJ�~%RDM Rob�ot� scove̖!+�ea��@Freq Anly�W'RemEp�An�'+�>7�Servo�@�p~{(SNPX b�bv�.SNCPCliKA<���"Libr�#Ο�k  Vt����o�`t*Pssag$�$R�a �#�ax+R�/ID]>'�MILIBP�*�?P Firm�":��P*SAcc40<;T�PTX�?(�eln��`m�+�s!�e;�or�qu� imulah�1Q1�u�pPa�a�:�30�1�s&�Pev�.'�� rid@ï�USB port- �0iP�@aL@w�?R EVNTj�|�nexcept�@`l�Y�w��H�MVC�1r�R�RKxV�0����h	����S��SC���;�SGEP�F�UI~x+Web Pl� �Ό��_�ĢP~DJAV�ZDT Applx�Ty*��EOAT6�� 4}&����!�Gri�d;�-A��iR��.�*o�AϺ"R�CP0120iC��,larm Caouse/j�ed�(�Ascii�QłL�oadS@��Upld��r?l� �1Gu�&d�)�P0B6yc� `�b��e�q@VRA/�0�@��$Jain1��r�{(NRTL���#O}nn e Heln8�/�E_.�}�z�`�tr��KROS Eth
�atI�e��j�"�$�64MB DRA9M��Q�FROZ�� �rcWeld�Pc8g�"tC5ell�,y=#sh�����c�{���� p1���ty� s ��A7W�R��p.�;k�8�A�2w-maie@ě�wM6����0qglu��pj�CP�hR�/��L��Sup���q�� �@Pcro�6����c��6@�uestF�rtcA6�x*�9/ �dv����� �///2/</i/`/ r/�/�/�/�/�/�/? ??.?8?e?\?n?�? �?�?�?�?�?O�?O *O4OaOXOjO�O�O�O �O�O�O_�O_&_0_ ]_T_f_�_�_�_�_�_ �_�_�_o"o,oYoPo bo�o�o�o�o�o�o�o �o(UL^� ������� � �$�Q�H�Z���~��� ����Ə����� � M�D�V���z������� ������I�@� R��v���������� �����E�<�N�{� r����������޿� 
��A�8�J�w�nπ� �Ϥ϶��������� =�4�F�s�j�|ߩߠ� ����������9�0� B�o�f�x������ �������5�,�>�k� b�t������������� ��1(:g^p �������  -$6cZl�� ������)/ / 2/_/V/h/�/�/�/�/ �/�/�/�/%??.?[? R?d?�?�?�?�?�?�? �?�?!OO*OWONO`O �O�O�O�O�O�O�O�O __&_S_J_\_�_�_ �_�_�_�_�_�_oo "oOoFoXo�o|o�o�o �o�o�o�oK BT�x���� �����G�>�P� }�t���������֏�� ���C�:�L�y�p� ��������ҟܟ	� � �?�6�H�u�l�~��� ����ίد����;� 2�D�q�h�z������� ʿԿ���
�7�.�@� m�d�vϣϚϬ����� �����3�*�<�i�`� rߟߖߨ��������� �/�&�8�e�\�n�� ������������+� "�4�a�X�j������� ����������'0 ]Tf����� ���#,YP b������� �//(/U/L/^/�/ �/�/�/�/�/�/�/? ?$?Q?H?Z?�?~?�? �?�?�?�?�?OO O MODOVO�OzO�O�O�O �O�O�O_
__I_@_ R__v_�_�_�_�_�_ �_oooEo<oNo{o ro�o�o�o�o�o�o A8Jwn� �������� =�4�F�s�j�|����� ͏ď֏����9�0� B�o�f�x�����ɟ���ҟ�����5�,�V��  H55�2F�l�21r�R7�8q�50r�J61�4r�ATUP��5�45��6r�VCA�Mr�CRIѧUI�F��28ҦNREv~�52ŦR63}�wSCHr�LIC��DOCV2�CSU�~�869��0��E�IOC�4q�R6=9ŦESET��ħ�J7ħR68}�M�ASKr�PRXY��7r�OCO��3Ю�q�����3ٶJ6֔�53U�H�LC�H��OPLG��0^�MHCR¶SP��MCS��0��55���MDSW���OP�MPR����0��PCM�R0`�ǚ���Z��51���51�0��PRSv��69ٶFRDѦ�FREQ~�MCN�r�93��SNBA���SHLB~�M�����2��HTC���TMIL~�U�T{PAm�TPTX��#ELq�Z�U�8�����}�J95��TUTv�95ٶUEV��wUEC��UFRѦ�VCCy�Oi�VI�P��CSC�CS�G�G�Ir�WEBn��HTT��R6��#誠��CG��IG���IPGS
�RCv��DG�H84���R66��R7��Rn�R53�68�E2�RȂ��4i��66E�4}�NVDv��R6\�R84��D0��F��AWS�ѧLI�ȸ�CMS�m�2 ��STY��T�O��7T�NNٶO�RSi�J�?�O]L@END~�L��S{FVRm�M�� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/�Z#  Hg552V'p!21v)�R78u,50v)J�614v)ATUP��*545�,6v)VwCAMv)CRI�+�UIF�+28�*N�RE�*52�*R6�3�+SCHv)LI�C5:DOCVv:C�SU�*869�+0^�*EIOC6;4u*�R69�*ESET��+�+J7�+R68ޅ*MASKv)PR�XY<7v*OCOB�<3�,u*@�,3UJ[J6�,53�:H�L�LCH5JOPLGz�+0uJMHCR6J]S�KMCS�,0K{55�*MDSWV[vdKOPdKMPReJtR0�L0�*PCM:�R0�[@�*P�K5�1�+51�\0�*P�RS�;69UJFR�D�*FREQ�*M�CNv*93�*SN�BAF;�KSHLB��jM�kR0E\2�*H{TC�*TMIL�,�:TPA�:TPT�X�jELujP�;8��+� �*J95%:T�UTeK95UJUE�V�:UEC5JUF]R�*VCC�|OZwVIPzCSC5z�CSG5:�0Iv)W�EB�*HTT�*Ra6D<c|� 5�CGT�{IG4�IPGS���RCzDGdKH8�4�*R66�*R7��;R�\R53�[68�\2uJR�L�0�\�4�66�4�*N�VD�:R6[R8�4uJD0��FӜA�WS�+LI�\�+C�MS�:"��*STY��TOU�7�<NN.UJORSZJ��&Jv3lOL4�END�*uL�{S��FVR�9 U(��� �2�D�V�h� z�������¿Կ��� 
��.�@�R�d�vψ� �ϬϾ��������� *�<�N�`�r߄ߖߨ� ����������&�8� J�\�n������� �������"�4�F�X� j�|������������� ��0BTfx ������� ,>Pbt�� �����//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?O O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h� zߌߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N�`�r������� ��������&8 J\n����� ���"4FX j|������@�//0/B/R)^ �STDY$LANGz$u)�/�/ �/�/�/�/�/??/? A?S?e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O�O �O__'_9_K_]_o_ �_�_�_�_�_�_�_�_ o#o5oGoYoko}o�o �o�o�o�o�o�o�1zRBTy&OPTNN`r����|��DPNx$ �� �2�D�V�h�z�������Q(��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬϾ����� ����*�<�N�`�r� �ߖߨߺ�������� �&�8�J�\�n��� ������������"� 4�F�X�j�|������� ��������0B Tfx����� ��,>Pb t������� //(/:/L/^/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�? �?�?�?�?�?O O2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�o�o�o�o�o�o &8J\n�� �������"� 4�F�X�j�|������� ď֏�����0�B� T�f�x���������қ�՟���)�;�M��99T��$FE�AT_ADD ?_	�������?  	Q��� ����ȯگ����"� 4�F�X�j�|������� Ŀֿ�����0�B� T�f�xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo�tot�DEMO �[��    Q��m�o�o�o�o�o& /\Se�� �����"��+� X�O�a�{��������� �ߏ���'�T�K� ]�w����������۟ ���#�P�G�Y�s� }��������ׯ�� ��L�C�U�o�y��� ����ܿӿ��	�� H�?�Q�k�uϢϙϫ� ���������D�;� M�g�qߞߕߧ����� ��
���@�7�I�c� m����������� ���<�3�E�_�i��� ������������ 8/A[e��� �����4+ =Wa����� ���/0/'/9/S/ ]/�/�/�/�/�/�/�/ �/�/,?#?5?O?Y?�? }?�?�?�?�?�?�?�? (OO1OKOUO�OyO�O �O�O�O�O�O�O$__ -_G_Q_~_u_�_�_�_ �_�_�_�_ oo)oCo Mozoqo�o�o�o�o�o �o�o%?Iv m������ ��!�;�E�r�i�{� ������ޏՏ��� �7�A�n�e�w����� ��ڟџ����3� =�j�a�s�������֯ ͯ߯���/�9�f� ]�o�������ҿɿۿ ����+�5�b�Y�k� �Ϗϡ���������� �'�1�^�U�gߔߋ� �������� ���	�#� -�Z�Q�c������ ����������)�V� M�_������������� ����%RI[ ������� �!NEW�{ �������/ /J/A/S/�/w/�/�/ �/�/�/�/�/??F? =?O?|?s?�?�?�?�? �?�?�?OOBO9OKO xOoO�O�O�O�O�O�O �O__>_5_G_t_k_ }_�_�_�_�_�_�_o o:o1oCopogoyo�o �o�o�o�o�o�o	6 -?lcu��� �����2�)�;� h�_�q�������ԏˏ ݏ���.�%�7�d�[� m�������Пǟٟ� ��*�!�3�`�W�i��� ����̯ïկ���&� �/�\�S�e������� ȿ��ѿ���"��+� X�O�aώυϗ��ϻ� ��������'�T�K� ]ߊ߁ߓ��߷����� ����#�P�G�Y�� }����������� ��L�C�U���y��� ����������	 H?Q~u��� ���D; Mzq����� �
///@/7/I/v/ m//�/�/�/�/�/? �/?<?3?E?r?i?{? �?�?�?�?�?O�?O 8O/OAOnOeOwO�O�O �O�O�O�O�O_4_+_ =_j_a_s_�_�_�_�_ �_�_�_o0o'o9ofo ]ooo�o�o�o�o�o�o �o�o,#5bYk �������� (��1�^�U�g����� ����������$�� -�Z�Q�c��������� ����� ��)�V� M�_������������ ݯ���%�R�I�[� ����������ٿ� ��!�N�E�Wτ�{� �ϧϱ��������� �J�A�S߀�w߉ߣ� �����������F��=�O�|�s��  ����������� �!�3�E�W�i�{��� ������������ /ASew��� ����+= Oas����� ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e�w������� ��џ�����+�=� O�a�s���������ͯ ߯���'�9�K�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�i  �h�a�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�w��� ������џ����� +�=�O�a�s������� ��ͯ߯���'�9� K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� �-�?�Q�c�u��� �����������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ� ����������'�9� K�]�o߁ߓߥ߷��� �������#�5�G�Y� k�}���������� ����1�C�U�g�y� ��������������	 -?Qcu�� �����) ;M_q���� ���//%/7/I/ [/m//�/�/�/�/�/ �/�/?!?3?E?W?i? {?�?�?�?�?�?�?�? OO/OAOSOeOwO�O �O�O�O�O�O�O__ +_=_O_a_s_�_�_�_ �_�_�_�_oo'o9o@Ko]ooo�o�o�a�`�h�o�o�o�o );M_q��� ������%�7� I�[�m��������Ǐ ُ����!�3�E�W� i�{�������ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳����� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q��� ����%7 I[m���� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q������� ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ�������� �+�=�O�a�s߅ߗ� �߻���������'�9�K�]�o������$FEAT_DEMOIN  �䫀�������I�NDEX�������ILECOMP \���������SETUP2 ]����  N� @���_AP2B�CK 1^� � �)��t���%j����������� i�����"��/X�� |��A�e� �0�Tf�� �=��s/� ,/>/�b/��/�/'/ �/K/�/�/�/?�/:? �/G?p?�/�?#?�?�? Y?�?}?O$O�?HO�? lO~OO�O1O�OUO�O �O�O _�OD_V_�Oz_ 	_�_�_?_�_c_�_
o �_.o�_Ro�__o�oo �o;o�o�oqo�o* <�o`�o��%� I�m���8�� \�n����!���ȏW� �{��"���F�Տj����w����N�PR�� 2g�*.VR���_�*���\�0 �D�.�ېPCL�u�>_�FR6:`���0�ůT�T���������%��දK�-�G*.Fޟ|�^�	���j���8�Ϳ\�ST�Mؿω����-���Q�\�Hτ��r�p/�A���]�GIF�π
���ϳ���Z�]�JPGdߎ��z�7�Iߌ��U�JS���_�����߼�%
JavaScript=�h�CS.��Ƃ�?�� %Casca�ding Sty�le Sheet�s��3�
ARGN?AME.DT��S��\���$�4�E����4�DISP*;�Q�0��I�[�����u�
TPEIN�S.XML�� �:�\��,�Cust�om Toolb�arM|�PASS�WORD��Q�F�RS:\�O��P�assword ?Config�,� �P��t� �9�]�/�(/ �L/���//�/5/ �/�/k/ ?�/$?6?�/ Z?�/~?�??�?C?�? g?y?O�?2O�?+OhO �?�OO�O�OQO�OuO 
__�O@_�Od_�O_ �_)_�_M_�_�_�_o �_<oNo�_roo�o�o 7o�o[o�oo�o&�o J�oC��3� �i��"�4��X� �|�����A�֏e� Ϗ���0���T�f��� �������O��s�� ����>�͟b��[��� '���K��򯁯��� :�L�ۯp�����#�5� ʿY��}��$ϳ�H� ׿l�~�Ϣ�1����� g��ϋ� ߯���V��� z�	�s߰�?���c��� 
��.��R�d��߈� ��;�M���q���� ��<���`������%� ��I��������8 ����n���!�� W�{"�F� j|�/�Se ��/�/T/�x/ /�/�/=/�/a/�/? �/,?�/P?�/�/�?i6��$FILE_D�GBCK 1^���s0��� < �)
�SUMMARY.�DG�?<<MD:��?OH0Dia�g Summar�yO:
CONSLOG�?�?�1HO�O�AConsol�e log�O;	?TPACCN~O�O�%�O_ETP �Accounti�n�O:FR6:�IPKDMP.ZIP<_@8
T_�_E�$PExcepti�on�_B[�0MEMCHECK�OeO�?�o�AMemor?y Dataoi6�4n )�QRI�PE{O�_�_�o#c�%[a Pack�et L�Oj4L��$��R[aSTAT��ouo�o %��bStatus<�k	FTP_ot�xg�Amme?nt TBD��g� >I)ETHERNE�oy�Q��$�AEther�n�`�@figur�a�_4�qDCSV�RF�{���-s�k� verify� all��j3M{4f�DIFF�������+��c��dif�f-���Qk�CHG01"�	����/qC�,؟�2�n�2����@��4�?�՟�u�3*�8�#��� J�߯�n�VTRNDIAG.LS䯕����<�'a�� Ope�L��a Anost�icIg��)�VDEV �DAT�=��,�>�0pVi�s_�Devicef�s�IMG ��_��譿BϩcشIma�g�q�UP��E�S���FRS:�\����AUpd�ates Lis�t��:0�FLEXEVEN�!�3��L�/q� UIF� Ev�q�oj2-�vZ)
PSRB?WLD.CMx�<<����ϝ@PS_ROBOWEL�X�:GIG^o+�6�|O�"fGigEh��r�j2N�@�)>@�HADOWJ�/��A���%cShad�ow Chang�e>Ke(dt��RCMERR������Z�%c�CFG �Errorްta�il�� a���cCMSGLIB R�9�K���g��8r���ic�����)��ZD�:��^!g7ZD{�ad ��{ ��NOTIp��=O�#eNot�ificM��j5,�AG?;B?_f? l�?�H��~ /�7/I/�m/��/ �/2/�/V/�/z/�/!? �/E?�/i?{?
?�?.? �?�?d?�?�?O/O�? SO�?wOO�O�O<O�O `O�O_�O+_�OO_a_ �O�__�_�_J_�_n_ o�_o9o�_]o�_�o �o"o�oFo�o�o|o �o5G�ok�o� ��T�x��� C��g�y����,��� ӏb��������(�Q� ��u������:�ϟ^� ����)���M�_�� �����6���ݯl�� ��%�7�Ư[�����  ���D�ٿ�z�Ϟ� 3�¿@�i�����ϱ� ��R���v��߬�A� ��e�w�ߛ�*߿�N� ���߄���=�O��� s����8���\��� ���'���K���X��� ���4�����j����� #5��Y��}� �B�f��1 �Ug���� P�t	//�?/��c/�p/�/z#�$F�ILE_FRSP�RT  ���� �����(MDONLY �1^�%z  
� �)MD:_�VDAEXTP.�ZZZ�/Q/(?7;�6%NO B�ack filey ?z$S�6P./ �??�?v/�?�?(/O �?+O=O�?aO�?�O�O &O�OJO�O�O�O_�O 9_�OF_o_�O�_"_�_ �_X_�_|_o#o�_Go �_ko}oo�o0o�oTo �o�o�o�oCU�o y��>�b��	��$VISBCK��(�!�#*.VD�
�T��pFR:\�#�ION\DAT�A\?��r�pV�ision VD U2���ȏڏ���� "���3�X��|���� ��A�֟e�������0� ��T�f�!������=� ���s����,�>�ͯ b�񯆿�'���K�� 򿭿ϥ�:�ɿK�p� ����#ϸ���Y���}��ߡϳ�Hߨ*LUI�_CONFIG �_�%6�S� $ 1��#�߰����������
��$$ |x:�<�N�`�r�� ��*����������� �5�G�Y�k�}���� ������������1 CUgy��� ����-?Q cu����� ��/)/;/M/_/q/ /�/�/�/�/�/�/�/ ?%?7?I?[?�/l?�? �?�?�?�?p?�?O!O 3OEOWO�?{O�O�O�O �O�OlO�O__/_A_ S_�Ow_�_�_�_�_�_ h_�_oo+o=oOo�_ so�o�o�o�o�odo�o '9K�oo� ���N���� #�5��Y�k�}����� ��J�׏�����1� ȏU�g�y�������F� ӟ���	��-�ğQ� c�u�������B�ϯ� ���)���M�_�q� ������>�˿ݿ�� Ϫ�$�I�[�m�ϑ� (ϵ���������ߦ� 3�E�W�i�{ߍ�$߱� ����������/�A� S�e�w�� ����� �������+�=�O�a� s��������������|��  x��$FLUI_�DATA `����L���>RESUL�T 2aLu ? �T��+� ������! 3EWi��~�� �����/!/3/�E/W/i/{/�-?��0���L�/�+����/�/??,?>? P?b?t?�?�?�?�?{ �/�?�?
OO.O@ORO�dOvO�O�O�O�O�� O �/�G�/_�/+_=_ O_a_s_�_�_�_�_�_ �_�_oo&_9oKo]o oo�o�o�o�o�o�o�o �o�O2�OV_} �������� �1�C�U�g�&o���� ����ӏ���	��-� ?�Q�c�"��F��j l�����)�;�M� _�q���������x�ݯ ���%�7�I�[�m� �������t�ֿ���� �Я3�E�W�i�{ύ� �ϱ����������ʯ /�A�S�e�w߉ߛ߭� ���������ƿ�� 4�^� υ������ ������'�9�K�]� ߁������������� ��#5GY�b� <��r���� 1CUgy�� �n����	//-/ ?/Q/c/u/�/�/�/j |��?�)?;?M? _?q?�?�?�?�?�?�? �?O�%O7OIO[OmO O�O�O�O�O�O�O�O _�/�/�/T_?{_�_ �_�_�_�_�_�_oo /oAoSoOwo�o�o�o �o�o�o�o+= Oa _2_D_�h_� ����'�9�K�]� o�������do��ۏ� ���#�5�G�Y�k�}� ������rԟ���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ���ğ&��J� �qσϕϧϹ����� ����%�7�I�[�� ߑߣߵ��������� �!�3�E�W��x�:� ��^�`��������� /�A�S�e�w������� l�������+= Oas���h�� ��� ��'9K] o������� ���#/5/G/Y/k/}/ �/�/�/�/�/�/�/� �(?R?y?�?�? �?�?�?�?�?	OO-O ?OQO/uO�O�O�O�O �O�O�O__)_;_M_ ?V?0?z_�_f?�_�_ �_oo%o7oIo[omo o�o�obO�o�o�o�o !3EWi{� �^_p_�_�_��_� /�A�S�e�w������� ��я����o�+�=� O�a�s���������͟ ߟ�����H�
� o���������ɯۯ� ���#�5�G��k�}� ������ſ׿���� �1�C�U��&�8��� \���������	��-� ?�Q�c�u߇ߙ�X��� ��������)�;�M� _�q����f���� ����%�7�I�[�m� ��������������� �!3EWi{� �������� ��> �ew��� ����//+/=/ O/s/�/�/�/�/�/ �/�/??'?9?K?
 l?.�?RT?�?�?�? �?O#O5OGOYOkO}O �O�O`/�O�O�O�O_ _1_C_U_g_y_�_�_ \?�_�?�_�_�Oo-o ?oQocouo�o�o�o�o �o�o�o�O);M _q������ ��_�_�_�F�om� �������Ǐُ��� �!�3�E�i�{��� ����ß՟����� /�A� �J�$�n���Z� ��ѯ�����+�=� O�a�s�����V���Ϳ ߿���'�9�K�]� oρϓ�R�d�v����� ���#�5�G�Y�k�}� �ߡ߳������ߨ�� �1�C�U�g�y��� ��������������� <���c�u��������� ������);�� _q������ �%7I�� ,��P������ /!/3/E/W/i/{/�/ L�/�/�/�/�/?? /?A?S?e?w?�?�?Z �?~�?�OO+O=O OOaOsO�O�O�O�O�O �O�OO_'_9_K_]_ o_�_�_�_�_�_�_�_ �?o�?2o�?Yoko}o �o�o�o�o�o�o�o 1C_gy�� �����	��-� ?��_`�"o��FoH��� Ϗ����)�;�M� _�q�����T��˟ݟ ���%�7�I�[�m� ���P���t�֯诬� �!�3�E�W�i�{��� ����ÿտ翦��� /�A�S�e�wωϛϭ� �����Ϣ��Ư�:� ��a�s߅ߗߩ߻��� ������'�9���]� o����������� ���#�5���>��b� ��N߳��������� 1CUgy�J� �����	- ?Qcu�F�X�j� |����//)/;/M/ _/q/�/�/�/�/�/�/ �??%?7?I?[?m? ?�?�?�?�?�?�?� ��0O�WOiO{O�O �O�O�O�O�O�O__ /_�/S_e_w_�_�_�_ �_�_�_�_oo+o=o �?O O�oDO�o�o�o �o�o'9K] o�@_����� ��#�5�G�Y�k�}� ��No��roԏ�o��� �1�C�U�g�y����� ����ӟ���	��-� ?�Q�c�u��������� ϯᯠ��ď&��M� _�q���������˿ݿ ���%�7���[�m� ϑϣϵ��������� �!�3��T��x�:� <߱����������� /�A�S�e�w��Hϭ� ����������+�=� O�a�s���Dߦ�h��� ����'9K] o�������� �#5GYk} ����������� /./��U/g/y/�/�/ �/�/�/�/�/	??-? �Q?c?u?�?�?�?�? �?�?�?OO)O�2/ /VO�OB/�O�O�O�O �O__%_7_I_[_m_ _>?�_�_�_�_�_�_ o!o3oEoWoio{o:O LO^OpO�o�O�o /ASew��� ���_���+�=� O�a�s���������͏ ߏ�o�o�o$��oK�]� o���������ɟ۟� ���#��G�Y�k�}� ������ůׯ���� �1�����v�8��� ����ӿ���	��-� ?�Q�c�u�4��ϫϽ� ��������)�;�M� _�q߃�B���f��ߊ� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� �������������� ��ASew��� ����+�� Oas����� ��//'/��H/
 l/.0/�/�/�/�/�/ �/?#?5?G?Y?k?}? <�?�?�?�?�?�?O O1OCOUOgOyO8/�O \/�O�O�?�O	__-_ ?_Q_c_u_�_�_�_�_ �_�?�_oo)o;oMo _oqo�o�o�o�o�o�O �O�O�o"�OI[m ������� �!��_E�W�i�{��� ����ÏՏ����� �o& J�t�6���� ��џ�����+�=� O�a�s�2�������ͯ ߯���'�9�K�]� o�.�@�R�d�ƿ��� ���#�5�G�Y�k�}� �ϡϳ��τ������ �1�C�U�g�yߋߝ� �����ߒ������ڿ ?�Q�c�u����� ����������;�M� _�q������������� ��%�����j ,������� !3EWi(�z ������// //A/S/e/w/6�/Z �/~�/�/??+?=? O?a?s?�?�?�?�?�? �/�?OO'O9OKO]O oO�O�O�O�O�O�/�O �/_�/5_G_Y_k_}_ �_�_�_�_�_�_�_o o�?CoUogoyo�o�o �o�o�o�o�o	�O <�O`"_$��� �����)�;�M� _�q�0o������ˏݏ ���%�7�I�[�m� ,��P��ğ����� �!�3�E�W�i�{��� ����ï������� /�A�S�e�w������� ��~�ȟ����؟=� O�a�sυϗϩϻ��� ������ԯ9�K�]� o߁ߓߥ߷������� ���п���>�h�*� ������������� �1�C�U�g�&ߋ��� ����������	- ?Qc"�4�F�X� |���);M _q����x�� �//%/7/I/[/m/ /�/�/�/�/��� ?�3?E?W?i?{?�? �?�?�?�?�?�?O� /OAOSOeOwO�O�O�O �O�O�O�O__�/�/ �/^_ ?�_�_�_�_�_ �_�_oo'o9oKo]o Ono�o�o�o�o�o�o �o#5GYk*_ �N_�r_���� �1�C�U�g�y����� ��������	��-� ?�Q�c�u��������� |ޟ���)�;�M� _�q���������˯ݯ ���ҏ7�I�[�m� �������ǿٿ��� �Ο0��T��ύ� �ϱ����������� /�A�S�e�$��ߛ߭� ����������+�=� O�a� ς�DϦ��|� ������'�9�K�]� o���������v����� ��#5GYk} ���r����
 ��1CUgy�� �����	/��-/ ?/Q/c/u/�/�/�/�/ �/�/�/?��2? \?�?�?�?�?�?�? �?OO%O7OIO[O/ O�O�O�O�O�O�O�O _!_3_E_W_?(?:? L?�_p?�_�_�_oo /oAoSoeowo�o�o�o lO�o�o�o+= Oas����z_ �_�_ ��_'�9�K�]� o���������ɏۏ� ���o#�5�G�Y�k�}� ������şן���� ���R��y����� ����ӯ���	��-� ?�Q��b��������� Ͽ����)�;�M� _����B���f����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ���p�������� /�A�S�e�w������� ����������+= Oas����� ����$��H
� ������� �/#/5/G/Y/}/ �/�/�/�/�/�/�/? ?1?C?U?v?8�? �?p/�?�?�?	OO-O ?OQOcOuO�O�O�Oj/ �O�O�O__)_;_M_ __q_�_�_�_f?�?�? �_�_�?%o7oIo[omo o�o�o�o�o�o�o�o �O!3EWi{� �������_o �_&�P�ow������� ��я�����+�=� O�s���������͟ ߟ���'�9�K�
� �.�@���d�ɯۯ� ���#�5�G�Y�k�}� ����`�ſ׿���� �1�C�U�g�yϋϝ� ��n������϶��-� ?�Q�c�u߇ߙ߽߫� �����߲��)�;�M� _�q��������� ���������F��m� ��������������� !3E�V{� ������ /AS�t6��Z� ����//+/=/ O/a/s/�/�/�/��/ �/�/??'?9?K?]? o?�?�?�?d�?��? �O#O5OGOYOkO}O �O�O�O�O�O�O�O�/ _1_C_U_g_y_�_�_ �_�_�_�_�_�?o�? <o�? ouo�o�o�o�o �o�o�o);M _q������ ���%�7�I�oj� ,o����dǏُ��� �!�3�E�W�i�{��� ��^ß՟����� /�A�S�e�w�����Z� ��~�ȯ򯴏�+�=� O�a�s���������Ϳ ߿񿰟�'�9�K�]� oρϓϥϷ������� ����Я�D��k�}� �ߡ߳���������� �1�C��g�y��� ����������	��-� ?����"�4ߖ�X߽� ������);M _q��T��� �%7I[m ��b�t������ /!/3/E/W/i/{/�/ �/�/�/�/�/�?? /?A?S?e?w?�?�?�? �?�?�?�?���:O �aOsO�O�O�O�O�O �O�O__'_9_�/J_ o_�_�_�_�_�_�_�_ �_o#o5oGoOho*O �oNO�o�o�o�o�o 1CUgy�� �o����	��-� ?�Q�c�u�����Xo�� |oޏ�o��)�;�M� _�q���������˟ݟ �%�7�I�[�m� �������ǯٯ믪� �Ώ0����i�{��� ����ÿտ����� /�A� �e�wωϛϭ� ����������+�=� ��^� ��ߔ�Xϻ��� ������'�9�K�]� o���RϷ������� ���#�5�G�Y�k�}� ��Nߘ�r߼����� 1CUgy�� ������	- ?Qcu���� ��������/8/�� _/q/�/�/�/�/�/�/ �/??%?7?�[?m? ?�?�?�?�?�?�?�? O!O3O�//(/�O L/�O�O�O�O�O__ /_A_S_e_w_�_H?�_ �_�_�_�_oo+o=o Ooaoso�o�oVOhOzO �o�O'9K] o�������_ ��#�5�G�Y�k�}� ������ŏ׏鏨o�o �o.��oU�g�y����� ����ӟ���	��-� �>�c�u��������� ϯ����)�;��� \����B�����˿ݿ ���%�7�I�[�m� ϑϢ����������� �!�3�E�W�i�{ߍ� L���p��ߔ����� /�A�S�e�w���� ���������+�=� O�a�s����������� ���� ��$����] o������� �#5��Yk} �������/ /1/��R/v/�/L �/�/�/�/�/	??-? ??Q?c?u?�?F�?�? �?�?�?OO)O;OMO _OqO�OB/�/f/�O�O �/__%_7_I_[_m_ _�_�_�_�_�_�?�_ o!o3oEoWoio{o�o �o�o�o�o�O�O�O ,�OSew��� ������+��_ O�a�s���������͏ ߏ���'��o�o
 ~�@����ɟ۟� ���#�5�G�Y�k�}� <�����ůׯ���� �1�C�U�g�y���J� \�n�п����	��-� ?�Q�c�uχϙϫϽ� �ώ�����)�;�M� _�q߃ߕߧ߹����� ������"��I�[�m� ������������ �!���2�W�i�{��� ������������ /��P�t6�� ����+= Oas����� ��//'/9/K/]/ o/�/@�/d�/��/ �/?#?5?G?Y?k?}? �?�?�?�?�?��?O O1OCOUOgOyO�O�O �O�O�O�/�O�/_�/ �OQ_c_u_�_�_�_�_ �_�_�_oo)o�?Mo _oqo�o�o�o�o�o�o �o%�OF_j |@o������ �!�3�E�W�i�{�:o ����ÏՏ����� /�A�S�e�w�6�Z ��Ο�����+�=� O�a�s���������ͯ �����'�9�K�]� o���������ɿ��ҟ ���� ��G�Y�k�}� �ϡϳ���������� �ޯC�U�g�yߋߝ� ����������	��ڿ ����r�4ϙ��� ��������)�;�M� _�q�0ߕ��������� ��%7I[m >�P�b������ !3EWi{� �������// //A/S/e/w/�/�/�/ �/�/���?�=? O?a?s?�?�?�?�?�? �?�?OO�&OKO]O oO�O�O�O�O�O�O�O �O_#_�/D_?h_*? �_�_�_�_�_�_�_o o1oCoUogoyo�_�o �o�o�o�o�o	- ?Qcu4_�X_� |_����)�;�M� _�q���������ˏ�o ���%�7�I�[�m� �������ǟ�蟪 ��ПE�W�i�{��� ����ïկ����� ܏A�S�e�w������� ��ѿ�����؟:� ��^�p�4��ϩϻ��� ������'�9�K�]� o�.��ߥ߷������� ���#�5�G�Y�k�*� t�NϘ��������� �1�C�U�g�y����� ����������	- ?Qcu���� |�������;M _q������ �//��7/I/[/m/ /�/�/�/�/�/�/�/ ?���f?(�? �?�?�?�?�?�?OO /OAOSOeO$/�O�O�O �O�O�O�O__+_=_ O_a_s_2?D?V?�_z? �_�_oo'o9oKo]o oo�o�o�o�ovO�o�o �o#5GYk} �����_�_�_
� �_1�C�U�g�y����� ����ӏ���	��o� ?�Q�c�u��������� ϟ�����8���\�j��$FMR2_GRP 1bj��� �C4  B�#�	 #��������E�� E�  �F@ F�5U�ܥ���L���M���Jk�K��v�H�,�H�k��?�  x ����9tQvH��8���6h�%<T��A�  p����BH��B��������@�����ʿ۽^��@UUU�U��۽>�]�>П���;r8	=�==E��<D��><�ɳ<��Ε�:�b�:�/'79�W�9�
@�8�8�9�ϑ�ܿ�������E7� E?p� D������D��  D�  C����#�~�_CFG {c��T ��[�m��!�NO ���
F0�� ��� �RM_CHK?TYP  {�#�p����K�}�ROM���_MIN��#��������X~�SS�B1�dj� ��/�#�&�O��a�'�TP_DEF�_OW  #�|��v�IRCOM������$GENOV_RD_DO��-�n��THR�� d��d��_ENB�� ���RAVC��e��#� �ȥF�nH E�� G�a H�� H�@Jh`�ψK�|�������� [��OU��k��������⸥<��2���&TV#�C�������j@)�#������p����h��SMT���l(���%�y�$HoOSTC1�1m��n$��-� 	OMOO#� �e����/ *�3/E/W/i/��/�  	anonymous�/�/�/�/�/? N`rO?�/� "/�?�?�?�?/�?O O'O9O\?�/�/�O�O �O�O�O?"?4?F?HO 5_|?Y_k_}_�_�_�? �_�_�_�_o0_fOxO Uogoyo�o�o�O�O_ �oo	P_-?Qc �_t�����o� :o�)�;�M�_��o�o �o�o������ %�7�~[�m������ Ə������!�3� z�����L������ï կ������/�A�S� e�����П����ѿ� ��<�N�`�r�Oφ��� �ϗϩϻ������� �'�9�\ϒ����ߓ� �߷����"�4�F�H� 5�|�Y�k�}����� ����������f�C��U�g�y����1EN�T 1n�� P�!���  �  ����,��Pt 7�[����� �:�^!3� W�{�� /�� 6/�Z//~/A/�/e/ �/�/�/�/�/ ?�/D? ?P?+?y?�?a?�?�? �?�?
O�?.O�?OdO�'O�OKO�OoJQUICC0�O�O�O_��D1	_�O�OX_�D2�Y_5_G_�_!ROUTER�_�_�_�_!PCJOG�_��_!192.�168.0.10��O�CCAMPRT,Io%o!9e1B`po�WfRT�_to�o�o �!Softwa�re Opera�tor Pane�l�o6o7��NAM�E !��!R�OBObo?S_C�FG 1m�� ��Aut�o-starte�d��FTP�� �q���H��1�C� U�g��������� ҏx�	��-�?�Q��#��֩����� ������(��L� ^�p�������9�ʯܯ � ��$�������� ����ן��ƿؿ��� ï �2�D�V�hϋ�� �ϰ���������?�Q� c�@�w�d߫��ߚ߬� �߅�������*�M� ��I�r������ �%�7�9�&�m�J�\� n�����Y�������� ��!���4FXj| ���������A� 0BT�� ����w//,/ >/P/������/ �/�/??(?�L? ^?p?�?�?�/9?�?�? �? OO$Ok/}/�/=O �?�O�/�O�O�O�O�O �? _2_D_V_yOz__��_�_�_�_�_zNp_?ERR oXz�_�fPDUSIZ � �P^�@�d�>6eWRD ?��uhA�  ?guest�Vvo��o�o�o�o�oGtSC�DMNGRP 2�p�u `��hA�P���VKt �	P01.05� 8MA   
��  3  Y�MpLpٝ�CK� ���U��?�����3uptp?�'����]}$oЦ���wDp�����Mp�Z@Z@U~]�����t�pup���Hp�}[�5�li@6i@	I=��zdASew��k_GROU pq*ip�b	�a8q�4��QUPD  �dEe���TYꌐm`TTP�_AUTH 1r�k <!iP�endan�gR���_��!KARE�L:*R�[�m�KC������z�ݟ˟�� �q�@��)�v�M�_� ����������˯ݤ!�CTRL sm�q>��Q
�QF�FF9Eh�\�hB�FRS:DEFA�ULT`�FA�NUC Web ?Server`�N� >�!�^opd	�ֿ������0�dWR_C�ONFIG t�{ `�aID�L_CPU_PC���QB�i@�� ;BH��MIN��Na~��GNR_IOa�Db�Ph��NPT_�SIM_DO�����STAL_SC�RN�� ���IN�TPMODNTOqL��˻�RTY��ܢ���VIS%�EN�B�����OLN/K 1ukr`�߀�����������M�ASTE���SLAVE vo�E�RAMCACH�E4�,�O'�O_CcFGv�ӎ�UO�����CMT_OPp���j��YCLu����y�_ASG 19wwPa
 �;� M�_�q����������������% ��N�UMCci
��I�Ps��RTRY_CN�����Cc����e �����x�T�j`�j`��P�?=�T� ��	�* <N`r��� ����/�,/>/ P/b/t/�//�/�/�/ �/�/?�/�/:?L?^? p?�?�?#?�?�?�?�?  OO�?6OHOZOlO~O �OO1O�O�O�O�O_  _�OD_V_h_z_�_�_ -_�_�_�_�_
oo�_ �_Rodovo�o�o�o;o �o�o�o*�oN `r���7I� ���&�8��\�n� ��������E�ڏ��� �"�4�ÏՏj�|��� ����ğS������ 0�B�џf�x������� ��O�a�����,�>� P�߯t���������ο ]����(�:�L�ۿ �ϔϦϸ�����k�  ��$�6�H�Z���~� �ߢߴ�����g�y��  �2�D�V�h��ߌ�� ��������u�
��.� @�R�d���������� ��������*<N�`r�_MEMBERS 2y��   u$�������	� RCA_�ACC 2z��   �[� V�5;ڀ"  �'!+C��B�UF001 2{�= �u0�  u0�(�N��s������V���2�X�U}��������$8$`$��$�$�$���� 9$F9$l�  �:�W"�  o��k���i$5�i$ݙ��$������� %ȭ � �%�$J�$p��$��$��$��U	�$.�$S�$y�$e��$��$ $�4U74]4�4�4��4���I4E�I4jI4�I4�I4��v2�����2 ��2��2��2��2 ����2��2��2 ��2��2��2  � !B B B  B ( B0 B8 �?!DB H DBP �W!Y!_!a! g!�o!tBx tB� � �!�B�4�!�B�4�!�! �!�B� �B� �B� �B � �B� ��!�B� �B � �B� �B 0�B0�B 	D1R 0R(0R00 R80R@0RH0�O1 TRX0TR`0TRh0TRp0TRx0�v3�?��3 �R��3�R��3�R� �3�R��3�R��3�R �C#Cb"&C b("6Cb8"FCMbH" VCdBgBg#vCub x"�C�#�C�b�T�# �C�b�"�C�b�"�C�b �"�C�#�C�b�"�C �b 2S�bd3&S%r (26S%r82FS%rH2VS ]rX2fS]rh2vS]rx2~tCFG 2|� 4 � �zJ < �t�qr�HIS�~ �� 2025�-12-�0 ;~7�I�[�m���������Ǐ0��l�1� ��$�6��H�Z�l�~��7�  �!��!��l"���� ������ 	��-�?�Q�c�u��� ��П��ϯ���� )�;�M�_��������� ��˿ݿ���%�7� n���m�ϑϣϵ��� �������F�X�j�W� i�{ߍߟ߱������߀��v�0���%�d ��^�p������� ����܏�$�6�H�Z� l�~�������6Iᤐ H⬐HⴐH�0�B� ,>Pbt�� �������( :L^p���� ��� //$/6/H/ Z/��g/�/�/�/�/ �/�/? ?2?i/{/�/ z?�?�?�?�?�?�?�? 
O���w�P�)��qO �O�O�O�O�O�O�O_ _��I_[_m__�_ �_�_�_�� P���b S ��N?`?&o8oJo\ono �o�o�o�o�oJ?o�o "4FXj|� ��o�o�o���� 0�B�T�f�x����� ��ҏ�����,�>� P�b�����������Ο������(�:��I_CFG 2=K� H
Cycle Timev��Busyp�I�dl}�t�minz@���Upy��w�Read���Dow���� ���t�Count>w�	Num t�u���l�#� P���P�ROGZ��=EG@�3�x����������ҿ��E�SDT_�ISOLC  �=I� ��J2�3_DSP_EN�B  ˳�.�INC �>� S��A   ?�  �=���<#�
|�u�:�o ����ϫ� Q����'�OB�N�C7���`���G�_GROUP 1݂�<��<A��s�Y9���?Xg�x� PQ�߳��߀�ߖ�����1� W�����G_IN_A�UTO��B�POS�RE���KANJ?I_MASK��^����RELMON #�=K+� Ry����!�3�E�W����R��Y�I� Ty���J��KCL_Lo�NU�M;���$KEYL?OGGING��B@�-�F�I�LANGUAGE =E� �DEF�AULT #+AL�G[��Y���� Qxl��P8��H�  � P'0X�W 
� Q� P޿��;��
�(�UT1:\g�� ������0GTfx� R(������  N_DISP �Xϯ������)CLOCTOL$  QDzC��q�:!�GBOOK ��4d�����r X��/�/�/�/�/�+` =@��9�&	X%��	5��^?{V"_BUFF 2��G z� P]E�? q"�?���?�?OO !ONOEOWO�O{O�O�O �O�O�O�O___J_��P�DCS � Y�d�y�<N?��a��_��_�_�_aTIO 2�m[ ��o5��!o1oCoUoioyo �o�o�o�o�o�o�o	 -AQcu������UER_ITM
�dO�*�<�N� `�r���������̏ޏ ����&�8�J�\�n�p����4'�rSEV��>��vTYP
�����������RS�T��_USCRN__FL 2�
mC���_������ȯگ쯌��/�TP��
��>.-NGNAM7ċ%��UPS_AC�RG���m�DIGI�w�F�m�_LO{AD��G %+��%REQMEN�U�-,MAXUA�LRM��z�.0�2F�
񲒱_Pv�z�� L#1�C���4�/�?�83��P �2�b+ ر6	�:���]  �Z��Ԥ��ϻ���� �X��5� �Y�<�Nߏ� z߳ߞ���������� 1��&�g�R��v�� �������	�����?� *�c�N�����|����� ������;&_ qT������ ��7I,mX �t�����/ !//E/0/i/L/^/�/ �/�/�/�/�/�/??�A?�DBGDEF �<�I�H�J?\0�_LDXDISA�X�*��SMEMO_{APR�E ?+�
 n1)8�?�?��? OO$O6OHO�F�RQ_CFG ��<�r3A *7@i��C*0<I�d%KLзO\On@�<����* P/R **:R*4�O X�O*66_H_u_l_~_ �_�_�_�_-?<�
o�p`�_1ol*o@j,(�_ �o�Tvo�o�o�o�o�o �o1UgN��r�����IS�C 1�+��@ � 3?-���s?C�.?|�g������_MSTR� ���ÅSCD 1��=������ 6�!�Z�E�~�i�{��� ��؟ß��� ��0� V�A�z�e�����¯�� �ѯ���@�+�d� O���s��������Ϳ ��*��N�9�Kτ� oϨϓ��Ϸ����� � &��J�5�n�Yߒ�}� �ߡ߳��������4� �X�C�h��y���������������MK�qA�ҍ�A0�$M�LTARMpB�:�G[� $cl0�����[0METPUܕ0���ډND�SP_ADCOLx��p0��CMNT�� ��FN������FSTLIˀ �Ҏq��A�|���POSCF?=PRPM���	�ST��1�ҋ 4�B#�
"a +	+-?�c u������#/ //Y/;/M/�/y!���SING_CHK�  !$MODAoC��Y�[��%�DEV 	�:	�MC:�,HSI�ZE�=���%TA�SK %�:%$�12345678�9 j?|5�'TRI�G 1�ҋ l [5�O�?Vi�?�?VmL6�YP71Ve�$�#E�M_INF 1���K`)AT?&FV0E0�?uM�)]AE0V1&�A3&B1&D2�&S0&C1S0}=dM)ATZuO�O�DH�O�O�A�?_�HA%_M__q_X_�_�_ [O�_O�O�O�O &o�OJo�_no�o3_�o _o�o�o�o�o�_�_4 �_�_o|�oAo��o ���o��0��T� f���=Oas� ��?��>��b�� �������o���򟥏 ��ɏ:�L���p����� O�Y�ʯ���կ�$� ןH�����1���U� ƿؿ����� �ۿ1��V�=�z��/NITO�RZ G ?;  � 	EXEC�1��2��3��4���5�ȍ0��7��8
��9���D�(��� (���(���(���(��� (���(�
�(��(�"Ҫ(�2/�2;�2G�2�S�2_�2k�2w�2���2��2��3/�3�;�3���!R_GRP_SV 1�JK� (�m��%T1_�D�:>��ION_�DB� ��-�  ��> �&���������'p�N ��,���)-ud�1#59�K�]���PL�_NAME !�[5���!De�fault Pe�rsonalit�y (from �FD)���RMK_ENONLY�/���R2A� 1�L�XLȆ���l d^� %7I[m�� �����!3EWi	�2���� ����//)/;/���e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o�o1oCoUogoyo
�< T/�o�o�o�o�o�o 1CUgy��o"�}
��
�P�� ��'�9�K�]�o��� ������ɏۏ���� �5�G�Y�k�}����� ��şן�����1� C��$�y��������� ӯ���	��-�?�Q��c�u����� F�nH F�� G3=�
�]��ƿؽ

�d\�����+� 9ǫ���d�]�|�gϠ��� �ȿϵ��� �������=ߓ���`�4p�
���	`�ϣ�����߆�:�oA���� ��
� OA�  2��,��� 
�
���0�������  �h  3�=�  GS���Ϫ�� ���������(�S�d�KRR��~�����?� | ����~|� @D�  ��?���{�?\���\��A�Ǐ�K%H� � ;�	l��	 �X8  ���������� �� � � l����K(��K(��K ��J��n�J�^J&	u������Wa��@Y�,@Cz@I�@Ɂ���:I�=�N���f��N����_� a������?�*  �ȯ  �9� H� �� ��\�?s8y��
�/\��x��� �M�!\����:���D
� [ Y��w�so�  ~Ї���H	'� �� �I� ��  �?�F:��È�È=�#�������]���@��F��9/Y�����)/HN�Б/  �'�&t� @2���@���@� @Z� @�C� C��_C��\C� C� �C����@@~1		�	� -� EB 3�?6��K5"�1g5\�Dz��?��?�?�?��?�2�l� í��E1E  �\��55\�p7A?�ffJ�EOWO��? �ЌO�K�18x\��O�J?��7$��C
(\��EP�HI0������Y#?L	 8D��1;�Cd;�p�f<߈<���.<p��<�?��J3��@�Y�������/�?fff�?0?&�PH@��׳R�N�@T싿U[�2�Q��C	 ���_��o�V��vOKo 6oooZo�o~o�o�o�o`�o�o\��UF��  M�oq�_�idt�`xC��E��\�?Gd G;�\� � �9�$�]�H���l� ~�����ۏƉn/�̏ -��N��u�菙���Ƚ�ϟ�����dOA ��!����W�B�{�FB��A|P��;�!kCk�0Яg�U����$����H�3�  �P���R��.40DE� ACx5��B������� �S�B�/�B"�}A��#�A��9@�dZ�?vȴS��~�����<)�+�� =�G��������q���
AC�
=C�������� ��p��Cc�¥��B=���f�f�{S�I����HD-�H��d@I�^�F8�$ D;q�oʭ���Jj��I���G�FP<���x�QpJnP�H�?�I�q�?F.� D�|\8� ���%��I�4�m�X� jߣߎ��߲������ ��3�E�0�i�T��x� ������������/� �S�>�w�b������� ��������=( :s^����� � 9$]H �l������ �#//G/2/k/}/h/ �/�/�/�/�/�/?�/�
?C?.?g?"�('��g�3:n?'Q���5W53�V��?�?�2���?�?�Q4M㇬�?�?�Q�=��O%O4Ue'��T9?M?IOmO�OP�O�O�L�P_RP�N���"_u?._X_C_<|_gY���(�_�_��_�_�_�_�_TAB� �_oFo1ojoUo�o5_`��o�o�o�k/�o��o+;aO��{fgy�������  2 Fn�HTFF��TFG=b�B�0����C9��"`�@��m����T@�E�� F�5��H C፰��ɏQK����E�h�1�a �o�0�B�QK?q�c�T�@TE�dT@T@r�i���
 Q� ��Ɵ؟���� �2� D�V�h�z������l�����;�~Y���$MR_CABL�E 2��H �x�QTP@�@Y�`�������%u��`�C�TAO8�tBx�@���V��`�M�TDO��1��H�>hQ�c�
P�
PCQ�6'�~ȅ�����"��2�1�C�)�HE�ٿ�7��T� Ko�G�YϾ�}��Ϲ� ��������N�I��k߀C�Uߺ�y���1��A ���"�4�TH��c�u�܇�TH*��**} ףOM ������%TBU��-%% 2345?678901����! ����T@�T@\�5T@TA
����not sen�t ��9�W�E�TESTFEC�SALGR  e�gRJ\�d��@�
,��P�PTDl��TG������
 9�UD1:\mai�ntenance�s.xmlY � ���DE�FAULT܌עG�RP 2��� � E�TE  �%�1st mec�hanical �check�TA���d��� �@�1CUgyTB��controller�����"�	//-/?/�cM�g/TB"8}#ʰ�"�/���/�/�/�/�/J*C�-?|/Q?��/?�?�?�?��?�C� ge�.� battery�?A?O�	n?COUO�gOyO�O�9�dui��able�O��p"�C��O'G2O_�_+_=_O_��4g�reas�O�Gf�B�S-�@�Q�_��O@�_�_�_oo�
�4�oiG�_�_�_��_�o�o�o�o�o�X�:�O�F��s<�@q&�
~oSew���Lt�?B�)�;�M�_���Overhaul`/�|��� x�p������ۏ����#��p$̏K�����z� ʏ����ß՟� 6��Z�l�~�4�e�w� ��������ѯ �2�D� �+�=�O�a������ 毆�
�߿���'� v�K�]Ϭ���п�Ϸ� ������<��`�r�G� ��k�}ߏߡ߳���� &�8��\�1�C�U�g� y��ߝ�������"��� 	��-�?���c����� �����������T� )x���_����� ���>Pb I[m��� (�/!/3/E/� �{/�j/��/�/�/ �/?Z//?A?�/e?�/ �?�?�?�?�? ?�?D? V?+Oz?OOaOsO�O�O �?�O
OO�O@O_'_ 9_K_]_�O�_�O�O�_ _�_�_�_o#or_Go �_�_}o�_�o�o�o�o �o8o\onoC�og y����o�"4 F�-�?�Q�c�u�� ���������p)�;���~�	 X=�0j�|���}�B ���� ϟ����)�;�M� _�q���������˯ݯ ���%�7�I�[�m� �������ǿٿ�����!�3�E�WϽ� }�݁?�  @~� ���ϨϺ�~���������~�*�+�** F�@  ������]�c�u߇�I�p�߽��������� ��E���5�G�Y��}� �������q���� �e���U�g�y����� �����������- ?Q������� ���]>���~��$MR_H�IST 2����q� 
 \��$� 2345678�901��?%��9~�����|� :/L/^//'/�/�/�/ o/�/�/ ??�/6?�/ Z?l?#?�?G?�?�?}? �?�?O O�?DO�?hO zO1O�OUO�O�O�O�O��D]SKCFMA�P  ��Rt��X�@ _�UONREL  ��Dq)QVREX_CFENB[W
'S�UtQFNC{_mTJOGOVLIM[Wqdq�PRKEY[W��U�U_PANpZX�R�RRRUN�\��[SFSPDT�YP�XfUSSIG�N[_mTT1MOT��_jQR_CE_�GRP 1���)SyU����o�C�o �o\d�o�o>P t+��a��� ��(�:�!�^���� ��{���o��Տ��ɏ�H���l�#�QQ?Z_EDITXd#W�LcTCOM_CF/G 1�]~U˟�ݟ� 
��_AR�C_xR[e�YT_MN_MODEXf{磚_SPL���VUAP_CPL�T��TNOCHEC�K ?[ �O ����ͯ߯� ��'�9�K�]�o���𓿥���D[NO_WAIT_LWg���`NT���[.��C�	�_ERR�a2	�YV���`�rτ�@��7Q�ϻ��.�O7�}�>�| V�a�d߯A<`S?��K�&��:P��0�PAR�AM8´[� 6RX�ϩ�^�X���� = ������� 1�C��O�y��g�����]��������)�LbODRDSP�S�Zf�XOFFSET_CAR��z�_��DISl�]�S_A�.�ARKXg��OPEN_FILE���Za򑢖
�OPTION_IO�_�Q���M_PRG %�Z%$*.��WmO����g��S_J6R��y 9�y	 ��Hy�J�C�?�RG_DSBL  i�)Q"��<�RIE�NTTOZP�ACY�9P(QA =�UN�/IM_D��&R���?�VC�LCT ��͞�r�d�Ed<j	;_PEX6���n�RAT6� d�U��d�UP �H��R �����!//)�$s�2�c��L�XL�2l{�w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�?�?�?�?�G2e/O O 2ODOVOhOzO�O�O�O^b�?�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏���O �(�:�L�^�p�����@����ʟܟ�$�� � �<�$�P)�f� x���������ү��� ��,�>�P�b�t�C� U�����ο���� (�:�L�^�pςϔϦ� �χ����� ��$�6� H�Z�l�~ߐߢߴ��ߐ�����������!�;�M�w�k�}� b��� � ���������z 
�4�*�<� N�l�r������R ��4���	�	`�x*<��:�o�Zl~���A�S  �	�,��U�����0�����  h��� =�  GS �A�����CU@�yd����C$K O�UN �)���)�HZ$� o| ���� @D�  !?��#�?�"�D�	�"!�E�  �;�	l"	 �X8  ��b!Y  � _� � lx"�~"��H<zH<W��H3k7G��CG���G9|��>/5��/�$��CC  C/� 4�� ��#(!?�#�*�  ��  �9*&0H&0&0�? ?�2?�BY�������^�H�� `?� �?�!�3���*�  �� ��0��0�  �0� F�O��%	'� � �<BI� � � ���&=��!�`OrKC!��  @�(��O��DȕI�O�&NX 
_  �' V�!I0CX C���\CU0CY0C�]?/_A_����@�@�)	�	� ~�- �'B� �VX �U��Q�U$"z�ob?'oo7o�]oHbIAl� í�LB�e}Q�e  E���R�A�!�=p�a?�ff��o�obo ��{Ia�8�-;z?��H�1!�*(�iuPrx`�io!h#h$�C?L�@��dHa;�Cd;��pf<߈<���.<p��<�1?Xz�/�g@��!���"� ?ff�f?�P?&��$@���,��N�@T�8���R�= I`%p�(���vT$�o ď���ӏ���0�� T�f�Q�����s�������[�}��ݟ>�٘C�	 E��:2Gd G;��-���y��� ��֯�������0�� T�?��O��E����ǿ %��a��$�6�H��j�	�oAϚ���@���ϻ��Ͽ&WA�pҰ	7;C��I����?X�?��w�~߷���99�P�:2L1H^>�PDE� C�U�Ļ��Կ�А�4�@I��8=B�/B�"�}A��#A���9@�dZ?�vȅ;���~���<)�+� �=�G��v䀽�q���
AC
�=C���������� ��p��Cc�¥��B=���ff��{8=I����HD-�H�d�@I�^�F8$� D;����̠�Jj��I�G�FP<����QpJnPH��?�I�q�F.� D��|��z� e��������������� @+dO�s ������* N9K�o�� ����/&//J/ 5/n/Y/�/}/�/�/�/ �/�/?�/4??X?C? |?�?y?�?�?�?�?�? �?O	OOTO?OxOcO �O�O�O�O�O�O�O_ _>_)_b_M_�_q_�_м_�_�_��(���33:�_�q��e�U�3�V�oo(b��4oFo��4M��`oro��=���o�o4Ue'��T9�m�i�o�o
(@.|i�P�rPr~������_�����y���(��;�`&�K�q�\���B�t� �������Ώ����0:�(�^�L�/d�n��������ڟȟn�{f ���(��L�:�p�~��  2 FnHn��F�Ж�G=��1B/`��C95Л����@!����
���E��� F����H C���B���o���{�������ÿ��?��ܱpp���������k��o�
 ʿ-�?�Q�c�u� �ϙϫϽ���������ߖ����\k�~�Y��$PARA�M_MENU ?��e� � DEF�PULSE��	�WAITTMOU�T{�RCV�� �SHELL_�WRK.$CUR�_STYLy�κ�OPTС��PT�B����C��R_DECSN��cu6�0� B�T�}�x������� �������,�U�P��SSREL_ID�  �e�q�d�U�SE_PROG �%_�%Q���e�C�CR��v�qg���_HOST !_�#!����T�p���'�� )c��_�TIME��v���~P�GDEBUGt��_�e�GINP_F�LMSK��	TR\��PGA�  ��j��CH��TWYPE\�h�P� J�������� �/9/4/F/X/�/|/ �/�/�/�/�/�/?? ?0?Y?T?f?x?�?�? �?�?�?�?�?O1O�WORD ?	_�
 	PR� ��MAI-�	�3SU��lCTEJ ��-H	��yBCOL���I�O.L�� ��`�����d�T�RACECTL �1��ei� pp�p"_!S�F_DT Q��eMP~PD � bsZ_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�o�o�o �o�o
.@Rd v������� ��*�<�N�`�r��� ������̏ޏ���� &�8�J�\�n������� ��ȟڟ����"�4� F�X�j�|�������į ֯�����0�B�T� f�x���V_����ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~������ � 2DVhz ��������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����߀�����"�4�F�P���$PGTRACE�LEN  Q� � ���Q��f�_UP _����������  ��f�_CFoG ����*P�������������x���  �����DEFSPD� ���O�x���f�H_CONF�IG ���}�� Q�Q�d\��&u� O�_�P����l{�Q��f�IN��?TRL ������8���PEA��K������[���f�LID�����	~��LLB 1�K�_ �|�Bk�sB4;�� |��TN��� <<{��  ?�~ �~����� 3Q7Ik����g/�/ 9/�2/o/b/t/�/���GRP 1� ��Q�A��333�P�A��D�@� D�� D@7 A@O-T`���09"9[�[�� �/v>>´u3W?@;Bx0�1?i?{?�?�?��?�
��?����?0OBN,O =?o=	7LGO�O CO}O�O�O�O�O_O�O�"_�O2_X_C_  Dz}S�_Q�
m_�_]_ �_�_�_o�_,ooPo ;oto_oqo�o�o�o�o��o z!P�
V7�.10beta1��� A��>/qB1��@�!,p�>y�#Cq;3���+q@�
=Sq>waG�+rm8cq>��z�!�!�!;q;t  ������Ap���2k��	�� -����o�5�oI��>l��V���z�ۏ��,p\��"��u0�����N� �F���Pq�!�p�r� B�B�m�_�B�H���Q�Q�L�|�����ǒ
�x˔x7��3������S����` =�_�;�k�\�o�u�_��A�������KNO?W_M  �����SV �K�r���_/�A�S����w�b�t���P�=��M��#�K� �;r	~��	�	� ���ύ��� ���"Pqx{b�g�XcΦ���MR�#�⽀1Ώ�X�5���˱-O�ADBANFWD����ST�!1 15˕��4��;� ;rQ���9�K�]ߎ߁� �ߥ������� ���� V�5�G��k�}����@�����������2%�8�8���<b�6��!�3L�^�p����4 ���������5��(�6EWi{��7�����8`��!�MA��4I��OVL/D  Aϭ/��PARNUM � (����SC-H� �
''�85)�G%UPD���R5�/��_CMP_0ذ�)��'թ$�ER_CHK�%�������&�/�+RqS���ס_MO��(8_?��_RES+_G$��A
��� �?�?�?�?�?�?OO OFO9OjO]O�O�O�Of7K�s<�?�Oh5�� �O�O�Oj3��_0_5_ j3D P_o_t_j3� �_ �_�_j3� �_�_�_j3�=o,o1oj2V 1��+���@k��p+2THR_IN�R������d�fM�ASS�o Z�gM�N�o�cMON_QUEUE �(ը���q��N� U��!N�fx/sEND84qR?NyEXE]Nu�s BE\p>/sOP�TIO;w[;2pPR�OGRAM %�z%1pko/0rT�ASK_I��~O?CFG �/��9�DATA۳�B�"�2������ ̏ޏ�����&�8�J��\����������i�IWNFO۳ц��!t r��!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w�җޔ�҆� �I8�. K�_<��B�����ECNB�Ƚ@��2���G<�2�Ȼ �X,		�!=�{��Oϸ�@��h�$3��!g�gɏd���_EDIT ��B�����5�WERF�L~x�c�RGAD�J ֬�A�  �?X &սa��2q�ñ���??�  Bz�X <g�X ��%S���Ș�M:Ֆ�2�H��	�H)pl�&�bB=P��UT@V����*
�/� *�*:���7�$<��]`A��8���@z�o����iX"R����`�������(��A]`������ �~�(�z�d�^�p��� ����������V R <6H�l��� �.�* � D��z�/�/ ���r//n/X/R/ d/�/�/�/�/�/�/J? �/F?0?*?<?�?`?�? �?�?�?"O�?OOO O�O8O�OtOnO�O�O �O�O�O�O�Of__b_ L_F_X_�_|_�_�_�_�_��	U�_o��Mo�oqd�t$ �o�kto��opo�o8�PREOF �H������
��IORITY��w�ƀ�MPDSaP�q��p�fwUT$�|����ODUCT!������OG��_TG��&��ʥr�HIBIT_DO����{TOENT �1۬� (!?AF_INE�pC�~N�!tcpN�>v�!ude���?!icm��;�֥rXYA�ܬ����)� "��������=� �,�i�P� ��t���ß���Ο�@��A�(�e�w�*�sA��H�p�yߺ�̯�ï>��J �"�/�,쩯�����ܬ�A~j�,  �>p���g�y�������C��Z�ݿ��������ENHANCOE ߘ���A���d�s�Z�  �D�v't�/As����PORT_NUM��s��]u�_�CARTRE��|�ׂSKSTA�w��SLGS@�����j�xpUn?othing{�\� n߀ߐ�B߳��������TEMP ��y��e��_a_?seiban�oK� �o[��l������ ��������G�2�k� V���z����������� ��1U@yd v������ +Q<u`�� �����//;/ &/_/J/�/n/�/�/�/ �/�/?�/%??I?��>�VERSIop�w��0 dis�able��`=SA�VE �z	�2670H844Z8F?�?!c��?�?��O 	<H�ronK	eOtse�O�O�O�O�O�J�LO"_���7]_�p 1���0iP9b�Us_�_�W p/URGE2�B�p	�؁WF�P��tH��v�W<��T{q��WRU�P_DELAY ����wvb_HOT %�u�rb�Vo��UR_NORMA�L5h�rEo�oigSE�MIyo�o�oqQS�KIPQS��bSx D?#@?GYk.}�u ��w������ ��>�P�b�(���t� ����Ώ��ޏ��(� :�L��p�^������� ʟ���ܟ�$�6����F�l�Z��������5�?$RBTIF�Tj~ҠCVTMOU�����ҠDCR�QS�y ��:uCL�CL	��A7�fy8s��F��@���~%��a5.~�A� �;�Cd;�p�f<߈<���.>�]�>П�򐿺�z���� ���,�>�P�b�tπ�ϘϪϼ������eR�DIO_TYPE�  X]Կ��ED�PROT_CFG� �w#�9TB�H�SE6��a2�nH� �ѱB�[� �ߝ�ѿ��u������ �ݞ�<��oc���v� �����������&� 4�R�W�ܥ���n��� ������������"D� Ih�jz��� ���.3R f �x���� �/*//N/�P/ �/t/�/�/�/�/�// ?+?�/L?�/p?^?�? �?�?�?�?�??O4? �?HO6OlOZO�O~O�O��O�O�? O_ޣ8�I�NT 2�8i�р�G;� O_a[��xο�_J�f�0 �_ �[�O�_�O�_�_�_3o !oWo=ogo�o{o�o�o �o�o�o�o/S eK�w���� ���+��O�a�G� ��s�������ߏŏ���'�ĮEFPOS�1 1��  x�Ou�T�|_�� ��Θh�z���� � 9�ԟ]������~��� R�ۯv�����#�5�Я ��}�h���<�ſ`� 鿄��Ϻ�C�޿g� ϋϝ�8�Jτ����� 	ߤ�-���Q���N߇� "߫�F���j����� ����M�8�q���0� ��T��������7� ��[�m���T����� ��t�����!��W ��{�:��p ��A�e  �$��Z�~/ �+/=/��$/�/p/ �/D/�/h/�/�/�/'? �/K?�/o?
?�?�?@? R?�?�?�?O�?5O�? YO�?VO�O*O�ONO�O rO�O_�O�O�OU_@_ y__�_8_�_\_�_�_ �_o�_?o�_couoo "o\o�o�o�o|o�o�)�o&_�cK�2 1�W�M�� ��o��7��4�m� ���,���P�ُt��� ��ҏ3��W��{�� ��:���՟p������ ��A�ܟ� �:����� ��Z��~�����=� دa����� ���D�V� h�����'�¿K�� o�
�lϥ�@���d��� ��߬Ͼ���
�k�V� ��*߳�N���r���� ��1���U���y��&� 8�r���������� ?���<�u����4��� X���|�������;& _����B�� x�%�I�� B���b�� /�/E/�i//�/ (/�/L/^/p/�/?�/ /?�/S?�/w??t?�? H?�?l?�?�?O�?�? �?OsO^O�O2O�OVO �OzO�O_�O9_�O]_��O�_gyt3 1� �._@_z_�_�_o"_ @o�_do�_ao�o5o�o Yo�o}o�o�o�o�o `K��C�g ���&��J��n� 	��-�g�ȏ��쏇� ���4�Ϗ1�j���� )���M�֟q�����ϟ 0��T��x����7� ��үm��������>� ٯ���7�������W� �{�ϟ��:�տ^� ����Ϧ�A�S�eϟ�  ���$߿�H���l�� iߢ�=���a��߅�� �߻����h�S��'� ��K���o���
���.� ��R���v��#�5�o� ����������<�� 9r�1�U� y���8#\� ��?��u� �"/�F/��/?/ �/�/�/_/�/�/?�/ 	?B?�/f??�?%?�?<�_�T4 1�_[? m?�?%OOIOO?mOO �O,O�O�ObO�O�O_ �O3_�O�O�O,_�_x_ �_L_�_p_�_�_�_/o �_So�_woo�o6oHo Zo�o�o�o�o=�o a�o^�2�V� z�����]�H� �����@�ɏd�Ə�� ��#���G��k��� *�d�ş��韄���� 1�̟.�g����&��� J�ӯn�����̯-�� Q��u����4���Ͽ j�󿎿ϲ�;�ֿ� ��4ϕπϹ�T���x� ߜ���7���[���� ߣ�>�P�bߜ����� !��E���i��f�� :���^�������� ���e�P���$���H� ��l�����+��O ��s 2l�� ���9�6o 
�.�R��?�45 1��?��� R/=/v/|�/5/�/Y/ �/�/�/?�/<?�/`? �/??Y?�?�?�?y? O�?&O�?#O\O�?�O O�O?O�OcOuO�O�O "__F_�Oj__�_)_ �_�___�_�_o�_0o �_�_�_)o�ouo�oIo �omo�o�o�o,�oP �ot�3EW� ����:��^�� [���/���S�܏w� � ��������Z�E�~�� ��=�Ɵa�ß���� � ��D�ߟh���'�a� ¯��毁�
���.�ɯ +�d�����#���G�п k�}���ɿ*��N�� r�ϖ�1ϓ���g��� ��߯�8�������1� ��}߶�Q���u��ߙ� ��4���X���|��� ;�M�_��������� B���f��c���7����[����� $6 1�/����j ����b���! �E�i�(: L���/�//� S/�P/�/$/�/H/�/ l/�/�/�/�/�/O?:? s??�?2?�?V?�?�? �?O�?9O�?]O�?
O OVO�O�O�OvO�O�O #_�O _Y_�O}__�_ <_�_`_r_�_�_o
o Co�_goo�o&o�o�o \o�o�o	�o-�o�o �o&�r�F�j ���)��M��q� ���0�B�T����ڏ ���7�ҏ[���X��� ,���P�ٟt������� ����W�B�{����:� ï^����������A� ܯe� ��$�^����� �~�Ϣ�+�ƿ(�a� ���� ϩ�D���h�z� ����'��K���o�
� ��.ߐ���d��߈����5�-7 1� 8����.������� �������N���r� ���1���U�g�y��� ��8��\��� }�Q�u��" ���|g�; �_���/�B/ �f//�/%/7/I/�/ �/�/?�/,?�/P?�/ M?�?!?�?E?�?i?�? �?�?�?�?LO7OpOO �O/O�OSO�O�O�O_ �O6_�OZ_�O__S_ �_�_�_s_�_�_ o�_ oVo�_zoo�o9o�o ]ooo�o�o@�o d�o�#��Y� }��*����#� ��o���C�̏g����� �&���J��n�	��� -�?�Q����ן��� 4�ϟX��U���)��� M�֯q���������� T�?�x����7���[� ������ϵ�>�ٿb�<H�Z�8 1�e�� !�[��������!߼� E���B�{�ߟ�:��� ^��߂ߔߦ���A�,� e� ��$��H���� ~����+���O����� �H�������h����� ��K��o
� .�Rdv�� 5�Y�}z� N�r��/�� �/y/d/�/8/�/\/ �/�/�/?�/??�/c? �/�?"?4?F?�?�?�? O�?)O�?MO�?JO�O O�OBO�OfO�O�O�O �O�OI_4_m__�_,_ �_P_�_�_�_o�_3o �_Wo�_ooPo�o�o �opo�o�o�oS �ow�6�Zl ~���=��a�� �� �����V�ߏz�� ��'�ԏ� ���l� ��@�ɟd�퟈��#� ��G��k����uχ�MASK 1������ӯ᧳�XN�O  ¯��MOTE  ���8�_CFG �?������A��*S�YSTEM*7�V�9.40107 ���7/23/2021 A �q����z�REPOW�ER_T   � $FLAG�r�����STA�RT�� , �ɶ$DSB_SIoGNALr�$ײ?UP_CND��7�?�RS232X���� � $CO�MMENT �$DEVICEwUSE��PEE�$PARITY���OPBITS��F�LOWCONTR�O��TIMEOU�*���CUS�M��A�UXT����INT�ERFAC8�TA�TUZ����CH�� t $OLD_>��C_SW �F�REEFROMS�IZ��n�ARGE�T_DIR �	$UPDT_M�AP�¹�TSK_wENB��EXP��z��!/�FAUL���EV���RV_D�ATA��  �$3�Ep�  � �	$VALUH�� 	/�GRP_ �Ų3�  2� �SC��
�  �$ITP_�E� $NUM�c�OUPr���TO�T_AXZ���DS}P��JOGLI��FINE_PC)�ny�OND��$���UM��K��_MIiR����P6�TN��APL���_EX�'�ԕф�������P=G<�BRKH�� �{NC��IS K� c�TYP��n���P��D8��� �BS�OC��8�N��DU�MMY166��S�V_CODE_O�Pv�SFSPD_�OVRDl�#�L�D����OR��TP �LE��Fd�����OV��SF�RUN���SF5�����oUFRAK�TOiĿLCHDLY��R�ECOV�����WaS��������ROv������_5�  � @��SD�NVE�RT��OFS��CP���FWD����ឦ�ENAB���T�R����_%�FD}O �MB_CM��z B��BL_M��(��-32=�V�����BЋ��G.A�A�M?�! ��o��_�ME ��M��x��T�$CA�е Dj��� HBK�����I�Ov� �IDX�PPA�
�	������DVC_DBG��E ��F�����]��g�]3�e��ATIOr�������UL�иy�AB��۰Y���З��F�h����_����S�UBCPU���S�IN_հW��1�,FWʲm�$HW_C1��"!� K&�F$AT��K��_$UNITw�q >j ATTRI�~"���CYCL��NE�CA��FLTR_2_FI��������LP��CHK�_��SCT�F_�j'F_t,�"�*FS8�Oo"CHA �(p>1Nx�=2RSD��`첇�
��� _Tl�PRO�n�EMP����k�T+2" K��+2F �6DIAG~ �RAILACS�M|�LO�����M7��PS��w� � ���PRGS�� I��AC9+�	��FUNCl���RINS_T����0�<Dm�RAM@��l��� eC���eCWAR���CBLCUR�zH�DA�K�!�H�HD�Au�fA�H�C�ELD@������C��oA�1��CTI	BU��K�$CE_RIA��V��AF	 P�CS,��IUT2�0C��f�@OIu DF_�LEc1����p�LM�QFA��HRDYYO���RG�@H_0����@�UMULS�E�P�'3nB$�J��J����FAN_ALMLV���aWRNeHAR�Dw���$�P��p@2�aS���O�_����A�U��R04��TO_SBR;�e�Ћjj �;DA�cMPINF¹��!�d�A�cRE	G�C�V�����d��DAL_��!�FLL%l�$M�@� ���f� K�%h,uCMf9NF�!�ON �j!e0�b/r8F�3��� ���� ���$Y�r����z�d���$ �4�EG7������q#AR�й��2�3�uܼ@A�AXE��RO�B��RED��WRd��h�_"���SYe���qj�D�SN�WRI���vJ STڰ�Ӆ��i���El!M��t8���ca��B����9\�3� OTO�aM���ARY��̂�1��W���FIJ���$�LINK�QGTH���T_������30���XYZp���"!/�OFF��R���ЀB�Ђ1Bq�������r�F�I� ��������1B��_J)�K������hX`����3F$6��|0�R��Cٰ0�D�U���3�P�3TU�R`XS3�ځ�bX]�� �FL�i��0�pQ�5���34���� 1M�K��M��!�5�5%	B'��ORQ�6��kC蘹��0G�O@�N	B��8���a�OVE��rM����s7��s7��r�6���5���5���4�ANB!�7�IQ�q��� v�fW�/��;����s���[���ER��oA	B�2E��3�	C��A��o ��]E�2؇�A��AAX��K��A�S! �XŹ1d��Qdɋ�c� ��cʹ�c��0cʞ�c���c�1+�cƗP`ɗP pɗP�ɗP�ɗP�ɗP �ɗP�ɗP�ɗP������ɯ �RC�DEBUB#$=AIc�2�����AB�7����V� A" 
��n�q ��F �*� 狡 籡  �� ��1 瞁 缁�OT��IR��r�LAB−�> KGROh� �Bl� B_�1 �z��3���`�����8��va��AND���@����va"� ��Jq��6��AE�� �NqT)`��h�VEL�1 ��r��1z���VP?Rr�#NA`|�-�CS1��%��3񤞂  �S�ERVEh�p	 q$^�i@��!��SPO�BP_�0T �!��򜱱p
�  $TREQ�b
-� �IR2
0'P�0_ � l'@�Q�&ERR���"I� v�N�TOQ����L�Pb�j���0G��%��A��RE�@ G ,��4N ���RA� 2 �d�+�'  �p$+��2yPR�̄pOC�A=  � uCOUN�T�� ��SFZ�N_CFG 4G �f�"TA�?#���ӡ� ��e�s ���M �R�q`����4� �FA6P��DV�X����H�r���� �P?b���HELpj� 5��B_B;ASA�RSR�f%@E�S1Q^ 1��^ 2�*3�*4�*5*�*6�*7�*8�Q!�RO�����NL��q�AB���0_ A�CK��IN#T_�uUX`�Pya9_P�U�Cb*ROU��P�M@�h>#�z`|�>�T�PFWD_KAR���aw RE���PP8��Ab@QUE�i+� ��k�C`VaI`���>#�o3w��f�SE�M��F
��PA�S�TY 4SO�0ldD�I,1�`���1=�wQ_�TM�cMANRQ�]F�ENDjd$�KEYSWITCaHo3�1?A�4HE��BEATM�3PE��pLE��1��HU҃3F�4�2SDDDO/_HOMGPO?a0EF��PRw��/�{�uC�@O�Qt �OOV_MԒ��Ev��OCM ��7
�����?#HK�q DH��g�Uo�2M�px�4W��FORC�c�WAR����?#O}M�p  @��T��u`U��P�p1�V�,p�T3�V4���T�p(O�0L�R���hUNLOJ0m�dED[a  ��SNPZpSk �0pADD���$SIZ�a$V�A���MULTI�P2?c�PA�Q? � $Y9@`HR���rS���C� ��fFRIFY"#S��0�YT�`NF`DODBU]�G��e�c�iX��Fqw@IA���》������_ �p� � ]`�TE�l�񢞃SGLoqT��]�&��s��F�pp�STMTj��sPS�EGn�BW�qtS�HOW�uZ!BAN�pTPT�������+�h�J�1 V�_G�; ��$PC��$��T�FB�QP-�SEP�0A+0/��D�~�� �hA00��p��Pw��P�w��Pw��Pw�5u�6�u�7u�8u�9u�Au�Bu��Pw�|�x��pBw�Fu���9���1���Gp9���1��11�ω1܉1�1��1��1�1�1*�1�7�2t�2��2��2���2��2��22�ω2܉2�2��2��2�2�2*�2�7�3t�3��3��3*��3��3��3��T٨܉3�3��3�U3�3�3*�37�U4t�4��4��4��U4��4��44ωU4܉4�4��4�U4�4�4*�47�U5t�5��5��5��U5��5��55ωU5܉5�5��5�U5�5�5*�57�U6t�6��6��6��U6��6��66ωU6܉6�6��6�U6�6�6*�67�U7t�7��7��7��U7��7��7��7ωU7܉7��7��7�U7�7�7*�77��1VP�@U� ! ��v"
��V��b�� x $gTOR�1%p  ���M	 RJ 1 +�Q_�<R����P�S�D�C�AY�s�_U8�`~�RYSL� �� � ]er{��dRg�@���@��4rVALU{60�6F���=F��ID_L`C�HI
I�R$FI�LE_]36'$$�S�P��SA� h�b E_BL�CK�3o�qxD_CPU�	^`�	R`��9K>`YopW3R � � PW�>� �`�LA�q�S���RUN8pG���@6�6�HW0X��.��T2�1_L}I�R   � �G_O�2�0P_gEDI�R�PT2�x!�i	0��`��`��TABUI����" $�91LgINE�sIAG_�Njp�`��SCޤP# �CL�LS �PT�RY�TB{C2a�$ �fp`{@8p9`�1xFTDH$CTDC8u�c aM�]&s!\'TH�`"�Q�$8�'R�!-`vPERVEC�$Cķ$Hq(!0�  �%X -$�!L�ENC�$C� :0R1A�0+b��W_T�i1�!#2)7MO��(eS�`ERTIA�m�/Q9!�� f;DE<v5�aLACE=RO��CC'co��@_MA�C`u6�5�7�1TCV�<�1�7TiA�:�5�:@M�t3F�E�3F�JP%AB�M@D�@J��_�Rt5aA�5�!2P`�pE�zAs3-`JK�FVK��AOQ�AHq�@�J��A�CJJ�CJJ�CAAL�C�@�C��@�FTq�B5�#
@N�1�<
P�;�0m��_��qp��� CFGb&{ `�GROU��(�qr9�N? C�ceP?REQUIR�"`@�EBU�c�!AF$Tv02%�Q� �V(!�F`.$' \��A�PPR�PCLm�
u$�N�XCLO���YS%�Yt5'"�f( �Mq �0	@RN8d_MG.qB`Ca��c LhA@�0MgBRK�KiNOLDKf�pR�TMOw�j{m<eJ�3P�D�0�C�0�C��0�C�0 S�06�e7��e}q�DR-%)�� �R	2�x(w�A6sPATH2w�KqAsKq8Gs(`�P(q��SCA��g�R6AaIN�"UCU0<1Z�pCO�UM�xY+0T J@�q�!�z�@��z�`�pPAYLO�A�gJ2L��R_	A��L� ����#�LeR_F2LS3HR�$P�LO��q�Q��s_��sACRL�_!1�u���w�tRH���m�$HLb��F�LEX�S�BJ,&* P�R=/O/�/��/V܀�%+ :�/ 6�0Q�h�?Q0�0??0<F1h��� ʗ??Q?c?u?�?�?��E�?�?�?�?�?�?O !O3OѨ�5GLC�Dސ@ �TOfOxOg�JT��ϡX{�HA�E=�%��E ��x��O�O�O�@�E�E �E�E __$_6Y� ܀IT, �8 V_h_z_�� ��AT㖍Q?@E�LQ���XJ�P+v�PJEx`CTR�q�ޑTN�ƅWHA_ND_VBm�ہ��t-�20Lf�$��SWۑ�!)c.� $$M5� 9i6�hab�warܔ�e��b��A �<f�٢EmAVl��hjAvkA��k��Wk� hjDvkDʅkPepGN�ST�jgV�wiV�N�hDY �PLf������ G� h�G�b���G%���r��eP�e�e�e�e�e�e�ur�>�t/ X�=�0r �T�
a�`�ASYMuu����Puv.K��}b��_ W���p�t�m��)������J��`$�pD:	C��_VI���
c� V_UN �� �ȳO�J�E� ��b��y������?@���`����G��0̄Ԅ�0 HR���0"�u�j"DI��`�SO�bvISS1 ذ��I��A�a y�������" DP��w 2 � -:�ME9���4D��T�PT' F�Rp!N�R��	 (�2!&)T( ;Q $DUMMY1�a�$PS_�RF���n$m&2`FLAKPYPw��"#$GLB_T[� ��% ��ڀ �����3 X�P�WqST�DA�PSBR6M�21_V�RT$S/V_ER5�O���#� 3CL� �"AR�Ol�qGL� EWLQ�4 4SP!$Y
ɲZɲWK3�@L�6ӡA��r9�-1U155� C�Ne0- $�GI��}$11 �4*4d0LQ6 qLSP�6��}$F��E�6NEAR3�N��F�90�TANC����JOGܗ��` 7D�$JOINT��J���-1MSETLQ8 E �7E�5��S����4��LQ9� � ��U9�?��PL?OCK_FOa�A�ސBGLV��GL�HTEST_XM��P>AEMP@�R8�B�"j@$U$�02F��25�Pd3�A6�Bh=�o@�A4�!CE8P|�3�@ $KAR��}M�TPDRA40T�1VECy�V@kIU�A7�AHEq@OTOOL��=SV��;REPIS3)�]R96�a�ACH$@�PE8JQO�p#\$3Oq��0SI�R  �@$RAIL_B�OXE��0RO�BO�D?�1HOWWARQ�Qj �QROLMu"�UE��T��Ru��PҐpO_F�v�!0HTML	5��q��" ��>��-0wQq:
O �R
"POC�;Kb��A`�n.0OU&B< 	t0�E4���j@֚bPOsa��PIP�FN1�SR�RwQ���AJ`!�CORDEaDo@{pi`�0XT�`��1)�Pq�O� �= D � OB�ѿ�o@wqV#� �r����SYSqA�DR�q TCH�� > ,C�E�Nz��AvA_�4�ttN�B�pVWVA~�? � P�12�PREV_R�T��$EDIT��vVSHWRv�P�&�p1�E1� D�����tȱ$HECADA	��s�KEE1P CPSP]D �JMP$pL�2ڀR5��@p쁪lvI�@S��C�N�EFP����TICK4��"M���H�J�{HN�!A @p8g�R�(�_GP���V���STYnr�QLO��!�pG���E�B�`
��pGzu%$�q�4=:� S��!$����!�%��&P��S�QUP���"�TE�RC ɱ[�S`�C �0� s�1�rǈ�4Q��O 
#�I�Z�$�1�%i!PR`�`v!Ւc��`PU���_DO�2spXS:"@K�AXI�c�AUR��R����P���2v1я�_4PDrEETE�PxB pz���Fz��A��}��]$9�W2ر	`p0S=R�Dl��[� ��j���}�ҩ������ �������������� ����2�(��V�f�6�C��D�CU���x*�0TSSC� � E h0DS�ŀQ\ SP�2�A	T�Б�摤�s�Y"�ADDRESGSB��pSHIF5b�A_W2CH�.qI� ����TU� Io� �FKbCUSTOTf� qVTBI�GerЌHF�ɓ_�
�J
 ��V�a���H 	\Y��h���̣�Z��C'㦒i��ʛf2���TXSCRE�E	rI��TICNA#3�0dԆ4(18F�F�J�J TY�0 ɒDq1� ���Cr����pRRO���0������nUEO�K# �r�]q{ S$1Dq'RSM���U�`o���uS_^3;�� +�>�Y��F�CdB�ޘ� 2J�UE�F�L�2~�ՐGMTL�!�� �a�A pBBL_�PW�C �M ����OX1��LEv���P�����RIGH��B�RD4l�CKGR�C #�T�`"��WIDTH�S�p��Q�!�GQ �UI`E9Y-`�N d<0"`��P炧PёBAC�K�u"��1�F�O�a��LAB�?�(�I�PhB$U�R�Q����I_�H>�� O 8V�0!_������RE0jB����X����O}��P��� 7�U�GRxB�QLUMG)�f�GERV�aTpo�P�0jv�Q�z�GE��0�1d��b�LP�o�	El���)������qP�	5�6�7�8�j���А�0%��[&qQbASZ�P�n�USR14R �<Y��U�2�Ê2F�O���2PRI��mx�P���TRIP�Qm�UNDON�S�0(��
��Q�	����BC�=� qT��cԑG �aT`居��OS:!�&RI����CQ��U�:?L3S>+"Ǆ�0�BU���V4/F/T�ƅN�OFF�@60W)�%\#O� �@U�`�$Z�$V�`GU>qP�!�B�#��'��SUB�ǂ �E_EXeENpVb��WOۡ� X{ ��WQA�pc&1��b�V_DBE3]0^�c	T- ��Y���1`��sOR�P�5RAU��"�4T�9jws1_�pO��Z | jxOWN|�{t$SRC���c�&�D�@�5��MP�FIބ��E�ESP ᑬ�|�UUv�QrcRp���3�p��[ `} �32{t��J�COP&�!$:��_@��0�A�a�EO2CT5�31AC31OC
��p�R��� \��SHAD�OW&�GS�A_UN�SCA&S�C[��CD�GD|QqEGAC��C����VC�C>t#]� �R=q64�$5PER��J\�H��S� C�`JUDRkIVǖP�_V���mT���PDDMY_UBYCRT
�+#4���I�|��q�XOA�R�P_�@ބ�RL�B�M��$r�DEY�osEX�`�ӒEMUb>�X��=d0�US%�0��_Rz�[�������\�Gw�PACIN��1�RGAvd�b��#�bQ#�bc�AREz�+!�"/S�b�p�^ ��y@G�PP�G��`�p0SR �p_ ~�@ ��d�2	�B��REIcSW�`_A$�a� >cӐOYl�QA~�Es��E��U��d �!��0SHK��`= ]z]���Bp���sEA���w30�0Eu�nuMRCV��a U�� O�M�0CH��	�r�#�c�rREF ���v�v�q4p� s�p h�z-��z-��{O��v��_�0�z���{@�S�15g�S���0R��b �!`��ri�t�U��OU0�N��bL��RS ]�e�2�^��e�'�Ԑ��_`E����f�UL���`F@CO� a/`,�NTACn�OB@m�(y�Py�8�L�S����S��(��P�wVIA26c ����HD����$JO�/���$Z_�UPL���Z�W��ڑ7���_LI�$EP,�#�@��ڑX�_�t_��ِ|DR��d 5E��PAP� E�CACHSLO!������0`��k�@CC0�M%Iw�F/�ѥT�ЦN��$HO�0�2��OCOMMhS�O� ��d�A��@�VP�b+pT�_SI	ZS^�Zp`Y��Z��O16�MP~�FAIj�G�t��AD����BMRE�βc�G�P�%`@�FASY�NBUF�FVRTaD ��c�6�OL��D_�#(�WQ#PC%_�PUc��Qbp��ECCU�hVEM�`��p�ϧVIRCற ����_DE�LA�cA���TAuG�R2aXYZ]�E�2aWq����ă�2��T5PbIM������k ĥGRABBr(!YIcNpLERW`9C!���F_D�PY��5��b֪�c��n���eR@��LAqSx�Yqn�_GEu�Af�A��"���T� A5QG@Q�eI�Կb,�ƀPBG��V��Q�PK�`��v��GI��N��Gr# �Ѡ�$۱��g���Sа��INe��@L"1v�h�B@�3{"PB5�J�I&`��A���@��d�s�_AC���@�"i�o����!P�YJiAD���a�T���j $>1IT��0n��U-C|VsSF|@�3k  ��B[y���UR�vSM�l��8ADJ�0�5eؐZDi�m D��)�AL�Ͱ� �(�PERI^�$�MSG_Q �$d������O2����n�M��1��#���XVR�o���T�_OVR�� �ZABCz5p�bf����
k���ACTV�S:� q � �$����CTIVB�IO�R��fQIT(S�bDV'@#
�av����AM� PS�B ǳ�B����LST`R�̐ �/_S�A���DCS;CH�2r L�1S����@#P��c�G�NA�'5c�R_GFUN����Z� 2Js[�$W$L�R�� �ZMPCFz5ts��hA��QWLNK�"
�M2a~{4u $���p�CMCM~`C��CCzA-!�P� �$JK#E$D I�Q"b"['O@g%O@E'0�p�t`"�'UX���UXEDa�&��V%�%�l%�!�!�)�!�'J F�TFZ�Q#4Yq	�=Z�v ���S ��%1Y1�D:�_ w 8�pR���U�A$HEIGHwcM�?(4�:��΀%0քx � ,G�$B8�_@U�jBSHIF��58R�V0�F����2[ C �F"zAK�-@bb�1 ���C>�DH5CE�hV��$1SPH�ER�P y ,�4�`8v?�9�`�P�Lc`N��˂ J����A�BO�WER �B�A��@�FSM_DRYf>�%�E�B%��A �O�M�B�`��N�JUM<�O�O�OY_�D�����iG�]S�IG�SPD=�}�|X�X��_�ZR��_�F�ې[��C�Q�C��QNGe�z� �:YH_�II_A�IRPU�`  :Z  :oa^r�8���@\k  �@�ISOLC  �lEkb�àla�edR�!k�0o�JOB�!Tf�g�Cjc�@;�Cts#��?�H�haH844  t~��y�@�E����Ox�@S23�2u� 1�E�S� LTE�� ?PENDAN�ps��a�a�|��oB@Mainte�nance CoKns0��0�"*��<�No Use �Z� �~�������ƏD�B�rN��r�a
e��qCHO� ��m�A		I��!�UD1:o��R�SMAV��? e��EaSR  �\kt �A��̐��TVv� e��I���^���V  2dv�Q�� Ds P 	 koo�e�^������E�� §���Я���*�� :�<�N���r�����̿ ���޿ �&��J�8� n�\ϒπϢϤ϶��� �����4�"�X�F�h� ��|߲ߠ��������� 
���T�B�x�f�� ������������� >�,�b�P�r�t����� ��������(8�^L��A�$SA�F_DO_PUL�S�pCq�p�CQsSC�AN� e�F�`S�C�@)��*ШQ�p�p
�a�d�q(Y�Y���� ��4 FXj|���`���/��E�25$�@)d5$�P!���) @��b{/�/�/�/d)x/ �Z��$�_ @�#T`�/?!?3?~@9T D��@? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO��O��v)p�O�O�O�G  
��;�o�DQ�ap��U
�u���Di��J0 � ��j� w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5�G����/p������� ��ʏ܏� �O�#%,� >�P�b�t���������Οӑ��0]RZS(U d]�1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ����Z��%�7�I�[� m�ߑߣߵ� ����� ���!�3�E�W�i�ԟ ��3"��������� ��'�9�K�]�o�}� ��������������  2DVhz�� �����
.`@Rdv��O O3�����// */</N/`/r/�/�/�/�/�/�/�*��/"?.,6��iR?�M�	123456�78ARh!B?!�� ���P�?�?�?�? �?�?�?O"O(A�KO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ |]:O�_�_�_�_�_�_ oo/oAoSoeowo�o �o�o�o~_�_�o +=Oas��� �������o9� K�]�o���������ɏ ۏ����#�5�G�Y� k�*�������şן� ����1�C�U�g�y� �������������	� �-�?�Q�c�u����� ����Ͽ����֯ ;�M�_�qσϕϧϹ� ��������%�7�I� [�m�,ϑߣߵ����� �����!�3�E�W�i�@{���������6�������.�@�\:Cz  B\�_   �M�2�� }��M�
���  	������������
�����Pb t������� (:L^p� ��5��� // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2?Da5:2��K2<]4� S5��  �m;�?q�s�j2|���t  t�h�9�?��(�3 `:2�j2�? Og�s�.�$�SCR_GRP �1*+*�4 � ���� F5	 �^A� fBwBpD�1L3�OG�Gp�O�O�OP������BDE� DP�� }CW�K.A�RC Mate �120iC 67w890��M-VP�A 8��M2I�AZQ�C
123�45[T�FO2  ,x0�� �VfA�F@UA�CUA.\1�AtJ�A�Y	�Roo(o:o�Lo\l��H�f@�TjGUB�o�O�o �o�o�F����oP�o=C8/{hGxxl`-X�IB�c�ƈ�r�t�AAt�  @����u�A@��p� ?��w�rHc���z��AF@ F�` )�1�(U�@�y�d��� ����ӏ����z}�q�r`"���1�C�B�Q� 揗�������ߟʟܟ � �9�$�]�H�����@-�C�O��دF7���կ
���q�q6�����G@�pJ�c��`��W�\�C����A�p��õ�o�e$а.Ĳ�� ���-���B�N�`�/� P��(�Ϥ�@��y��������J_ІT�;��S�5@EC�LVL  ������RѰQ@N�L�_DEFAULT|V�J��P�j�HOTSTR�v�ѱ��MIPOW�ERFU�X���ެ�WFDOw� ���4AERVENT� 1	]�]ѣ� �L!DUM_E�IP���j!?AF_INEv�;�C�!FT�j��1��!�o�� ��}���!RPC_OMAIN�����&���VIS�����r�!OPCU�As���a���!7TP��PU��$��d��
!
PMON_PROXY�'�e��V��$ �f�E�!RDM_'SRV�$�g��G!R�T
%�h��:!
��Mm!�i�)�!RLSY3NC��8u��!ROS���y4�/!
CE��MTCOM/'�k�/j/!	3"CON�Sk/&�lY/�/!>3"WASRC�'��m�/?!3"US�B?%�n�/N?!GSTM��h?#�o=?��?��?��?�=��I�CE_KL ?%��� (%SVCPRG1�?/JE2/O4O@3WO\O@4O�O@5�O�O@6�O�O@7�O�O@HwT?_:L9G_L[D t_A!O�_AIO�_ AqO�_A�OoA�O <oA�OdoA_�oA 9_�oAa_�oFA�_ FA�_,FA�_TFAo |FA*o�FARo�FA zo�FA�o�FA�oD� FA�ol�nA�?�2@ O@����>A �$�� H�3�l�W���{���Ɵ ���՟���2��V� A�h���w�����ԯ�� ����.��R�=�v� a���������п��߿ ��<�'�`�Kτϖ� �Ϻϥ��������&���8�\�G߀��:_D�EV ����MC:��4�����GRP 2��՞�@bx 	�� 
 ,�� ���	���,��P�7� I��m��������� ���(�:�!�^�E��� ���߸�o������� ��6H/lS�w �����  D��9z1��� ����/.//R/ 9/v/�/o/�/�/�/�/ �/?]*?<?#?`?G? �?k?}?�?�?�?�?O O�?8OO\OnOUO�O yO�O�O?�O�O_"_ 	_F_-_j_|_c_�_�_ �_�_�_�_�_ooBo To;oxo�Omo�oeo�o �o�o�o,Pb I�m����� ���:��o^�p�W� ��{��������Տ� ��6�H�/�l�S����� ��Ɵ�����S� �ן D�V�=�z�a������� ԯ����߯�.��R� 9�v���o������� ����*�<�#�`�G� �ϖ�}Ϻϡ������π���8��1�n�u�d �u�	\ߥߐ���`������� �%� �<E�L����^�
� ^�n�|�f������ ����2��Z���D�2� h�V�x�z�������� (���
@.dR t����� ��� <*`��� P�L���// 8/z_/�(/�/�/�/ �/�/�/�/?R/7?v/  ?j?X?�?|?�?�?�? �?*?ON?�?BO0OfO TO�OxO�O�?�O�O�O �O�O_>_,_b_P_�_ �O�_�Ov_�_�_�_�_ o:o(o^o�_�o�_No �o�o�o�o�o�o 6 xo]�o&�~�� ���>d5�t� h�V���z�����ԏ� ��:�ď.���>�d�R� ��v����ӟ���� ��*��:�`�N���Ɵ ���t�ޯ̯��&� �6�\�����¯L��� ��ڿȿ���"�d�I� [��4��|ϲϠ��� ����<�!�`���T�B� d�f�x߮ߜ������ 8���,��P�>�`�b� t����������� (��L�:�\������ ������� ��$ H��o��8�4� ���� bG� zh����� �:/^�R/@/v/ d/�/�/�/�//�/6/ �/*??N?<?r?`?�? �/�?�?�?�?�?�?&O OJO8OnO�?�O�?^O �O�O�O�O�O"__F_ �Om_�O6_�_�_�_�_ �_�_�_o`_Eo�_o xofo�o�o�o�o�o&o Lo\o�oP>tb ����o�"�� �&�L�:�p�^���� ������܏� �"� H�6�l�����ҏ\�Ɵ ���؟����D��� k���4�����¯��� ԯ
�L�1�C������ d����������$�	� H�ҿ<�*�L�N�`ϖ� �Ϻ����� Ϫ��� 8�&�H�J�\ߒ��Ϲ� �ς��������4�"� D���ߑ���j���� �������0�r�W���  �������������� J�/n���bP� t����"F �:(^L�p� ����/ /6/ $/Z/H/~/��/�/n/ �/j/�/?�/2? ?V? �/}?�/F?�?�?�?�? �?
O�?.Op?UO�?O �OvO�O�O�O�O�O_ HO-_lO�O`_N_�_r_ �_�_�__4_oD_�_ 8o&o\oJo�ono�o�_ �o
o�o�o�o4" XF|�o��ol� ���
�0��T�� {��D�����ҏ���� ��,�n�S������ t�����Ο���4�� +���ޟL���p��� ��ʯ��0���$�� 4�6�H�~�l����ɿ ������ ��0�2� D�zϼ����j����� �����
�,߂Ϩ�y� ��R߬ߚ��߾����� �Z�?�~��r��� ��������2��V� ��J�8�n�\�~����� ��
���.���"F 4jXz���� ���B0f ���VxR�� �//>/�e/�./ �/�/�/�/�/�/�/? X/=?|/?p?^?�?�? �?�?�?�?0?OT?�? HO6OlOZO�O~O�O�? O�O,O�O __D_2_ h_V_�_�O�_�O|_�_ x_�_o
o@o.odo�_ �o�_To�o�o�o�o�o <~oc�o,� �������V ;�z�n�\������� ��ڏ���ʏ�Ə 4�j�X���|����ٟ ��������0�f� T���̟���z��ү �����,�b����� ȯR������ο�� �j���aϠ�:ϔς� �Ϧ����� �B�'�f� ��Z���jߐ�~ߴߢ� �����>���2� �V� D�f��z������� ��
���.��R�@�b� �������x����� ��*N��u�> `:����& hM��n�� ����@%/d� X/F/|/j/�/�/�/�/ /�/</�/0??T?B? x?f?�?�/?�??�? O�?,OOPO>OtO�? �O�?dO�O`O�O_�O (__L_�Os_�O<_�_ �_�_�_�_ o�_$of_ Ko�_o~olo�o�o�o �o�o�o>o#bo�oV Dzh���� �����R�@�v� d������ ����� ���N�<�r����� ؏b�̟���ޟ �� �J���q���:����� ȯ���گ��R�x�I� ��"�|�j�����Ŀ�� �*��N�ؿB�ԿR� x�fϜϊ������&� ����>�,�N�t�b� ���Ͽ��ψ������ �:�(�J�p�ߗ��� `��������� �6� x�]�o�&�H�"����� ������P�5t�~���$SERV_M�AIL  ~��t �ZOUTPU}Ti�}@^RV 2��;  w  (D<�^SAVE�x	�TOP10 2>�	 d z�0 BTfx���� ���//,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�?�? O0O$O��YP�[�FZN_CFG ;��w����dAGRP 2�nG� ,B �  A�@~�D;�� B�@�  B�4�RB21��HELLgB���� ��G_&[%RSR&_'_9_ r_]_�_�_�_�_�_�_ �_o�_8o#o\oGo�o��o�n�  ��tb�o�o�o�b�o b��orp��g
�b2�d�l�mOr�F�HK 1�K ������ ��(�#�5�G�p�k��}�������ŏ׏�LOMM �O'��B�FTOV_ENB�i��grOW_R�EG_UIG�\IMIOFWDL����E|�WAIT�D�Hy�B��� h�ܱ��TIMh����۟VAh ��|�_�UNITC���	L]Ca�TRYh���^ MON_AL�IAS ?e�� he/������̯ ڪ�����!�3�ޯW� i�{�����J�ÿտ� ��϶�/�A�S�e�w� "ϛϭϿ���|���� �+�=���a�s߅ߗ� ��T����������� 9�K�]�o��,��� ��������#�5�G� ��k�}�������^��� ������CUg y$������ 	-?Q�u� ���h��// )/�M/_/q/�/./�/ �/�/�/�/�/?%?7? I?[???�?�?�?�? r?�?�?O!O�?2OWO iO{O�O8O�O�O�O�O �O�O_/_A_S_e__ �_�_�_�_�_|_�_o o+o�_Ooaoso�o�o Bo�o�o�o�o�o' 9K]o��� �t���#�5�� Y�k�}�����L�ŏ׏ ������1�C�U�g� y�$�������ӟ~��� 	��-�?��c�u�����������$SMO�N_DEFPRO�G &����ա &�*SYSTEM*�����$SPD_L�ĤRECALL �?}թ ( �}��A�S�e�w����� /���ҿ��������+copy m�c:diocfg�sv.io md�:=>192.1�68.56.1:24292�m����Ϥ�51�frs:�orderfil�.dat vir�t:\temp\@H�Z����߬�-��*.d������p߂���ߧ�xyzrate 11J�\�Q� c����﫲8����?mpbackI��߸w��� }/1�db9�*F�X�a����l���3x1�:\�� ;�������v�������41�a9�K���f��� 	.�@�����u� ���G��b� *�����`�q���� 9K���//&8 �\m//�/��Q/ ��/�/?"4�X i?{?�?��C?�h? �?O�?0/B/�/�?wO �O�O�/IO�/dO�O_ _,?�?�Ob?s_�_�_ �?;_M_�?�_oo(O :O�O^Ooo�o�o�O�O So�O�o�o$_6_�_ Z_k}��_�_E�_ ��� o2oDo�� y�����oK��of��� 	��.�Ώdu��� ���=�O����� *�<�ŏ`�q������� ��U�ޏ���&�8� ˟\�m��������G� ڟ����"�4���Կ i�{ύϠ���M�֯h� ��ߞ�0�ÿT���w� �ߛ߮�?�Q����� �,�>�����s��� �ϼ�W����������$SNPX_A�SG 2����<�� 7 0+�%��d��  ?�-�PAR�AM <�^F� �	R�Pg��+�g����� ��/�OFT_�KB_CFG  �)�B�,�OPIN_SIM  <���#5?/��RVNORDY_�DO  �����QQSTP_DS�B����$�SR� <� � &�����=�/��TOP_ON_E�RR^-�PTN� <�6��A RING_�PRMpVCNT_GP 2<�:��I�x 	���+�~���(�VD>eRP 1�����<�/(/:/L/ ^/�/�/�/�/�/�/�/ �/ ??$?K?H?Z?l? ~?�?�?�?�?�?�?O O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o co`oro�o�o�o�o�o �o�o)&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�{�x����� ����ҟ�����A� >�P�b�t��������� ί����(�:�L� ^�p�������Ϳʿܿ � ��$�6�H�Z�l� �ϐϢϴ���������PRG_COUN�T���6�EN�BK�M;���H�_�UPD 1�T  
��*�ߤ� ����������'�"�4� F�o�j�|������ ��������G�B�T� f��������������� ��,>gbt ������� ?:L^��� �����//$/ 6/_/Z/l/~/�/�/�/ �/�/�/�/?7?2?D? V??z?�?�?�?�?�? �?O
OO.OWOROdO vO�O�O�O�O�O�O�O�_/_*_<_�_IN�FO 1��sfЈP	 __�_�_�_�Y@(���@^.D?���q��_�_oo�=oEd D���URD�  C4 � ´Pobm�YS�DEBUG Ё���VPdiّ`SP_PwASS �B?�k�LOG }V.��  VPEh\_�  �e�VQU�D1:\�dc^�b_MPC�m��Qc���q� ��1vSAV �i/�1a�alr�uxSV({�TEM_TIME� 1�g�� �0VP��t	��&}T�MEMBK  ��e��`�oe�w����X|f�� @��TSЩ�Ώތ��d����a 1k@�G�Y�k�}�0o�� ��şן���TSxc� +�=�O�a�s�����������eů���� � 2�D�V�h�z������� ¿Կ���
��.�@��uSK<�A�+�P���X�ϤϘ�=VP"C���b�A����� �� &�8�h�zߌ߀���VQ� �����������5��ʀB�g�y�����VP$����˯�� ��1�C�U�g�y��� ������������	�-?QE�T1SV�GUNSPD�e �'�e�t 2MO�DE_LIM � �y�bp2} ��!�moABUI_EDIT "���SCRN #��m�SK_OP�TION�`D��a��_DI�`ENB�  �ţe>BC�2_GRP 2$�cţc���Qx`C���hBCCFG 3&m�| ���`�$o!//1/ W/B/{/f/�/�/�/�/ �/�/�/??A?,?e? P?�?t?�?�?�?�?�?�O�?+OOOOaOiD LL{OMO�O�O;O�O�O �O__>_�~^_F�3P f_�_z_�_�_�_�_�_ �_o
ooRo@ovodo �o�o�o�o�o�o�o <*`Npr� ��x�@����"� �F�4�V�|�j����� ď���֏���0�� @�B�T���x�����ҟ ������,��P�>� t�b������������ ���.�@�^�p���  �������ܿʿ �� $��H�6�l�Zϐ�~� �Ϣϴ��������2�  �V�D�fߌ�z߰ߞ� ���������
��R� @�v�,��������� `�����<�*�`�r� ��R�������������  J8n\� ������� 4"XFhj|� ����� //0/B/ �f/T/v/�/�/�/�/ �/�/?�/,??P?>? `?b?t?�?�?�?�?�? �?OO&OLO:OpO^O �O�O�O�O�O�O�O_  _6_�N_`_~_�_�_  _�_�_�_�_�_ o2o DoohoVo�ozo�o�o �o�o�o
�o.R @vd����� ����(�*�<�r� `���L_����ޏ��� ��&��6�\�J����� ��r�ȟ���ڟ���  �"�4�j�X���|��� ��֯į����0�� T�B�x�f�������ҿ ������� �>�P�b� ࿆�tϖϼϪ���������$TBCSG_GRP 2'����  ���� 
 ?�  )�;�%�_�I߃� m�߹ߣ������	��)�d � |��?��	 HC꽀��>���:��[ff��C�L��!�8X�d�.�33��C�%�L�d�f�0�&�^&�>���F�\L��Ȭ���BL���B$��9���(���L�8^�p���  @���� ��������0M�*x��?333�~�	V3.�00!�	m2ia�	*� �� ���� ��(���z	 &�'   nB �\n�J2	�*���~CFG ,���� Ц�r�<��� !//*��//U/@/y/d/ �/�/�/�/�/�/�/? ???*?c?N?�?r?�? �?�?�?�?O�?)OO MO8OJO�OnO�O�O�O �O!�;��O�O_�O?_ *_O_u_`_�_�_�_�_ �_�_oo�_;o&o_o Jooo�o���Ϻo���o �o�o8&\J �n������ �"��2�4�F�|�j� ����ď���֏��� �B�0�f�x�8ϐ��� L��ҟ���,�� P�>�`�������h��� ��ί��(�:�L�^� ���p���������ʿ  ��$��H�6�l�Z� |Ϣϐ��ϴ������ ��� �2�h�Vߌ�z� �ߞ�������
ﴟ"� 4�F���v�d���� ��������*�<�N� �r�`����������� ���� &J8n \������� �4"XFh� |������
/ //T/B/x/f/�/�/ X��/�/�/�/??>? ,?b?P?r?t?�?�?�? �?�?�?OO:O(O^O pO�O�ONO�O�O�O�O �O_ _6_$_Z_H_~_ l_�_�_�_�_�_�_�_  ooDo2oTozoho�o �o�o�o�o�o�o�o
 @�/Xj|&�� �����*��N� `�r���B�����̏�� ܏��&����\�J� ��n�����ȟ��؟�� �"��F�4�j�X�z� |���į���֯��� 0��@�f�T���x��� ��ҿ俎��ϔʿ P�>�t�bϘφϨ��� ����������L�:� p�^ߔߦ߸��߄��� ���� ��H�6�l�Z� ��~���������� ��2� �V�D�f�h�z� ������������
 ,R@v�"Ϡ� \���<* `N����x� ���/8/J/\/n/ (/�/�/�/�/�/�/�/ �/�/4?"?X?F?|?j? �?�?�?�?�?�?�?O OBO0OROTOfO�O�O �O�O�O�O__�2_ D_V_ _�_t_�_�_�_ �_�_o�_(o:oLo^o�o�opo�o�o�o�n s �`�c �f��b�$TBJO�P_GRP 2-��e� / ?��f	 r's�/.|��`X?8  �rrDt�  � � �� l�r�c @��`?r	 �C�} �vf  C�w?q�rL���v�q�q��u�qz��q>��=�ZC��p�p��p��?C�  BȺw��"��~�@w�v�X�3�33T��x�p=�7�LC�f��Z�D0�p	����C��pŅ�A��r>�33����s��y<�҉C�\�t��pC�CHȞ�?�
�LR�ԁD��qڌ��x�t��x@p<_X��B$�s@�q �����ßF�X�ڌ�\��� �����~�p?�ffC����[�ޟ�r�����g��Ҩ���@Y�@pB� ֣߯񯔝4��"�� >�H�y�T�f������� οؿ	����(�B�,�P^�hϙ�,���f����u	V3.00�Esm2iaDt�*��Dt�a���� �E�'E�i��FT�F"w�qF>��FZ�� Fv�RF�~�MF��F����F��=F����F�ъF���3F���F��{G
G�dG�G#�
�D��E�'
EMKE����E�ɑE��ۘE��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF��u�<#�
<Kt�����0��oT�����f��?���v�}ESTPA�RS���h9psHR�O�ABLE 10*.y���d*��Q hP��*�*�*��g�a*�	*�
*��*���a*�*�8*���i�RDIq�8q���������J�OR�d�n���������j�SP�6s �w� ������ +=Oas��� ��}O S7r��) ��	-��������!�3�j��NUM [ �e8q�p��` ����j�_CFG 1�+�#�q�@ pIMEBF_�TTU�%6sb�6V�ER�� !563R� 12y� 8$���b�`�1 �`/  z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O_�O�O =__*_@_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o5"8�FXj|�J�b1_��!L6@V5L�MI__CHAN+7 V5} �sDBGLVu��-5V5K��pETHERAD ?Y�O������h�xz�D��pROUTI0!��!��̏��?SNMASKD�V3>U�255.
������,���L�OOL�OFS_DIU���u.�ORQCTRL 3i;���ߪ�T��Ο�����(� :�L�^�p��������� ʯܯ�����!��E��I�PE_DETA�I"�o�PGL_C�ONFIG 9��)�!��/ce�ll/$CID$/grp1I���ѿ���Ͻ󀕏2�D� V�h�zό�ϰ����� ����
ߙ�.�@�R�d� v߈��)߾������� ���<�N�`�r�� ��%���������� ���J�\�n�������.}9�������" 4�!6�\;�8�� �����2�! 3EWi���� �����///A/ S/e/w//�/�/�/�/ �/�/�/?+?=?O?a? s?�??�?�?�?�?�? O�?'O9OKO]OoO�O O�O�O�O�O�O�O_ �O5_G_Y_k_}_�__ �_�_�_�_�_o�_1o�CoUogoyo�o�o����User V�iew ��}}1�234567890�o�o�o(0tX�p��P���i2�i -o������K]�b3u:�L�^�p� �������c~4)��  ��$�6�H���i�c~5ݏ����Ɵ؟���[��c~6��V�h�z�@�������ѯc~7E� 
��.�@�R�d�ï��c~8����п������w�9�?� l�Camera �j��~ϐϢϴ�������Eq���&��o@��R�d�v߈ߚߐ�   X�tym������ �2� D���h�z���߰��� ������
�1��X�(� ��V�h�z�������W� ������C�.@R dv�/�܉�� ��
��@Rd �������� /���{0/B/T/f/x/ �/1�/�/�//�/? ?,?>?P?�Y�D��/ �?�?�?�?�?�?�/O *O<O�?`OrO�O�O�O �Oa?/���QO__*_ <_N_`_O�_�_�_�O �_�_�_oo&o�O/� ���_ro�o�o�o�o�o s_�o_o8J\ n��9oKg9� ��	��-��o>�c� u�������Ϗ�����	Z�0��@�R� d�v�����A���П� ����*�<�N�`�� �_�a����˯ݯ� ����7�I�[���� ������ǿٿ��Z��� p�%�7�I�[�m��&� �ϵ���������!� 3�E��&�9��ϑߣ� �������ߒ��!�3� ~�W�i�{����X� jեH����!�3�E� W���{����������� ������j�+�� i{����j�� �V/ASew �0j�}; ��� ////�S/e/w/���/�/�/�/�/�/�  �$?6?H?Z? l?~?�?�?�?�?�?�;   �/? O2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�o�o�o�o�o�o�&8J\�<  }
�(  �0( 	 l�� ������� ��2�h�V���z���vz
J �D/���� �/=�O�a�s������ ���ӟ�,�	��-� ?�Q�c���������� ϯ����)�p�M� _�q���������˿ݿ �6�H�%�7�Iϐ�m� ϑϣϵ�������� �V�3�E�W�i�{ߍ� �ϱ���������� /�A�S�߬߉��� ����������+�r� O�a�s���������� ����8�'9��] o������� �X5GYk} ������/ /1/C/U/�y/�/�/ ��/�/�/�/	??b/ t/Q?c?u?�/�?�?�? �?�?�?:?O)O;O�? _OqO�O�O�O�O O�O �O_HO%_7_I_[_m_8_�O��@ �R�_��_�_�S�W�p���)frh:\tp�gl\robot�s\m20ia\�arc_mate�_1`c.xml �_6oHoZolo~o�o�o0�o�o�o�h���o	 -?Qcu�� ����o���)� ;�M�_�q��������� ˏ�܏��%�7�I� [�m��������ǟޏ ؟���!�3�E�W�i� {�������ïڟԯ�� ��/�A�S�e�w��� ������֯п���� +�=�O�a�sυϗϩ� ��ҿ������'�9� K�]�o߁ߓߥ߷���:�X!Q �_�P�<< �P ?�������&�T�:� \��p�������� ����>�$�V�t�Z��l������F�@(��$TPGL_OUTPUT <�A��A��  ��#5GYk} ������� 1CUgy������Є��2345678901� ��
//./6#�B� ]/o/�/�/�/�/O/�/@�/�/?#?5?�*}?? g?y?�?�?�?G?Y?�? �?	OO-O?O�?MOuO �O�O�O�OUO�O�O_ _)_;_�O�Oq_�_�_ �_�_�_c_�_oo%o 7oIo�_Woo�o�o�o �o_oqo�o!3E W�oe����� m���/�A�S�� ���������я�{� ��+�=�O�a���o��������͟ߟw��� $$��'� �G�9�k�]������� ��ׯɯ�����C� 5�g�Y���}�����ӿ@ſ�����?�}�рY�k�}Ϗϡϳ���@��������� ( 	 A�/��S�A� w�eߛ߉߫߭߿��� ����=�+�a�O�q� ��������������'�]�K�����  <<4� ���� ������% 7���hz�� ����V�.� dvP��
� �|�/*//N/`/ �H/�/�/B/�/�/�/ �/?r/�/J?\?�/d? �?l?~?�?�?8?�?O �?�?FO O2O|O�O�? �O�O^O�O�O_�O0_ B_�O*_x_�_$_�_�_ �_�_�_T_�_,o>o�_ botoNo`o�ooo�o �o�o�o(^p �ot�@���� �$���Z��F��� ��|�Ə؏6���� � ��D�V�0�b������ ԟn�ܟ
����@� R���v���"�t�����������)WG?L1.XML��;���$TPOFF_�LIM ��������I�N_S]VQ�  ��c��P_MON =���e�����2�E�STRTCHK' >��c�V�L��VTCOMPAT�x��g�VWVAR� ?��%�|� Kٿ =������M�_DEFPR�OG %ǹ%�Tϛ�J�_DISP�LAYX�Ǿm�IN�ST_MSK  �� ��INU�SER����LCK����QUICKM�EN%߯�SCRE�D����tpsc���_�d�c��u�_y�ST��c�R�ACE_CFG �@��%���	�F�
?���HNL� 2A|�u���,�  R��*�<�N�`�r��������ITEM �2B� �%$�12345678�90����  =<����-�5�  !;�C�O����F��� �������C���g�y� B��]��m�	 -GQ�u!G Y�}��) ��/q/��� =/�/��/�/%/�/I/ [/$?/??�/c?u?�/ �?�/O?�?3?�?W?O )O;O�?GO�?�?�?aO O�O�O�OSO_wO�O �O_7_�O�_�__�_ +_=_oa_!o�_EoWo �_mo�_�_�oo�o9o �o�o�o�o�o�o�o C�o���5�Y k}��M�s���� ����1����g�'� 9���E���ӏ������ �۟�Q��u�ǟP� ��k�ϟ{�������� ;�M�_�ٯ��/�U�g� ˯���������I� 	���'ϣ���~�ٿ ��������3���W�iϔ2߾�S��C��7�ψ  ��7� 8�ю߅�
 ���������f�UD1:�\����I�R_G�RP 1D��?� 	 @��=� O�9�o�]�����������������<:�%�?�  U�g� Q���u����������� ����)M;q_0����	����G�SCB 2ES� @�=Oa�s�����=�U�TORIAL �FS���/B�V_C�ONFIG G�S��ы���w/'-OUTPUT HS�h ���/�/�/ �/�/?!?3?E?W?i? {?�?�?e!�/�?�?�? �?O!O3OEOWOiO{O �O�O�?�O�O�O�O_ _/_A_S_e_w_�_�_ �O�_�_�_�_oo+o =oOoaoso�o�o�o�_ �o�o�o'9K ]o����o�� ���#�5�G�Y�k� }������ŏ׏��� ��1�C�U�g�y��� ������ӟ���	�� -�?�Q�c�u������� ��ϯ����)�;� M�_�q���������˿ ݿ���%�7�I�[� m�ϑϣϵ�Q/c%�/ ����)�;�M�_�q� �ߕߧ߹��߾���� �%�7�I�[�m��� ������������!� 3�E�W�i�{������� ��������/A Sew����� ���+=Oa s������� //'/9/K/]/o/�/ �/�/�/�/�/��/? #?5?G?Y?k?}?�?�? �?�?�?�/�?OO1O COUOgOyO�O�O�O�O �O�?�O	__-_?_Q_ c_u_�_�_�_�_�_�_ �Ooo)o;oMo_oqo��o�o�o�o�o�o������o�a�o 9��]o���� �����#�5��_ Y�k�}�������ŏ׏ �����1�C�T�g� y���������ӟ��� 	��-�?�P�c�u��� ������ϯ���� )�;�L�_�q������� ��˿ݿ���%�7� I�Z�m�ϑϣϵ��� �������!�3�E�V� i�{ߍߟ߱������� ����/�A�R�e�w� ������������ �+�=�O�`�s����� ����������' 9K\�o���� ����#5G�V�$TX_SCREEN 1Iu��`�}�V�������Ev�4/F/X/j/ |/�///�/�/�/�/ ??�/B?�/f?x?�? �?�?�?7?�?[?OO ,O>OPObO�?�?�O�O �O�O�O�OiO_�O:_ L_^_p_�_�__�_/_ �_�_ oo$o6o�_�_ lo~o�o�o�o�o=o�o ao 2DVh�o���$UALRM_MSG ?v�� �Y
�� ��%��I�<�N�l��r�����Ǐ��돟uS�EV  �}���rECFG �Kv�  �Y@�  AM� �  B�Y
  �`v��������ȟ ڟ����"�4�B�)��GRP 2L3�; 0Y	 j�����pI_BBL_N�OTE M3�T��l`�{b?���DEF�PRO�p%�{ (%ߏ�b ��-�� Q�<�u�`�������Ͽ຿�޿ϕ�FKE�YDATA 1N<vv�p B�Y @�{ύ�ʠj����Ϡ�,("���Y ��"�	�F�-�j�|�c� �߇����߽������ 0��T�;�x��q�� ����������,�[���<�c�u������� ��`Q�����
. @��dv���� M��*<N �r�����[ �//&/8/J/�n/ �/�/�/�/�/�/i/�/ ?"?4?F?X?�/|?�? �?�?�?�?e?�?OO 0OBOTOfO�?�O�O�O �O�O�OsO__,_>_ P_b_�O�_�_�_�_�_ �_�_�_o(o:oLo^o poG��o�o�o�o�o�o �_$6HZl~ �������  �2�D�V�h�z�	��� ��ԏ���
���.� @�R�d�v�������� П������*�<�N� `�r�����%���̯ޯ �����8�J�\�n� ����!���ȿڿ��� �"ϱ�F�X�j�|ώ� ��/����������� ��B�T�f�xߊߜ߮�څd����`����������#�5��,!�f����q� ������������ >�%�b�t�[������ ����������:L 3pW���o�� � $3�HZl ~���C��� / /2/�V/h/z/�/ �/�/?/�/�/�/
?? .?@?�/d?v?�?�?�? �?M?�?�?OO*O<O �?`OrO�O�O�O�O�O [O�O__&_8_J_�O n_�_�_�_�_�_W_�_ �_o"o4oFoXo�_|o �o�o�o�o�oeo�o 0BT�ox�� �������,� >�P�b�i�������� Ώ��򏁏�(�:�L� ^�p���������ʟܟ �}��$�6�H�Z�l� ~������Ưد��� �� �2�D�V�h�z�	� ����¿Կ���
ϙ� .�@�R�d�vψ�Ϭ� ��������ߕ�*�<� N�`�r߄ߖ�%ߺ��� �������8�J�\� n���!������������"��p$��>�p���M�_� q�I������,��� �����0T; x�q����� �,>%bI� m�����// �:/L/^/p/�/�/�� �/�/�/�/ ??$?�/ H?Z?l?~?�?�?1?�? �?�?�?O O�?DOVO hOzO�O�O�O?O�O�O �O
__._�OR_d_v_ �_�_�_;_�_�_�_o o*o<o�_`oro�o�o �o�oIo�o�o& 8�o\n���� �W���"�4�F� �j�|�������ďS� �����0�B�T�+/ x���������ҟُ�� ��,�>�P�b�񟆯 ������ί�o��� (�:�L�^������� ��ʿܿ�}��$�6� H�Z�l����Ϣϴ��� ����y�� �2�D�V� h�z�	ߞ߰������� �߇��.�@�R�d�v� ����������� ��*�<�N�`�r���� ������������&�8J\n��i����i���������,/F�jQ�� ������// B/T/;/x/_/�/�/�/ �/�/�/�/?,??P? 7?t?�?e��?�?�?�? �?O(O:OLO^OpO �O�O#O�O�O�O�O _ _�O6_H_Z_l_~_�_ _�_�_�_�_�_o o �_DoVohozo�o�o-o �o�o�o�o
�o@ Rdv���;� ����*��N�`� r�������7�̏ޏ�� ��&�8�Ǐ\�n��� ������E�ڟ���� "�4�ßX�j�|����� ��į�?�����0� B�I�f�x��������� ҿa�����,�>�P� ߿tφϘϪϼ���]� ����(�:�L�^��� �ߔߦ߸�����k� � �$�6�H�Z���~�� ���������y�� � 2�D�V�h�������� ������u�
.@ Rdv���� ���*<N` r�������/٠+�٠���-/?/Q-)/s/�/_&,q?�/i?�/ �/�/?�/4??X?j? Q?�?u?�?�?�?�?�? OOOBO)OfOMO�O �O�O�O�O�O�Oկ_ ,_>_P_b_t_��_�_ �_�_�_�_o�_(o:o Lo^opo�oo�o�o�o �o�o �o$6HZ l~����� ���2�D�V�h�z� �����ԏ���
� ���@�R�d�v����� )���П������� <�N�`�r�������7� ̯ޯ���&���J� \�n�������3�ȿڿ ����"�4�_X�j� |ώϠϲϹ������� ��0�B���f�xߊ� �߮���O������� ,�>���b�t���� ����]�����(�:� L���p����������� Y��� $6HZ ��~�����g � 2DV�z ������u
/ /./@/R/d/��/�/ �/�/�/�/q/??*?�<?N?`?r?I�t;}�I�����?@�?�=�?�?�?�6,�O &O�OJO1OnO�OgO�O �O�O�O�O�O�O"_4_ _X_?_|_�_u_�_�_ �_�_�_o�_0ooTo foEϊo�o�o�o�o�o �/,>Pbt ������� �(�:�L�^�p���� ����ʏ܏� ���$� 6�H�Z�l�~������ Ɵ؟����� �2�D� V�h�z������¯ԯ ���
���.�@�R�d� v��������п��� �ϧ�<�N�`�rτ� ��%Ϻ��������� ��8�J�\�n߀ߒߤ� {o���������"�)� F�X�j�|����A� ��������0���T� f�x�������=����� ��,>��bt ����K�� (:�^p�� ���Y� //$/ 6/H/�l/~/�/�/�/ �/U/�/�/? ?2?D? V?�/z?�?�?�?�?�? c?�?
OO.O@ORO�? vO�O�O�O�O�O�O����K������__1]	_S_e_?V,Qo�_Io�_�_�_ �_�_o�_8oJo1ono Uo�o�o�o�o�o�o�o �o"	F-j|c ��������� 0�B�T�cOx������� ��ҏ�s���,�>� P�b�񏆟������Ο ��o���(�:�L�^� p���������ʯܯ� }��$�6�H�Z�l��� ������ƿؿ�����  �2�D�V�h�z�	Ϟ� ���������χ��.� @�R�d�v߈�߬߾� ��������*�<�N� `�r��������� �����8�J�\�n� ��������������� "��FXj|� �/���� �BTfx��� =���//,/� P/b/t/�/�/�/9/�/ �/�/??(?:?�/^? p?�?�?�?�?G?�?�?  OO$O6O�?ZOlO~O �O�O�O�OUO�O�O_  _2_D_�Oh_z_�_�_ �_�_Q_�_�_
oo.oh@oRo)�Tk�)����}o�o�myo�o�o�f,�� *N`G�k� �������8� �\�n�U���y����� ڏ�ӏ���4�F�%� j�|�������ğ�_� ����0�B�T��x� ��������үa���� �,�>�P�߯t����� ����ο�o���(� :�L�^��ϔϦϸ� ����k� ��$�6�H� Z�l��ϐߢߴ����� ��y�� �2�D�V�h� �ߌ����������� ���.�@�R�d�v�� �������������� *<N`r�[�� ����	&8 J\n��!�� ���/�4/F/X/ j/|/�//�/�/�/�/ �/??�/B?T?f?x? �?�?+?�?�?�?�?O O�?>OPObOtO�O�O �O9O�O�O�O__(_ �OL_^_p_�_�_�_5_ �_�_�_ oo$o6o�_ Zolo~o�o�o�oCo�o �o�o 2�oVh@z����� �{��� ��������3�E��, 1�v�)�������Џ�� �ۏ�*��N�5�r� ��k�����̟ޟş� �&��J�\�C���g� �����گ����"� 4�CX�j�|������� ĿS������0�B� ѿf�xϊϜϮ���O� ������,�>�P��� t߆ߘߪ߼���]��� ��(�:�L���p�� ��������k� �� $�6�H�Z���~����� ������g��� 2 DVh������ ��u
.@R d������� �˯/*/</N/`/r/ y�/�/�/�/�/�/? �/&?8?J?\?n?�?? �?�?�?�?�?�?�?"O 4OFOXOjO|O�OO�O �O�O�O�O_�O0_B_ T_f_x_�__�_�_�_ �_�_oo�_>oPobo to�o�o'o�o�o�o�o �o:L^p� ��5��� �� $��H�Z�l�~����� 1�Ə؏���� �2���$UI_INU�SER  ����S���  3�7�_M�ENHIST 1�OS�  �( `����(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1r����	����9 ����936ҟg� y�����,���Ưد� ��� ���D�V�h�z� ����-�¿Կ���
� ϫ�@�R�d�vψϚ� ��;���������*� ��N�`�r߄ߖߨ߸��Gѧ�G������� ,�>�A�b�t���� ��K�������(�:� ����p����������� Y��� $6H�� l~����Ug � 2DV�z ���������
/ /./@/R/d/g�/�/ �/�/�/�/q/??*? <?N?`?r??�?�?�? �?�?�??O&O8OJO \OnO�?�O�O�O�O�O �O�O�O"_4_F_X_j_ |__�_�_�_�_�_�_ ��0oBoTofoxo�o �_�o�o�o�o�o�o ,>Pbt��' �������:� L�^�p�����#���ʏ ܏� ��$���H�Z� l�~�����1�Ɵ؟� ��� �ooV�h�z� ��������ԯ���
� �.���ϯd�v����� ����M������*� <�˿`�rτϖϨϺ� I�[�����&�8�J� ��n߀ߒߤ߶���W߀�����"�4�F�1����$UI_PAN�EDATA 1Q����|�  	�}X������������� ) ���;���J�\�n��� ��������������� "	F-j|c�������4�� C�2�7I[ m���(��� �/!/3/E/�i/P/ �/t/�/�/�/�/�/? ??A?(?e?w?^?�?�6~���?�?O O&O8O�?\O��O�O �O�O�O�OAO�O_�O 4__X_j_Q_�_u_�_ �_�_�_�_o�_0oBo �?�?xo�o�o�o�o�o %o�oiO,>Pb t��o����� ��(��L�^�E��� i�������܏Ooao� $�6�H�Z�l������� Ɵ؟���� ��� D�+�h�z�a�����¯ ԯ����߯�.��R� 9�v��������п� ����k�<ϯ�`�r� �ϖϨϺ�!������� ���8�J�1�n�Uߒ� y߶��߯������"� ����X�j�|���� ���I�����0�B� T�f����q������� ������,>%b I���/�A�� (:L�p� ������ /g $//H/Z/A/~/e/�/ �/�/�/�/�/?�/2?0?V?��}�g?�? �?�?�?�?�?)�?O �OKO]OoO�O�O�O O�O�O�O�O�O#_
_ G_._k_}_d_�_�_�_��_�_�_����$�UI_POSTY�PE  �� 	 o�^o-bQUICKM_EN  <kKo�ao/`RESTOR�E 1R�  ��_B��o�c�o�m ,>Pbt�� ������(�:� L��oY�k�}����ʏ ܏� ���$�6�H�Z� l�~�!�����Ɵ؟� ����	����V�h�z� ����A�¯ԯ���
� ��.�@�R�d�v�!�+� �����˿����*� <�߿`�rτϖϨ�K� �������߿�!�3� E߷πߒߤ߶���k� �����"�4�F���j��|����lgSCR�E|`?�m�u1sc�`u2���3��4��5��6���7��8����TAT8m� �c�%j�USER������TL����ks���4��U5��6��7��8���-`NDO_CFG� S<kw0v1-`P�D0�j���Noneoba�_I�NFO 2T� �`0%��/� ^A��w�� ���$HZ�=~elOFFS�ET W<i �S��`[����/ 2/)/;/h/_/q/�u/ �/�/�/�/�/?.?%?�7?I?�+�o�=�?�?
�?�?L���WOR/K X�?�?�O+O�`�UFRAME  �5�����RTOL_ABRqT|O��BENB�O~�HGRP 1Y�i��aCz  A� �C�A���O__'_9_ K_]_o[�F{`U�H��~�KMSK  �5��KNyA%	��%e?o�E_EVNĜ@�T��f��2Z�
 h��U�EV�@!td:�\event_u�ser\o``C7�eo�?U�F�=Y`SP�^acgspotw�eld�m!C6 �o�o�o���T!�_to 2gw�Q VD� �z���)��� �q����@�R���ݏ ̏������I�8�m� �*���N�ǟٟ����@���3�ޟ�5fW@32[k��18.����� ��ί௻��� �:�L�'�p���]��� ����ܿ�ɿ�$����H�Z�5�kϐϢ��$�VARS_CON�FI��\� FPvS����CMR�B;2b��YU��	��B%1: �SC130EF2� *.�2�S䙒(���P�5U���?U�P@PpsPȣ�' OO����L耱����������mUA�U��U�h B���p� ht��ߕ��߹���� �����%��"�[��� <���|�����z��������IA DcM��,�		d1DeFTG��P �g �8R�TSYNC� �Di�HazWINU�RL ?�
Ђ���'�SIONTMO�U o �?=b�dS۳�S۵�P�A FR:}\A\DATA�  �� M�C�LOG�  � UD1�EX��(�' B@ ����~�/��6/| � n6  �������VO'��  =���͌!&�� �>�TRAIN�T"4�"rd�#p�%�(D��4�d��eDk (���),=��,? 6?H?Z?l?�?�?�?�?��?�?�?�?O O9_�GEhfDk�`(��
�@(��B\G��REkg�Iұ�L�EXgDh���1-�e/VMPHASOE  De�l����RTD_FIL�TER 2iDk �O��}�G_Y_k_ }_�_�_�_�_�_�_� 2_o)o;oMo_oqo�o�o�o�o6SHIF�TMENU 1j^;
 <),%)/R���oT+ =�as���� ���>��'�t�K��	LIVE/S�NA��%vsf�liv�N����A � U����menu��ď^�#�5�Ad�ehk��hMOhml�N�z��ZDT��m�O(�<� }@�$�WAITDINE�NDL�h���OK�  �؜J�S��ڙTIML��2�GğT��w���W�%�W�D�ؘRELE�A��d���GY��_ACT����)ؘ�_� n!	�%�7�����;�RDIS�����$XVR��Ao�N�$ZA�BC��1p�� 	,� ��2��1��@�VSPT q�M\�!$
"�"��a��nτ�#�DCS�CH�@r!E�۲I-P��s���� ��2�D��MPCF_OG 1t�ɶ0��X����R�MP�u���!p�����߲��`  �!$?b���#!D�� D����H���	� �-��Q�>�{�����
�f���C4  ´!�3� �w�k�e� w�������_�q��#"A6��$ٴe��@v���8_CYLIND�Qwm� �&? ,(  *���!#�����  0B�e�� p����/J +/��a/H/�/l/���/�/03xES� Ă�?(<K�Q?@<?u?��?�?�ǖ�1�A��ZSPHER/E 2yj�/�? o/�?1OOUO�/�?�O �O/�O`OFO�O�O_ _tOQ_c_�O�O�__ �_�_�_�_:_o)o;o6ݰZZ%� �d�