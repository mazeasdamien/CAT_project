��   ��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����CCPTP_�CFG_T  �L h$DAT�A_PATH �!$OUTPU�T>5$PART�_NAMEC $�EDGE\!$C�LR_VDB_BUF  $x�_SIZ 9V�ER�DEV_I�D�H �VIS_�RES���P_D�T�POS_OF�S_ENB�TA�R_D� �CHK�_f �DEBUG�_MOD` � MAX_FC_PN���&CUV)S�EG)LAPTPP_� XfH�f�As� L�WAIT_TM �$ABV_PT�H���RETRsEA� �CNS� ��JUMP_LE�N_�$CURQV)f�T'T)�MAd	'ABOV�E_��$TO�L_WPR_CH�X_!b EXP%S�AT 2�ERR_H���-��q�(�q_PROXE N�ON� OPqCF%_S R��$RW�$�DI��$LI�D?EACT_F/3�5XID6�6J8 e9LOC6 ȧ5�P��ANs0�$X5!A���4�_C'CO��5F�IR��0H�SQ�� Xh_#f['�E`H@!p��$N_� 9L�!�ACH:I��L� �DYN_CO SW�;H�Xp�!�: �ALL�
�EP�TH@�
�D�F�NU��C��A8� �FBASFH@&�XYZWSH@�I��010Z�SPUS I@�FZI#U�oV�H#oGAIN�FXYCQ��F�P�Y�P�5n� R6�MI
 EC���Xk,S� �0NGI1�+c22f�L1a�'cIa?a� S .`_C   `b|Iaib ��&|:1 L �38N3�6�TOTx`�8�c��AVG!�$$�FINI�j2�G ��iF�jV�F�6�Q��3��dU�D� ~`
�&sENT�~`$ #yz�b��#�vaf`� mk�q``bST� � ? 
����$s ASS ? ����q���Z��Z�p� SIO�N�x  �XK�qIRTU�AL��q'2 �Z�!FR:\) �\����5UD1:_������q����q!������� ���� �� N��u0o  �&� d����&���1�  @@�@�E�?��BH<H�W��  >g�^�a�d���^�ʂ*����Ĉ��ğ��BȠϟ���f�^�A��D�z������ԛ��?�c�F�s�r�F�K�j�Q,"�Z���2����8������ ��ϯ��󯲯�)�;�M�  ;�:�`I�P�����
�ſ����߽� �"�4�F��j�|ώ����1234?567890���� ������������0� B�T�f�xߊߜ�