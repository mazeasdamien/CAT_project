��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1�TU4QQ���AR�x1R� � /$TIT91� �� � �Td�T0�ThP�TU5�V6�V7�V8�V9�W0�W�WOQ�U�W�gQ�U�W1�W1�W1��W1�W2�R�SBoN_CF�!@$<!J� ; ;2�1�_CMNT�$�FLAGS]�C�HEK"$�b_O�PTJB � ELL�SETUP � `@HO8@9 P�R�1%�c#�aREPR�hu0D+�@���b{uHM9 MN�B;16 UTOB�J U�0 }49DEVIC�STI/@�� �@b3�4pB�d�"VAL��#ISP_UNI�tp_DOcv7�yFR_F�@|%u13���A0s�C_WAx�t,q�zOFF_T@]N�DEL�Lw0pdq�1�Vr?^q��#S?�o`Q"U��t#*�QTB��bMyO� �E � �[M�����RE�V�BIL���!X�I� v�R  �!D�`��$NOc`M�|����ɂ/#ǆ� �ԅ��ނ�@Ded �p E RD_E���h�$FSSB�6�`KBD_SEV�uAG� G�2Q"!_��2b�� V!�k5�p`(��C�00q_ED|� � � t2d�$!S�p-D%$� ��#�B�ʀ_�OK1��0] P_C�� ʑ0t��U �`LACI�!�a�Y�� ��qCOMM� # $D
� ��@���J_�\R BIGALL;OW� (Ku2:-B�@VAR���!|�AB   �BL�@� � ,K�q��r�`S�p�@M_O]�˥��CCFS'_UT��0 "�A�Cp'��+pXG��b�0� 4� IMCM ��#S�p�9���i �_�"t\b���M�1 h$�IMPEE_F�s���s��� t����D_(�����D��F��� �_����0 aT@L��L�DI�xs@G�� �P�$I�'�����CFed XF@GRU@��Mb��NFLI�\Ì@U�IRE�i42� SgWITn$`0_N�`�S 2CF�0M�' �#u�D��!���v`����`J�tV��[ E��.p�`��>�ELBOF� � շ�p`0���3����� F�2T��A`��rq1J1��z _To!��p��g����G� �r0WARNM�p#tC�v`�ø�` � COR-�UrFLTR��TR�AT9 T%p� $ACCVq��� ��r$ORI�_&��RT��S<��HG*�0I���TW��A��I'�T���H9K�� �2028�a1��HDR�2��2�2J; S���3���4��5��6��7
��8��9��׀
 �2� @� TRQB�$vf��'�1�<�c_U<�G� COec  <� P�b�t�x53>B_�LLEC��}!~�MULTI�4��"u�Q;2�CHI�LD��;1ذO�@T�� "'�STY 92	r��=��)2��������ec# |@r056$J ђ��`����uTO���E^	EXTt����2��22"����$`@D	�`&��p������(p�"��`% �ak�����s�����A&'�E�Au��Mw��9 �% ��TR>�� ' L@�U#9 ���At�$J�OB����P��}IG��( dp��� ���^'#j�~�L��pOR�) tf$�FL�
RNG%Q@�TBAΰ �v&r� *`1t(��0 �x!�0«+P�p�%4��*��͐U��q�!�;2MJ�_R��>�C<QJ�8&<J D`5CF9���x"�@J���P_p�7p+ \�@RO"pF�0��I9T�s�0NOM��>Ҡ�4s�2�� @U<PPTgў�P8,|Pn�ć0�P�9�͗ RA����l�?C�� �
$�TͰtMD3�0TD��pU�`�΀+AYHlr>�T1�JE�1 \�J���PQ��\Q��hQ�CYNT�P��PD'BGD̰�0-���PU6$$Po�|�u��AX����TAI�sBUF,�O!�A�1�. ����F�`PIV|�-@PvWMuX�M�Y�@�VFvWSI�MQSTO�q$7KEE�SPA��  @?B�B>C�B�2��/�`=��MARG�u2��FACq�>�SLEW*1!0����
�4ذs�CW$0'����pJB�Ї�qDE�Cj�e��s�V%w1 Ħ�CHNR�;MPs�$G_@�g�D�_�@s��1_FP�5�@TC�fFӓC@�Й���qC��+�VK��*��"*�JRx���SoEGFR$`IOh!v�0STN�LIN>�csPVZ�z�Ц@�D2����r 2��hr�r��1��3` + ^?���եq�`��q|`������t��|aSI!Z#�!� �T�_@%�I��qRS�*s���2y{�Ip{�pTpLpF�@�`��CRC����CCTѲ�Ipڈ�a8���bL�MIN��aP1순���D<iC �C/���!uc�OP4�n �j�EVj���F��_
!uF��N����|a�֔=h?KNLA�C=2�AVSCA�@�A�WQ�a�4�  cSF�$�;�Ir�Kঠ'��05��	 D-Oo%g��,,m�����ޟ��RC�6� n���sυ��U��R�0HANC���$LG��ɑDQ�$t�NDɖ��AR۰N��aqg��ѫ�X��ME��^�Y�[PS�RAg�X�AZ�П���:rEOB�FCT��A���`�2t!Sh`0ADI��O��y�s"y�n!@�������~#C�G3�t!��BMPmt@�Y8�3�afAES$���v��W_;�BAS#?XYZWPR��*��m!��	y�U�87/  ƀI@d��2�8\�p_C:T����#��_L
 � 9K ���C�/�(z�J�LB�$�3�xD��5�FORC��b�_AV;�MOM$*�q�SaԫBP`Ր� y�HBP�ɀE�F�����AYLOAD&$�ER�t&3�2�X�rp�!ҁ�QR_FD��� : T`IH�Y3��E�&��Ct���MS�PU
$0(kpD��9 �b��;�B�	EVId�y
�!_IDXY�$���B@X�X�<&�SY5� � �HOPe�<��AL�ARM��2W�r}rR9_�0= hb P�nq�`M\qJ@$PiL`A&�M#�$�` ��� 8�	���V�]�0�U�qU�PM{�U���>�TITu�b
%�![q�BZ_;�.��? �B pQk���6NO_HEADE^az��}ѯ��`� �����dF�ق�tc`����@�@��uCIGRTR�`��ڈL���D�CB@4�RJ�� 1�[Q���A�2>�&��OR�r��O����T`UN_OO�Ҁ�$����T������I�VaCnp�DBP�XWOY���B��$SKADR��DB]T�TRL��C���րfpbDs��~�DIJj4 _�DQ}���PL�qwbWA���WcD�A��A�=�2�UMMY�9��10�VIȾ ����D;[QPR�� 
M�Z���gE O�Y1$�a{$8��L)�F!/��
����0G�G/��9�PC�1H�f/3#PENEA@T�f�I�/���RE�COR`"JH y@ �E$L�#F$#PR���+jp���nq�_D$�qPROSS]�
���R�r�` >u�$TRIG96�PAUS73ltETgURN72�MR:�eU 0Ł0EW$�~�SIGNALA��QR$LA�З5�1�G$PD�H$PDİ�AI�0�A�C�4�C��DO�D�2�!��6GO_AWA�Y2MOZq�Z��,CS��CSCB�g�K Իa#���E+RI�0Nn�T�`$�����FCBPL�@QBGAGE���P��ED`|BD�wA[CD�OF�q�[F0�FoC��MPM�AB0XoC�$FRCIN��2Dk��@��O$NE�@�FD�L8�� L� �����=��Rw�_��P>� OVR10����lҠ�$ESC_|�`uDSBIO��p��pTe�E�VIB�� `s��Z��V��p�SSW��$�VLY�:�Lk��X���ѣ�0bQ����USC�P��qA=�	Q��MP1%e@&S*`�(bt`'c5۳ESUd��-cWg&S Wg?cWd����Wd��Wd<.���AUTO$�Ya҃�ac�SB����-d���&SwB[��GB�f_$VOLT�g ���  �GAOD!��q���@:�ORQ�ҀKra�$DH_THE&0�Rgp� <qtnwALPHnt��o��w0 Vp]�$�.�Ra�[��s�5�`r�CQ�#BUD�S� F1M���sV
��;��L�b�tk���BRTHR��L��T`�Z���Vɖ��D)E  �1��2�⋅ ��������kѯ�a� �Tt0V�ꆸ������@̈Я�-�"�N~���sS2����INHB��ILTG0ɡ�T?� �3$�w��E��PqQxQ��TqPe��0Y�AF}�O�ນ��ڗ ��qPڳē����bPܙ���PL?���3���TMOU��ēS��� � ��s�/�S18���O��Aܙ��I����CDqIƑ˩o�STI��գ�O:ҋ�,0���AN��Qg�S��+r�#x$�����w�1_����PRA�P`�vC����MCN�eQe�����VER�S��r�oPIw�F�PåǲШ۷G.�DEN��G>�����F�2H�Ƿ�M�7�F��_�MN�D̠,���@�d�{ƭa����OB����U˱z���DI ���#���3�����A��w�Fx���3�O�N�5��Q��VAL��CR[�_SIZp��b�;Qn�REQ�R�b��]2b���CH q�΂�ڃ�Ռ�����:�n�S_U��X��wW�FLG���wU$CV�iMGP�QδFLXP�923R�u�L��EAL�P-�C	�F+rT��W��� �R��c���NDMS�7� ��K>S�P_M'0h�STWv������AL�P���Q����U���U�IAG@,�o��d�U�-�T"	A-`� ���A��� ��H`��Q`��6��Pq_D&��1s��.�P��F�"2�T�� ?7 1A>���#�#L��?`_=i @@>LD�pc�F�0�FRI�0 `Ѐ��1}Ѳ�IV\1�*�^1�U�P`��a��C�L!W��
`L=S&-c&&S�C.w��  L���!����d�Q$w!�҇��$w��p��
�P�5RSM��P���V0h � r�l�d^2AW�a_TRp�}�8@NS_PE�A����< ��$�SAVG�8�6G]%���CAR �`�!�$���"CRa���$ d�#qE�@��"STD���!Fpo��'QOF0��%��"RC���&RC۠�(F�2A�R#7����%, gMA�Q_�a��
QQ��al2��%u4Ib�r7I�R�9�wQ�7�8M/��!C:pR�  �p�2F<�SDN�a0 � W2QM P $Mi��s$cA �$C�cm�9���4���AT�0CY_ �N LS!IG1@x'yB��y@@H2Y��NO����SDE�VI�@ O@�$�RBT:VSP0�3�CuT�DBY|�A�	W`3CHNDGD�AP H@GRP�HE iXL�U��VSЌFx2� DL1p aQ6ROp��FB�\]�FEN�@��S���ChAR d�@DyOd�PMCSb���P薇P�R��HOT�SWz42�DMpEL�E�1/ex\8`�RS T�@���r� hf��`OL�GHA�Fk�Fs�����C�A@�T � $MD�LUb 2S@�E ���q�6�q	0�i�c�e
�cJ��	uݢ�#~X5t+w�PTO��� x�byU DSLAVS�� U  ��INAP �	V�ЊyA_;�wENUAV $R��PC_�q�2 1bLp�wpp B�pSHO+� W ���A�a�qB�2�r�v�u�v�b�_CF� X�` ,f��r�OG� gE��%D�h��p2C�Iߣi�MA��D��x AY?�W� p�N3TV	�D�VE�0@�SKI��T�`g?Ň2�� JZs�! �Cꆻ��f�_SV</ �`XCLU��H����ONL��'�Y��T��OT:eHI_�V,11 APPLY���HI4`;�U�_M�L�� $VR�FY8�	�U�M{IGOC_I���J 1/d��߃O�@X�LSw"�`@$DUMMY�4���ڑ�Cd L_TP���kC��^1CNFf���E��@HT�y� D_#UQ_��ݥ�YPCP��=�� ������uJ �ҟ Y +�
0R�T_;P��uNO�CCb Z�r�TAE���=�פ�DG��@[ D�P_B�Ae`kc�!I��_��H�t~T��E \�pyAb=cARGI�!�$���`[��SGNA] ��`U���IGN�Տ��� ���V������ANNUN��&�˳�EU�<J'�ATCH���J��B��u^ <`@g�����:c$Va������ᑴaE�F] I�� _ �@@FͲITb�	$TOTi �C�O��c� @EM�@NIF�a`tB��c��ùA>���DAY@CLOAD�D\�n���� �EF7�X�I�Ra��K���O�%��a�ADJ_)R�!@b��>�H2��"[�
 c�%��`a�͠MPI�J��D��qA��?�Ac 0� �х�� ��Z�ϡ��Ui ��CTRLܖ Yp d��TR�A8 ?3IDLE_�PW  �Ѡ��Q��V��GV_���`c ��o�;Q@e� �1$��6`<cTAC�-3��P�LQ�Z�Rdz\ A-u:ɰSW;�A\���/Jղ�`b�K�OH�(OsPP; �#IRO� ��"BRK��#AB  �������� _ ���F���`d͠, j@�S�RQDW��MS��P6X�'z��IF�ECAL�� 10^tN��V��豊�V�(0}f�CP
��Nr� Yb�0FLA_#f�OVL ��HE��>�"SUPPO��ޑ�\�L�p��&2XT�$Y-
Z-
W-
���/��0GR�XZl�q�$Y2�CO�PJ�SA�X2R��*r�!���:��"�rI�0)��f `�@CACH�E��c��0�s0L}AZ SUFFI, C��q\��哹6��QMSW�g� 8�KEYIM[AG#TM�@S���n
2j�r���ROC�VIE��~�h ��aBGL����`�?G� 	Q���i��m!`STπ!� �����n����/EMAI�`N��`A��`Z�FAU� �jH�"�qa��U�3�qq� }�k< �$I#�US�� �IT'�BUF`�r�DNB���SUBu$��DC_���J"��"SAV�%�"k�������';��P�$�UOR	D��UP_u �%��8OTT��_B`��8@�LMl�F4��C7AX�@Cv���Xu 	��#_uG��
 @YN_��R�l6���D�E��UM����T��F���caC�DI`BED%T)@C��~�m�rI��G�!c�&��l`���-�P��FZP n (�pSV� )d\��ρ���2ΰ��o�� ����>"$3C_R�IK��kB���hD{pRfgE.(AD�SP~KBP�`�II�M�#�C�Aa�A��UЂG���iCM! IP`��KC��� �DTH� ȷS�B*�T��CHS�3�CBSC��� ���V�dYVSP�#[T_D^rcCONV�Grc�[T� �Fu F�ቐd0�C�0j1��SC5�e�]CMER;dAFBgCMP;c@ETBc� p\FU D�Ui ��+�~�CAD�I%P702#@O��B�qWӏ�SQ��QǀSU��MSS�1ju�4`��TB�Aa��A�1r�� "�Й��4�$ZO@s���l�U�6�&��eP���eCN�c�l��l�l�iGRO�U�W)��S c�MN�kNu�eNu�eNpR|b|�i�cH�pi��z
 �0CYC���s�w�c���zDEL�_D��RO�a���qVf���v{�O�2���1���t��:R�ua�.#�� ���AL� �1s@ˢI1¡�J0�PB��,렒�ER^�T�Gbt ,!@��5��aGzI1LcR1s 
�0&ԠNO��1u����H�����P����Cڠ	�����!���J0��0vH *	�L U�1#J�Q��V
�[�7A z���z��z�n�z�Ѩz�Fz�7w�8w�9Pw���y���1��1��U1��1��1Ě1њU1ޚ1�2��2�����2��2��2��2�Ě2њ2ޚ2�3J��3��3����3��U3��3Ě3њ3ޚ�3�4���EXTF��1w6�.(�0�f�0��U�0ŷ�e.�FD�R5�xTU V�E��?1���SR��R�E�F���OVM�~C)�A2�TROVf2�DT� R�MXa��IN2���Q�2�IN	Dp�r�
���0�0�0�Gu1��[�G`��{�D_�[�RIV�P��oGEAR~AIOr�	K"N�0�y�p��5`@�a�Z_MC�M� ���F��U�R�Ryǀ��!?3 ��p?nЋ�?n�ER�v�Gme��!�P��zIj:�PXqB�RI0%�>`�#ETUP2_� { ���#TDPR�%TBp�������K�"BAC�2| QT��"�4)�:%	`t^B��p�IFI���� Mc���.�PT|��I �FLUI��} � ��K UR�c!���B�1SPx NE�EMP�p�2$��]S^�?x��Jق�0
3VRT���0x/$SHO��Lq�6 ASScP=1��PӴBG_�������FORC�3" �i�d~)"F%UY�1�2\�2
A�h� p� |��N�AV�a��������S!"��$VI�SI��#�SCM4S�E����:0E�V�O���$���M����$��I��@��FMR2��� �5`�r�@ �� �2�I�9 F�"��_���LIMI�T_1�dC_LM�������DGCLFl����DY�LD����5������F  ���D u	 T�sFS0Ed� P���QC�0$EX_QhQ1i0�P�aQ53�5��GoQ��g� ����RSW�%�ON�PX�EBUG���'�GRBp�@U��SBK)qO1L� ��POY 
)�(�P��M��OXta`KSM��E�"�0�����`_E � x
@F���TERMZ%9�c%�aORI�1_ Y�c%d�SMepO��B_ �|&.�`�(�c%��e:�UP>� ?�� -���b����q#� ���G<�*� ELTO��p�0�PFIrc�1Y���P�$�$�$UFR�$��1L0e&� OTY7�PT4q��k3NST�pPATz�q4PTHJ�a�`EG`*C�p1AR�T� !5� y2$2R�EL�:)ASHFTPR1�1�8_��R�P�c�& � $�'@�@� ��s�1 @I�0�U�R G�PAY�LO�@�qDYN_�k���.b�1|��'PERV��RA��H��g7��p�2�J�E-�J�R�C���ASYMFgLTR�1WJ*7����E�ӱ1�I��aUT�pbA�5�F�5aP�PlC�Q1FOR�p�M��GRI!����W��/&�0F0�a H��Ed� �m2N���5`OC1!?�$OP����c��c���bRE�P�R.3�1a�F��3e���R�5e�X�1(�e$PWR��_���@�R_�S�4��et$3U�D��.�Q72 ����$H'�!�`AWDDR�fHL!G�2(�a�a�aT��R��U�w� H��SSC����e-��e���e��S�EE��HSCD���� $���P_"�_ B!rP����}T!HTTP_���HU�� (�OB�J��b(�$�fL�Ex3pWq�� �� ���ะ_��T�?#�rS�P��z�KRN�LgHIT܇5��P ���P�r������PL���PSS<�ҴJQUERY_FLA 1��qB_WEBSOC���HW�1U����`6PINCP	U���Oh��q�����d���d���� �I�HMI_ED� T� �RH�?$��FAV� d�Ł��wOLN
� 8��yR�@$SLiR�$INPUT_�($
`��P�� �؁SLA� ����5�1��C���B��IO6pF_AuS7��$L%�}w%�A��\b.1��0���T@HYķ������Qh�UOP4� `y�ґ�f�¤�������`PCC
`���#���aIP_M�E�񵁗 Xy�I�P�`�U�_NET�9���Rĳs�)��DSP(�Op=��BG�����M��A��� lp:CTiAjB�pAF TI�`-U��Y ޥ�0PSݦBUY IDI�rF ���P�q�� �y0��,����Ҥ�N�Q�Y R��IRCA|�i� � ěym0�CY�`EA������񘼀�CC����R�0�A�7QDAY_<���NTVA�����$��5 ���SCA�d@��CL���� ���𵁛8�Y��2,e�o�N_�PCP�q��ⱶ��,�N�����
�xr���:p�N� �2��Ы�(ᵁ�p���xr۠LABy1���Y ��UNIR��Ë ITY듭��e�ւR#�5���R�_URL���$AL0 EN��ҭ� �;�T��T_U��A�BKY_z��2DI�SԐ�kSJg�����P�$���E��g�R���З A�/���J����FLs��7 Ȁ|���
�UJR� ���F{0G��E7��J7 O^ R$J8I�7�H�R�d�7��E�8{��H�APHIQ�S��DeJ7J8�B��L_KE*� � �K��LM�[� � <X�X�Rl�u���WATCH_VA��o@D�tvOFIELc��cy��L��4� � o1Vx@��-�CT[�9�m�� ��LGH���� $��LG_SIZ�t�z�2y�p�y�FD��Ix���+!�� w�\ ����v��S��� 2��p�������\ ��h�A�0_gCM]3NzU
RFQ\v�v�d(u�"B ��2�p����I��+ �\ ��fv�RS���0  ��ZIPDUƣp�L)N=��ސ�p��z6���f�>sD�PL�MCDAUiEA`Fp���TuGH�R�.OGBOO�a��� C��I�IaT+���`��RE����SCR� �s��D�I��SF0�`RGIO"$D�����T("$�t|�S�s{�W$|��X��JGM^'MN3CH;�|�FN��a&1K�'uЅ)UF�(1@n�(FWD�(HL�)STP�*V�(%Г(,��(RS9HIP�+��C[T�# R��&p:'^9U=q�$9'�H%C�d���"Gw)�0PO�7��*��#W}$���)E]X��TUI�%I�� �Ï���rCO#C� N*�$S��	)���B@�NOFAN1A|��Q
�AI|�t:��EDCS��c�CT�c�BO�HO�GS����B�HS�H(IGN������!O���DDEV<7LL�ѩ�|��­Ц(�;�T��$��2�p������#A
���(�`�{�Y���POS1�U2�U3��Q	��2�@�Ш ��{�PtD�����&q)��0�d��VST�ӐR�Y��B@ ` _�$E.fC.k��p<p=fPf���4�ѩ LRТ� ��x�c �p��<�Fp�d��?"�/_ �����Kqx&���c �MC7�� ���CLD�PӐ��TRQLI0#ѽ�ytFL��,r��5s8�D�5wS�LqD5ut5uORG���91HrCRESERAV���t���t���c~�� � 	u095t5u��PTp���	xq�t�vRCLMC�������q�q�M��k�������$DEBUGMA�S��ް��?U8$T�@��Ee�g���MF�RQՔ� � �j�HRS_RU�7��a��A��k5FgREQ� �$/@x�OVER��n�t�V#�P�!EFI�%�a��g��d���tǯ \R�ԁd�$9U�P��?A��SPS�P��	߃C���͢a��U\�l��?( 	�MI;SC� d@�QkRQ��	��TB �� Ȗ0A՘AX����ؗ�EXCE�SjҔЪ�M��\���W����ԝ���SC>�P � H��̔�_��Ƙǰ]���
�MKHԳK�J� �m�B_K�FLIC��dB�QUIREG3MO��O˫3���ML�`MGմ @�`��T���a#NDU�]��>���k�G�Df��INAsUT���RSM>�a��@N�r]3-��p�5�PSTL\�� �4X�LOC�VRI�%��UEXɶANG�uBu�R�ODA��ŷ�������MF O����Y�b@�e4Ŝ2k�SUP�e��F�X��IGG� � �A��c���c Q6�dD�%�b|�!`�Ȁ!`��|��3w�ZWa�T!I��p�a M��[��� t��MD��I��)֟@���H8ݰM��DIA��ӂ��W,!�wQ�1�D��)��O���]��[ 0�CU��VPА�p���!_V��ѻ� ��P�S�X�5�	�����P��0N��ЍP��KES2���-�$B� ����ND2x����2_TX�d�XTRA�C?�/��qM�|q�`�Pv�`�XҰ�Pt SBq`^�USWCS��T��<	���PULS��A��NSޔ��R��JOIN��H��~`j�=��b��b�����P�=��$��b$���TA����S���S�HS�ME��SCF�aPJ���R��PLQ� 
M��LO��н.�L��^����8��Ҹ����0�RR2���O 1��eA�q/ d$��Iΐ+��G�A2+/� ;�PRIN�w<$R SW0"��a/�ABC�D_�J%�¡u��_J3:�
�1SPܠe�u�P��3��р`
u��J/���r�q�O8QIF��CSKAP"z{�{�J���QL2LBҰ�_AZ�r�~ELxQ��OCMP���T���RT�����c1�+���P1��t>@�Z�SMG0���=�JG�`SCL<�͵SPH_�@���%V�u� RT�ER`  �< A_�@G1"�A�@c���\$DI�
"23U�DF�}!LWn�(VELqIN�b)@� _BL�@u��$ G�q�$�'�'�%`<��� ECHZR/�TS�A_`����E�}`<����5�Bu�Ht1}`_�� �)5 D2d%��A4I��N9t&FR�DH�A���ÀP�$V `�#>Aa$��Ͳ�$Q���R}ӆ��H? �$BELvᵆ><!_ACCE�!c�x�7/��0IRC_] ���pNTT��S'$PS�rL�d� /Es��F{�@F
��9gGCgG36B���_�Q�2�@�A���17_MGăDD�A]"ͲFW�`���3�EC��2�HDE�KPPA�BN>G��SPEE �B�Q%_pB�QY�Y�|�11$USE_��,`Pk�CTReTYhP�0�q P�YN��AAe�V)хQM����ѷ��@O� YA�TINCo�ڱ�B�DՒ�WG֑ENC����u��.A�2Ӕ+@INPO�Q�I6Be��$NT|�#�%NT23_�"ͲIcLO� Ͳ_`��I�_�if� _�k�? ȼ` ej�C400fMOSI�A���ОA䃔�PERCH  �c��B" �g��c��lb =�����oUu@�@		A6B(uLeT	~��1eT�ljgv�fTRK@%�AY��"sY��q 6B�u�s۰�]��RU��MOMq�ՒY�MP�^��C�s�CJR���DUF �BS_BCKLSH_C6B )����f���St�H��R�R��QDCLALM�-d���pm0��CHK����GLRTY ���d��Y��)Üd'_UM]�ԉC��A�!�=PLMT� _AL�0��9��E� .� ��#E)�#H� =�0�Q3po�xPC�ax�HW�頿EׅCMC�E��@�GCN_,N�D�Ζ�SF�1�iV oR��g<!��0r���7CATގSH)�, �DfY��f��7A����܀PAބ�R_P݅�s_ �v��X�s����JG�T]��Y�����TORQ�UaP��c�yPOU`��b��P%�_W�u �t��1D��3C��3C�UIK�IY�I�3F�`6�����@VC�00RQ�t��1���@ӿ��ȳJRK������UpDB M��UpM�C� DL�1BrGR�VJ�Cĭ3Cĳ3$�H�_��"�j@q�COS~˱~�LN���µ �ĭ0�����u�����ē��Z���f$�MY���؊���>�TH�ET0reNK23��3hҧ3��CBm�C5B�3C! AS� ��`u��ѭ3��m�SB�3���x�GTS$=QC������������$DU��Kw�B�%(��%Qq_��a��x�{�K���b(��\сA`Չ��p�{�{�LCPH~�g�Aeg�Sµ ��������g������֚�V��V��0��UV��V��V��V��UV	�V�V%�H��@������G�����H��UH��H	�H�H%��O��O��OV	��O���O��O��O��O*	�O�O�Fg����	�����SPBA?LANCE_-��LE��H_`�SP�!1��A��A��PFULCElTl���.:1��UTO_<����T1T2��22N���29`�!�q�nL�=B�3�qTXpO�v 
A4�INSEG�2�aREV��`agDIF�uS91�8'6t"1�`OB.!t��M��w2�9`��,�L�CHWARRCBA	B�� ��#�`-ФQ 5�X�qPR��&���2�� 
�""��1neROB͠CR0r|5�����C�1�_��T � x� $WEIGH��P`$��?3àI̡Qg`IFYQ�@LA�G�Rq�S�R �RBILx5OD�p�`V2ST�0V2P!t�W0P�11�&1/0�30
�Px�2�QA  2řd^[6DEBUg3L_@z�2�MMY9&E� Nz�D`$D�_A�a$�0��O� � �DO_:@A.1� <B0�6��m�Q�B�2�0N�-cdH_p`�P��2O��� �� %"��T`"a��T/!�4�)@TICKh3| TE11@%�C ��@N͠�XC͠R?��Q�"�E��"�E8@PROMP��SE~� $I�R��Q��R;pZRMCAI)��Q�R4U_r0C2S; �q�PR8�7COD�3FU�Pd6ID_[�vU R!�G_SUFFu� �l3�Q;Q�BD�O�G �E�0�FGR r3�"�T�C�T�"�U�"��Uׁ�T8D�0�B0Hnb _FI�19*c7ORD�1 50�2�36V�+b�Q1@$�ZDT}U 1�0;E��4 *:!L_N�AmA�@�b�EDEF_I�h�b�F�d�E�2��F�4�F�c�E�e�FISP��PAKp�Ds�C�d��44בi��2�D�"�It�3D�O|#OBLOCKEz���S�O�O�Gq�R�PUM�U�b�T�c�T�e�T !r�R�s�U�c�T�d�R �6�q�S� ���U�b��U�c�S�Z��X�@P@` t�@qe�)@W�x4���s 1TE�<D��( l1LO�MB_��ɇ0V2V�IS;�ITYV2A���O�3A_FRI��a SIq�Q!R�@��@�3�3V2�W��W�4����_e��QEAS^3�Rϡ���_�[p:R�4�5��6_3ORMUL�A_Iz���TH]R^2 �Gtg�30�f��<8�5COEFF_O�A	 ��A���GR�^3Sg0BCAnO/C$��]30�1�GRP� � �G $�p�YBX�@TM~w���u�B�s��bCER, Tttsd$`7�  �LL�TSpS~�_SVNt�ߐĸ�$`�@��$`� ���SETUsMEA*P�P��W0�1+b>/0� � h��  @ڐo�l�o�cqDz��b�@cqq`t�P�G��R�� Q\p�*q[p��>�c NPR�EC>at��ASKy_$|�� PB1?1_USER�e"��{ ���VEL@���{ 0�$Ō!I]`���MT�ACFG>���  �@@ =O�"NORE-0l@,o�V�SI.1�d��6��"UXK�fP!��D�E�� $KE�Y_�3�$J3OG��0SV���0���!��}�SW�"�ah\aS�ՐT|�GI����| ^�� 4 �h��'d2�!XYZ�c���31�_ERR#�� 8Ԡ�A�fPV�d��1����/$BUF��X�����MOR|�� HB0CUd�lA�!��GQ�\aB�,"!a$� ���a��u��?��G~�� � $cSIՐ���VO��<T�0OBJE_���ADJU)B��EL�AY���%�DR�O�U.`=ղВQ0b=��T���0���;BDIR���; I�"�0DYNW�2��T���"R���@�0�"��OPWORK����,%@SYSBUy�SOP��ޑ�U�; P�pN�<��PA�t�>�"��OP�PUd!0�`!�Ľl�IMAGw��B0y�2IM�Õ�I�Ne�d��RGOVCRD��-��o�Pq����0��J�Os���"L�pBa���o�PMC�_Ee`���1Ny M� A�21�2T���S�L_��� � $OVSL�ǫ�?qD�`��2�" -�_�� k�P��k�Pu���2�C� �`�Ź�^��_ZER�D��$G�� 82=���� @*����%Oh`RI��� 
 JP8+��=!/��L��ح�T� �0A�TUS��TRC_T���sB��}f�s�9s�1Re`��� !DFAm����L���"`��0a� ޱ��XEw {�����C0�vUP��+p	qPX�P�j�43 � ��PG\���$SUBe�%�qe9JMPWAIT ,z}%LO��F�A�RCVFBQ�@x"�!qR�� �x"ACC� �R&�B�'IGNR�_PL9DBTB2�0Pqy!BWbP�$2w�Uy@�%IGT�P=I��TNLN�&2�R��rL�NP��P�EED \HADCOW�06�w��E[pq4jO!�`SPDV!� LbAz�`�07�3UNIr��02"!R��LYZ`� �o/PH_PK���e�RETRIE9{�q���0'P;FI"�� �G`�0�D 2�g�DB�GLV�#LOGS�IZ��EqKT�!Ud��VDD�#$0_T�
G�MՐCݱ��|@eM�RvC}�3�CHECAK0���0O�V!�kЙI��LE(!��P�ArpT�2K�W��0I�P2V!� h $ARIBiR� c�a�/�O�P8�ӐATT ��2�IF|@z�Aq4S��3UX����PL9I2V!� $g���OITCHx"[�W ��AS9�wSLL�BV!�� $�BA�DYs��BA�M!���Y9�PJ�5��Q��R6�V�Q_�KNOW�Cb��UF��AD�XV��0D�~+iPAYLOAt���Ic_��Rg�RgZ�OcL�q��PLCL=_�� !7��bP�QB��d���fF�iAC֠�js��d�I�h!Rؠ�g�ҢdB���љJ��q_J�a#���AND��Ĳ.t�bؤaL!q�PL0AL_ �P�0���QTրC��DNcE����J3CpWv� TPPDCK������>P�_ALPHgs�s�BE��gy|��K�1�� � �\��HoD_1Oj2ydDP�AR�*��;��&���TIA4U�5:U�6��MOM��a����n���{�Y�B� A�Da���n���{�PUB��R��҅n�҅{��/2�Wp��W � � PMsbT� �BxQ���� e$PI��81���TgJ��niJ�IV�Id�Ir��[��3!��>!��r�Ӫ�U3HIG�SU3�%�4� �4�%� ���"����!x
��!�%SAMP����^��_��%�P4s ю���[ 	ӝ� 3 ���0���&�C��� ��^��Sp��H&0	�IN�SpB�������"��6��6�V�GA�MM�SyI�� E�Tْ��;�D�tA�
�$ZpIBR!62I.T�$HIِ_���$C�˶E��ظAҾ���LWͽ�
���7Ơ��rЖ,0�qC�%C�HK��" �~I_A�����Rr� Rqܥ�Ǚ��ԥ���Ws� �$�x �1���I7RCHk_D�!� RN{��#�LE��ǒ!,���x���90MSWF�L�$�SCR((1#00��R@��3]B�րç��a����َ0��P�I3A9�METHaO����%��AXH��XX0԰62ER)I��^�3��R�0$u�	��pF{�_���$?ⲣ1�L�L�_�a�OOP����wᲡN��APP:���F��`�@{���أRT�V�OBp�0T����;��� 1�I��� ��lr���RA�@MGA1o���SSV-�w�P_@CURg��;�GRO[0S_�SA�Q��Y�#NO�pC!"�tY�� Zolox�������!b��,��&�DO�1A���A ����Х��A���A"�0WS�c L"h�*�� � ��YQLH�qܧ��SrZ�]B�o�=�q�Ô�q_�C1��M_W���g���c�M� �`Vq�$Ap�x1o�3"�PMJ�,�� �'A� 9�!YWi:�$�LWQ |ai�tg�tg�tg{t� �N`���S��JSpX�0O�sRqZ���P� *�� ���M��������������PX��� ��5L�q_~R� |�q#(Y����& n��&{�Y�Z��'�&t���Q��D�#0��@�}`�$PQ�PMO�N_QUc� �{ 8�@QCOU��n%PQTH��HO�n^0HYS:PES�RF^0UEI0O��0O|T�  �0PGõz�RUN_TO�r@Oْ.�� PE`�5C��A<�IND}E�ROGRA�nP� 2g�NE_NO�4�5IT��0�0�INFO�1� p�Q�:A��$PA�B� (��SLE�QݖFAѕF@�6� OySy�T� 4�@�ENAB��0PT�ION.S%0ERV�E���G���1{BGC]F�A� @R0J$�Rq�2���R�H�O�G "�EDITN�1� �v�K�jޓʱE�NU0W�*XAUTu�-UCO�PY�ِN\����M�ѱNXP\[q�PRU�T9� _RN�@OUC�$G�2�T����$$CL`?0[��&������Г �P�S�@�X��PXK�QIGRTU��_�PA� _WRK 2 e��@ 0 � �5�QMoYh\Jo|m |l	�`�m�o��`��o�o�f�e�l}�aI�[ct'`BS�*� �1�Y� <7����� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P��b�t���������srC�C��LMT?0����s  dѴIN�ڿ�дPRE_EXE��)�Ƅ0jP���za'`DV��S��@e)�%s�elect_macro����kϤ�qt�IOCNVVB�� 5��P��USňw����0V 14kP $$p��a�|�`?���߰>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ ���$�ѰLARMRE?COV ^������LMDG ��Ь�LM_�IF ��d�(SYST-32�3 Collab�orative �speed li�mit (TCP?) ) ed���� ���9�K�]�o���, 
 ��C��8TEL�EOP ǘLIN�E 0ǑAUTO� ABORTED�ǘJOINT 1�00 %�����$!���1���A���ROG-057� Power F�ail Reco�v��memory� is cleaAr쏹�˯ң��Ѱ�NGTOL  �@� 	 A  � ��ѰPPIN�FO �� �f�L�^�p����  ������k���ۿſ �����5��Y�C�i���%���ү������ ����'�9�K�]�o���ߓߙ�PPLIC�ATION ?�t��|��Handli�ngToolǖ �
V9.40P�/17���
8g834ؒ��F0�	�549��������7DF5�О�Ǔ�None��F{RA�� 69����_ACTIVE�1�  �� �  \��ސMOD���������CHGAPO�NL�� �OU�PL[�1	��� �>�B�T�f���CU�REQ 1
�� � Tp�p�p�	 ��������l��������������i3l�wp����^H��A�t
HTTHKY�FX v|��*< N`������ ��//&/8/J/\/ �/�/�/�/�/�/�/�/ �/?"?4?F?X?�?|? �?�?�?�?�?�?�?O O0OBOTO�OxO�O�O �O�O�O�O�O__,_ >_P_�_t_�_�_�_�_ �_�_�_oo(o:oLo �opo�o�o�o�o�o�o �o $6H�l ~������� � �2�D���h�z��� ����ԏ���
�� .�@���d�v������������TO�����DO_CLEAN�|��E�NM  �� p�������ɯ�ۯv�DSPDRY�RL���HI��o�@ ��G�Y�k�}��������ſ׿����ϻ�MAX��,�����=��X,�<�9�<���PL�UGG,�-�9���P�RC��Bm�q��6�(ϗ�O����SEGF�K���� � m��G�Y�k�}ߏ�����LAP$�7ޡ�� ����+�=�O�a�s������� �TOT�AL_ƈ� �USE+NU$�1� �������RGDISPWMMC�d�C�&O�@@�1�O"�D���-�_STRI�NG 1��
��M��S���
��_ITEM1��  n������� �� $6HZl ~��������I/O S�IGNAL���Tryout M�ode��Inp�NSimulat{ed��Out`OVERR!�� = 100��In cyclT���Prog A�borj��JS�tatus��	H�eartbeat���MH Fauyl��Aler� !/!/3/E/W/i/{/8�/�/�/ (��� (����/??&?8?J? \?n?�?�?�?�?�?�?��?�?O"O4OFO�/WORИ�~A�/XO�O �O�O�O�O __$_6_ H_Z_l_~_�_�_�_�_8�_�_�^PO��� "`�KoEoWoio{o�o �o�o�o�o�o�o /ASew��bDEV%n�p9o�� ��#�5�G�Y�k�}� ������ŏ׏������1�C�PALT �-j��OD�������ȟ ڟ����"�4�F�X� j�|�������į֯X�GRIB������� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�z�����R�-�� &����������"�4� F�X�j�|ߎߠ߲�������������PREGn�W���0�~�� ������������ � 2�D�V�h�z����������$�$ARG_�~@D ?	����� � 	$$	+[]�$:	���SBN_CONGFIG�XW�qRCII_S?AVE  $z�m��TCELLSETUP 
�%  OME_I�O$$%MOV�_H� ��REP���#��UTOBA�CK� 	t�FRA:\D�c .D�z '`�9D�w� �s � 25/�11/29 20�:26:16D��;D���#//h��C/j/|/�/�/�/�/D�X/�/??(?:? L?�/p?�?�?�?�?�? �?g? OO$O6OHOZO �?~O�O�O�O�O�O�O����  c_F_�\ATBCKCTL.TM�)_;_M_�__q_8INIm��j~CMESS�AG� �Qz �[O�DE_D� �j��XO�p�_@PAU�S6` !� ?, 	�; <:oHg,		2olo Vo�ozo�o�o�o�o�o �o 
D.Pz}d~`TSK  mxw}_CUPDT�P�Wd�p�VXWZD_ENB�Tf
�v�STA�U�u��X�ISX UNT 2t�vwy � 	�p��P�v��� ��C l .��D�R�  /�������Q��m������R�.�1o����[ #�g o� ��y������,�/�M[ET��2@��y �PQ�A�d�A��1AZ��A�;�A]ˢA��F��>z��>�%;>$�H<��ԡ?��>�}��5�SCRD�CFG 1�Y ��w ����%�7�I�pD�Q�	ܟ������ϯ ��Z��~�;�M�_��q�������6���FG�R9��p�_ԳPNA�� 	FѶ_�ED�P1��� �
 �%-PEDT-¿ R�v����E�<�GE�D��;9/�>���  ����2�����B�  ����{�����j�����3��#� �G�Y���@G�ߠ�6�����4� �����Yި��Z�l������5K������ Y�t���&�8���\���6��d��Y�@� ���(��7�S 0wY�w��f����8�W��{�I Z��C/��2/���!9{/��//LZݤ/�?V/h/�/�/��CR ���?�?Tn?�? ?�2?�?V?԰!�NO_�DEL�ҲGE_�UNUSE޿дI�GALLOW 1��   (�*SYSTEM�*
�	$SER�V_GR[�@`REG�E$�C
��@�NUM�J�C�MP�MU?@
�LA�YK�
�PM�PAL�PUCYC10 N3^P!^YSULSU_�M5Ra�CLo_�TBOX�ORI�ECUR_��P�MPMCNV6V�P10I^�PT4DLI�p�_�I�	*PROGRA��DPG_MI!^Ko]`AL+ejoTe�]`B�o�N$F�LUI_RESU`9W�o�O�o�dMR�N�@�<�?�;M_ q������� ��%�7�I�[�m�� ������Ǐُ�����!�3�E�W�2BLAL_OUT �K����WD_ABO�R:PcO��ITR_�RTN  �$��빸�NONSTO��� lHCCF�S_UTIL ��̷CC_AU�XAXIS 3$� h}�j�|������ƽCE_RIA3_I`@�נ���FCFG �$�/�#��_L�IM�B2+� ��8p� 	��B\T���$8p
Ԡ��)[�Z�%�/�����[�����.R���!$�����L��(
5������PA�`GP 1H�����A�PS�e�w�6�CC� �C7��J��]��p�������� C�����������������é�̩�ձ�ߪ���������;L���PCk�������U�������������ɱ���������� D� D�!�!�!�!� m��&?��HE@�ONFIpC�G�_P�P1H� +EH��ߟ߱�����������C�KPAU�S�Q1H�ף  IR�S�H�A��e�� ������������� E�+�i�{�a����A?Iץ�MؐNFoO 1���� �3��$4�A����Aԫ���g2�@C�0���B�J��*� D�@B�Qs�A��*C�2�/?��kBG��Pb�O�� � ��LLECT_�!�����EN+`�ʒ����NDE�#��/�1234567890�"�A���/ҵHw��#) j��<i{��;� �/��/`/+/=/ O/�/s/�/�/�/�/�/ �/8???'?�?K?]? o?�?�?�?�?O�?�:�$� ��IO &��"S�▒O�O�O�O`GT-R�2'DM(��^�?�NN�(oM Z���_MOR)q3)H��7ىU3��Y�_�_��_�_�_�[bR�kQ*JH�,S�?<�<Ѡ<c�8pKFd���P,��;ϒo�o�o˿��o�oœh�UY@�E�oS �wsja�PDB�.���4cpmi�dbg3��Рs:���>uqpz��v/  ��>x���}.��}�`��|�<�mgP���t��~�f������@u�d1:�?��XqD�EF -��zC)�*�cO�buf.txtJ��|K�[`��/DM��>����R�A��MCiR20�_{RCd���hS21b����G���CzA��d4�EI�jA���]\ �F]� �B�e;t�H��j�C1�aCN�/�I؂�DH󇳜�LڒY�E�E�>��MSo�F��&�ġ�����f23FDLD�	>	P!� Y2��}��yc
�@�x9� C�Ĵ�  D4G�E����  E%q��F�� E�p��u�F�P E���fF3H ?��GM��Ъ>5�>�33��?��xn9�q@�Q5�����RpA?a��=�L��<#�QU��@,�Cϒ���RS�MOFST +xi�����P_T1Ɠ�4DMA =ք�M?ODE 5dm�@c��	Q�M;���%��?���<�M>��Ͷ�/TESTc�2i�`�ER�6�O�K�CN�QAB���n� 8��\�n�CdB���C�pp����	P:;d�QS ��ՠ ������4�I7R>���>B8m5�$�RT_c�PRO/G %j%��d�|1�h@NUSER���x�KEY_TBL�  e�����	�
�� !�"#$%&'()�*+,-./(:�;<=>?@AB�Cc�GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������>���͓���������������������������������耇���������������������8�LCK��F�y��OSTAT��2�X��_ALM�����_AUTO_DO��E�FDR 3�:i�2h&q[~��� BUO�SYST-322� Auto st�atus che�ck time out ���i�$TELEO8|�i� ��)q�A�ʜ@Ĭ������?�ڛ�MsB�õ��?*?���?Mf=�o�TR��-����D.�B����C���B�yN�*p�4�N�4�J5Hj5H���>�i�BJ�d�B�F�	PZ��[~�b bt����5/��M*F�B�G�A+$����@R��J�}�BQ�H����������2�>��@�@����&��CBxHCKH<B��6>Tbt ��/��u�US�H?Z?l?i�$7?�?:��  mϸ?�?p���?�?O O�?,OfOxO�M6?�O �O�O~?�O	_�?*_$_ BOD_6_p_~_T_�_�_ �_�_�Oo)o;o�OLo qo_�o�o�_�o�o�o �o�o�oFXo ��No���o�� ��@�N�$�b�x� ����n������ A��b�\�z�|�n��� ����ʟ���(�֏O� a�s������T�ʯį ��֯����2�H� ~���>���ɿۿ��� ϼ�2�,�J�L�>�x� ��\Ϛϰ����Ϧ�� 1�C��T�y�$Ϛߔ� �ϴߦ��������� N�`�߇���V߼� ���������H� V�,�j�������v��� ��$I��jd ���v����� 0��Wi{&� �\�����/ &/�:/P/�/�/F�/ �/�/��/?�:?4? R/T?F?�?�?d?�?�? �? O�/'O9OKO�/\O �O,?�O�O�?�O�O�O �O�O
_ _V_h_O�_ �_�_^O�_�_�O
oo "_$ooPo^o4oro�o �o�o~_�o	�_, Q�_rl�o�~� ����&�8��o_� q���.����dڏԏ ��� �.��B�X� ����N�ǟٟ럖��� !�̏B�<�Z�\�N��� ��l����������/� A�S���d���4����� ¯Ŀ�����Կ�(� ^�p���ϩϻ�f��� �Ϝ���*�,��X� f�<�zߐ����߆��� �#���4�Y��z�t� �ߔ����������� .�@���g�y���6�� ��l�����������( 6J`��V�� ����)��JD bdV��t�� �/�7/I/[/l/ �/<�/�/��/�/�/ ?�/?0?f?x?&/�? �?�?n/�?�?�/OO 2?4O&O`OnODO�O�O �O�O�?__+_�?<_ a_O�_|_�O�_�_�_ �_�_�_ o6oHo�Ooo �o�o>_�o�ot_�o�o o�o0>Rh ��^o����o� 1��oR�L�jl�^��� ��|���Џ���?� Q�c��t���D����� ҏԟƟ ���"�8� n���.�����˯v�ܯ ���"��:�<�.�h� v�L�����ֿ迖�� !�3�ޯD�i���τ� ���ϖ����ϴ���� >�P���w߉ߛ�FϬ� ��|�����
����8� F��Z�p���f��� ������9���Z�T� r�t�f�����������  ��GYk�| �L������� �*@v�6� ��~�	/�*/$/ BD/6/p/~/T/�/�/ �/�/�?)?;?�L? q?/�?�?�/�?�?�? �?�?�?OFOXO?O �O�ON?�O�O�?�O�O O__@_N_$_b_x_ �_�_nO�_�_o�Oo Ao�Obo\oz_|ono�o �o�o�o�o(�_O aso��To�� �o�����2�H� ~���>��ɏۏ�� ��2�,�J�L�>�x� ��\����������� 1�C��T�y�$����� ��������į�� N�`��������V��� ῌ�������H� V�,�jπ϶���v��� �߾�$�I���j�d� �τ�v߰߾ߔ����� �0���W�i�{�&ߌ� ��\������������ &���:�P�����F�� ����������:4 R�TF��d�� � ��'9K��\ �,������ ��
/ /V/h/�/ �/�/^�/�/�
?? "/$??P?^?4?r?�? �?�?~/�?	OO�/,O QO�/rOlO�?�O~O�O �O�O�O�O&_8_�?__ q_�_.O�_�_dO�_�_ �O�_�_ o.ooBoXo��otc�$CR_F�DR_CFG };re�Q?
UD1:�W�P:�aJ�d  �`�\��bHIST 3<�rf  �`  w?�R@tuAtB�bC�PU,pDtEtItUg�Ppotw�_���bINDT_E�N6p�T��q�bT1_D�O  �U�u�sT�2��wVAR 2m=�gp hq�  �4�f�4��R�5H4��5H�m[��RZ�`S�TOP��rTRL?_DELETNp�t� ��_SCRE�EN re�r_kcsc�rUw��MMENU 1>~��  <�\%�_��T��R��S /�U���e�w�ğ���� ��џ�	�B��+�x� O�a�����������ͯ ߯,���b�9�K�q� ������࿷�ɿ�� ��%�^�5�Gϔ�k�}� �ϡϳ��������H� �1�~�U�gߍ��ߝ� ��������2�	��A� z�Q�c������� ����.���d�;�M� ��q�������������YӃ_MANUA�L{��rZCD�a�?�y�rG ����R�f"
�"
?�|(��PdTGR�P 2@�y�cB� � s��~� �$DBCO�p�RIG���v�G_�ERRLOG 	A��Q�I[m� �NUMLI�M�s��u
�P�XWORK 1B�8���//��}DBTB_�� CC%���S"�� �aDB_AWA�Y��QGCP Ϋr=�ןm"_AQL�F�_�Yz�����p�vk  1D
�Ap
��/"�/�%?/(_M�pqw,@}�=5ONTIM�����t�_6�)
��0�'MOTNE�NFpF�;RECO�RD 2J� y�-?�SG�O��1 �?"x"!O3OEOWO�8 _O�O�?�OO�O�O�O �O�O(_�OL_�Op_�_ �_�_A_�_9_�_]_o $o6oHo�_lo�_�o�_ �o�o�o�oYo}o2 �oVhz��o� �C�
��.��R� �K��������Џ?� �ߏ�*�����+�b� t�㏘�����Ο=�O� ����:�%���p�ߟ 񟦯��O�ǯ�]�� ����H�Z������� ��#�5����ϩ�i"�TOLERENC�v$Bȿ"� L���� CSS_CCS_CB 2K�\0"?"{ϰϟ��� 7��
����@�R�d�3߈ߚ�"�x����� ����'�9�K�]�o� ������������� �#�5�G�Y�k�}��� ������������ 1CUgy���C ������VR�LL]�La�m1|T#2 C��C��F�^ A��C�pC���#�0��� 	 A�̃�B���?�  �$����\0c袰�0��B�ƀ`#s�K/]/o/�ϓ/�/�/s/�/�/��K��KP����5ѹ�0�����CȦ�D�/��/`?;�@��O?�?�?�?�0AF��?{F�A  OO�7�1���9M	AB
AZOdBAE�9$OP�O�O�Oi:P��`�@�0�DJCA�� @��
X8-.
[#_   M?�>O�ڴ�q_�_�_�_:W�A<o:[< ǲ/o�/�_+oPo0boto�eACHC�V��WB$�Dz�cD �`�a=/�o�oo�oW$�a.+!��2=t,y �J?�.s�s�js�w �yj�������Q�Qs�@`��$� ����A����Bމ�o ��'�9��_]�o�N� ��r���ɟ۟_�B��ʄ��YZ>`��(��B�O�A�i��@-D�=g=�8��w�Z�l�~����`_м¯ ���
���̯9�,�]� o��� �H�����ٿ� ���ƿ3�E�W�iϬ� ��$ϱ����� Ϟ�� ��/�A�S߶�w�V�h���ߌ��S���ߐ� _�f	��H�?�Q�~� u���������� ��D��-�g�q��� ����������
 @7Icm��߾�  ����� )M@qdv� ������// I/P�m/�v/�/�/�/ �/�/�/�/?3?*?<? i?`?r?�?^/�?�?�? �?�?O/O&O8OJO\O �O�O�O�O�O�O�O�g�	  Q��P�s �P+C4p*p�p6U\6P\C9p/pG�� ]V^PM]�6P��:P�>P�VJ_�
^P�bP�fP�Vr]v���p Q
k���_�oo�id1Q&oNo �;o_co�oˏUUA�   �o�k1Q@�C  �o�k�b������p �� �1��6�w1C���CA�cPfL��?#�c�>�{���`�cP�@@�d��r�`�B�cP>�s�qC�Ϋp����b�t<��o?�PH�)S�B�tq�q�p�r�`B���eIC�&�Q�4( �oz�UU��:�P�A�j��@-F�=f�c�8���Q�-R����0��}¿�`B��8b@y��`ځ`  ?�p����U�[?����}t��$���$DC�SS_CLLB2� 2M���p�P�^?�NSTC�Y 2N��?�  ��� ����ʟ؟���� � 2�D�Z�h�z��������¯ԯ��SA�DEV�ICE 2O��!�$��4&V�h��� ����˿¿Կ���
� 7�.�[�R�ϑϣϵ������4(A�HNDG�D P��*�Cz|�A�LS 2Q��_�Q�c�u߇ߙ߫������?�PARAM RP��1�`�&տRBT 2T��/ 8�P<C�'pG �qi�l��sF@"�R��(qI�X���0�pB CW  ��B\x�N��`Z��&���%��)���X�@j��p����zq�����B �(s,�F�p��V��q���b��B ��4&c �S�e�l�4+�����H1~�����D�C�$Z|��b���A,� �4�u@�X@��^@w���]�B���B�cP%���C4�C3�:^C4��n��� ��p8�-B�{B��A����� l��C��C3�JC4jC3��yn�+�3 Dff 2�A PB W4+@:�]o�W�� ���/�/P/'/ 9/K/]/o/�/�/�/�/ ?�/�/�/?#?5?�? Y?k?�?�?�o�?�?O �?6O!OZOlOWO�O�E s�?�?�?�O�O_�O �OL_#_5_G_Y_k_}_ �_�_�_ o�_�_�_o o1o~oUogo�o�o�o �o�owO D/A ze����O�o�o 
��o��R�)�;��� _�q����������ݏ �<��%�r�I�[�m� �������ǟٟ&�8� �\�G���k������� گů�����F�� /�A�S�e�w�Ŀ���� ��ѿ�����+�x� O�aϮυϗϩϻ��� ��,���b�t�ﯘ� �߼ߧ��������� :��C�U߂�Y�k�� ����������6�� �l�C�U�g�y����� ������ ��	- ?Q������ �@+dvQ� ������� *///%/r/I/[/�/ /�/�/�/�/�/&?�/ ?\?3?E?�?i?{?�? �?U�?�?"O4OOXO CO|OgO�O{��?�O �?�O�O0___f_=_ O_a_s_�_�_�_�_�_ o�_oo'o9oKo�o oo�o�o�o�o�o�O :%^I�������H�$DCS�S_SLAVE �U���	����z_4D�  	��AR_MENU V	� �j�|�������ď��BY�� ��~?�S�HOW 2W	� � �b�aG�Q� X�v���������П֏���� @�:�d�a� s����������߯� �*�$�N�K�]�o��� ����̯ɿۿ��� 8�5�G�Y�k�}Ϗ϶� ����������"��1� C�U�g�yߠϝ߯��� �����	��-�?�Q� c��s��������� ����)�;�M�t��� �������������� %7Ip�m�� ��������! 3ZWi���J ����//DA/ S/e/��/��/�/�/ �/�/?./+?=?O?v/ p?�/�?�?�?�?�?�? ?O'O9O`?ZO�?�O �O�O�O�O�OO�O_ #_JOD_nOk_}_�_�_ �_�_�O�_�_o4_.o X_Uogoyo�o�o�o�_ �o�o�ooBo?Q cu���o:��~�CFG X)��3�3q5p��FRA:\!�L�+�%04d.CS�V|	p}� ��qA g�CHo�z@v�	����3q�����́܏� ���4��JP����q�p1� �RC_�OUT Y���C��_C_�FSI ?i� .����� ��͟�����>�9� K�]���������ίɯ ۯ���#�5�^�Y� k�}�������ſ�� ���6�1�C�U�~�y� �ϝ����������	� �-�V�Q�c�uߞߙ� �߽��������.�)� ;�M�v�q����� �������%�N�I� [�m������������� ����&!3Eni {������� FASe�� ������// +/=/f/a/s/�/�/�/ �/�/�/�/??>?9? K?]?�?�?�?�?�?�? �?�?OO#O5O^OYO kO}O�O�O�O�O�O�O �O_6_1_C_U_~_y_ �_�_�_�_�_�_o	o o-oVoQocouo�o�o �o�o�o�o�o.) ;Mvq���� �����%�N�I� [�m���������ޏُ ���&�!�3�E�n�i� {�������ß՟���� ��F�A�S�e����� ����֯ѯ����� +�=�f�a�s������� ��Ϳ�����>�9� K�]φρϓϥ����� ������#�5�^�Y� k�}ߦߡ߳������� ���6�1�C�U�~�y� ������������	� �-�V�Q�c�u����� ����������.) ;Mvq���� ��%NI [m������ ��&/!/3/E/n/i/ {/�/�/�/�/�/�/�/�3�$DCS_C�_FSO ?����71 P ??T? }?x?�?�?�?�?�?�? OOO,OUOPObOtO �O�O�O�O�O�O�O_ -_(_:_L_u_p_�_�_ �_�_�_�_o oo$o MoHoZolo�o�o�o�o �o�o�o�o% 2D mhz����� ��
��E�@�R�d� ��������ՏЏ�� ��*�<�e�`�r��� ������̟����� =�8�J�\�������?_C_RPI4>F? �������3?�&��o����� >SLү@ d������%�7�`� [�m�Ϩϣϵ����� �����8�3�E�W߀� {ߍߟ���������� ��/�X�S�e�w�� �����������0� +�=�O�x�s������� ������'P K]o����� ���(#5Gp k}�����Q�� �/6/1/C/U/~/y/ �/�/�/�/�/�/?	? ?-?V?Q?c?u?�?�? �?�?�?�?�?O.O)O ;OMOvOqO�O�O�O�O �O�O___%_N_I_ [_m_�_�_�_�_�_�_ �_�_&o!o3oEonoio {o�o�o�o�o�o�o�o FASe�������>�NOC�ODE ZU���?�PRE_CHK \U���pA �p�< ��pU�]�o�U� 	 <Q����� ���ۏ�Ǐ�#��� �Y�k�E�����{�ş ן��ß����C�U� /�y�����s���ӯm� ��	���?��+�u� ��a�������ɿ�Ϳ ߿)�;��_�q�K�}� �ϝ������ω���%� ���[�m�Gߑߣ�}� ���߳����!���E� W�1�c��g�y����� ���������A�S�-� w���c����������� ��+=asM _������ '�]o	�� ����/#/� G/Y/3/e/�/i/{/�/ �/�/�/?�/?C?9 Ky?�?%?�?�?�?�? �?	O�?-O?OOKOuO OOaO�O�O�O�O�O�O �O)_____q_K_�_ �_a?�_�_�_�_o%o �_Io[o5oGo�o�o}o �o�o�o�o�o�oE W1{�g���_ ����/�A��M� w�Q�c���������� Ϗ�+���a�s�M� ��������ߟ��� '���3�]�7�I����� �ɯۯ������� G�Y�3�}���i���ſ ��������1�C��� +�yϋ�eϯ��ϛ��� ������-�?��c�u� Oߙ߫߅ߗ������� �)��M�_�U�G�� ��A����������� ��I�[�5����k��� ����������3E Q{q���] ����/Ae wQ������ �/+//7/a/;/M/ �/�/�/�/�/��/? '??K?]?7?�?�?m? ?�?�?�?�?O�?5O GO!O3O}O�OiO�O�O �O�O�O�/�O1_C_�O g_y_S_�_�_�_�_�_ �_�_o-oo9oco=o Oo�o�o�o�o�o�o�o __M_�ok� o������� �I�#�5����k��� Ǐ��ӏ��׏�3�E� �i�{�5c���ß�� ���ӟ�/�	��e� w�Q�������ѯ㯽� ϯ�+��O�a�;��� �����Ϳ߿y��� �!�K�%�7ρϓ�m� ���ϣ���������5� G�!�k�}�W߉߳ߩ� �����ߕ��1��� g�y�S������� �����-��Q�c�=� o���s��������� ����M_9�� o����� 7I#mYk� �����!/3/) /i/{//�/�/�/�/ �/�/�/?/?	?S?e? ??q?�?u?�?�?�?�? OO�?%OOOE/W/�O �O1O�O�O�O�O__ �O9_K_%_W_�_[_m_ �_�_�_�_�_�_o5o o!oko}oWo�o�omO �o�o�o�o1U gAS����� �	����Q�c�=� ����s���Ϗ�o��� ���;�M�'�Y���]� o���˟����۟� 7��#�m��Y����� �������!�3�ͯ ?�i�C�U�������տ �������	�S�e� ?ωϛ�uϧ��ϫϽ�������$DC�S_SGN ]�	�E��-����30-NOV�-25 17:1{7 ��29R�O20:2^�x�x� [}�t�ԁq�т�xҚك�JѨ��EƼÞ� ���ǖ�  1�H�OW ^	�� x�/�V�ERSION �=�V4.5�.2��EFLOG�IC 1_���  	�����C���R�%�PROG_�ENB  ���:�{�s�ULSE � X��%�_A�CCLIM������d��WRS�TJNT��E��-�EMO|�zя�$����INIT `�2����OPT_�SL ?		�	�
� 	R575���]�74b�6c�7c�50��1���C�����@�TO  �L��� �V�DE�X��dE�x�P�ATH A=�A�\k}��HC�P_CLNTID� ?�:� �D�ռ��IAG_�GRP 2e	�����z�	 �@�  
ff?aG����B�  2��/�x8[I@c�ς�!�7@�z�@^�@
�!���mp2m15� 8901234�567���� � ?��?��=q?��
?�޸R?�Q�?_��?�����(�?�z��|�x�@�  A_�cAp !7A�8�8_�B4�� ���L�x�
�@��@��\@~��R@xQ�@q��@j�H@c��
@\��@U?�@Mp��/�/'$�; �O)H���@Ct >d 9���@4�/\)@�)� #t {@��/�/�/�/�/~P'?���?����_ ?}p�?�u?n{?vs ?\�Q�?� ?2?D?V?h8�
=K?����0w5��z�H?p�h��?^�R�?�?�?P�?�?h8��t0�e��@�?��0�;@&O8OJO\OnO P'�$_�_Y_k_�O ?_�_�_�_�_�_s_�_ �_1oCo!ogoyoo�o ��Bj"� �2{1�@"/?���f�t0�d�"5!�
u4V��u"�B3t�A>u���?@[q��@`�,=q�=b���=�E1>�J��>�n�>���H"<�o �z�Ss�q��� �xѽC�@<(�Uz�K 4�� ����A@x�?*�o��m *�P�b���tn���2����Ώ�����i>J;��&�bN2�"O��G�N��o@�@�v���0����@�ffr!l ��3�3���(��"C��� ƒI�C�H�)C.dBت"8"����'���"~�A?�&"K�X���pf�B��@�p��������p��<����?蕼����?啼��m<��i<���J���V���RD�@BQs_�A��*x�> � �����0��N�T�����C2�/??��kB�D�#� ����ȿ���׿�����?,�<�o��CT�_CONFIG �f��|��egY��STB_F_TTS��
�頺��О�}���1�M�AU������MSW�_CF��g�  �# ��OCVIEWf��h!�-��� s߅ߗߩ߻��ߟ�a� ����,�>�P���t� �������]���� �(�:�L�^������ ��������k� $ 6HZ��~��� ���y 2D Vh������,�v�RC�i���!���/S/B/w/f/�/�/�/��SBL_�FAULT j�*6��!GPMSK����'��TDIAG� k��-�������UD1:� 6789012345I2��=1�Ǥ�P\υ?�?�?�?�?�? �?OO'O9OKO]OoO��O�O�Od696���r
�t?�O|�TRECP"?4:
B44_[7��s? p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o��o�O�O�O�o7�UMP_OPTIO=��.�aTR����)�uPME��Y�_TEMP  _È�3BC�gp9�B�QtUNI�����gq�YN_BRK� lL�7�EDI�TOR�a�a@�r_~
PENT 1m)�  ,&TELEOP^P ���=�pPSNA�:�&MTPG�p +�=��/��I�z����� ۏ����5��Y� k�R���v���ş��� П����C�*�g�N� v������������ޯ���?�Q���EMGDI_STAzu�V�gq�uNC_IN�FO 1n!��b���X���������vn�1o!� ��o(����
�d�oU� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߽߫��� u���� 
��*�B�*�P�b�t� ������������ �(�:�L�^�p����� ����2������� 9�CUgy��� ����	-? Qcu������ ��//1;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?m?? �?�?�?��?�?�?O )/OEOWOiO{O�O�O �O�O�O�O�O__/_ A_S_e_w_�_�_�_�? �?�_�_o�_3O=oOo aoso�o�o�o�o�o�o �o'9K]o ����_�_��� �+o5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� �ӟ���	�#�-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ���7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� �����������%�/� A�S�e�w����� ��������+�=�O� a�s������������� ���'9K]o �������� #5GYk}� 	������/ 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?��?�? �?�?/O)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�?�_�_�_�_O�_ !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew��_�_� ���o�+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ������ɟ۟�� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߝ��߹������� ���%�7�I�[�m�� ������������� !�3�E�W�i�{��߇� ���������/ ASew���� ���+=O as�������� ��//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?�� �?�?�?�?��?OO 1OCOUOgOyO�O�O�O �O�O�O�O	__-_?_ Q_c_u_�?�_�_�_�_ �?�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m�_ u����_��� !�3�E�W�i�{����� ��ÏՏ�����/� A�S�e�������� u������+�=�O� a�s���������ͯ߯ ���'�9�K�]�w� ��������ɿ���� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g߁��ߝ߯� ��ۿ����	��-�?� Q�c�u������� ������)�;�M�_� y߃������������� %7I[m ������� !3EWq�c�� �������//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? i{�?�?�?�?��? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_�?s?}_�_ �_�_�?�_�_�_oo 1oCoUogoyo�o�o�o �o�o�o�o	-? Qk_u����_� ����)�;�M�_� q���������ˏݏ� ��%�7�I�cQ�� �������ٟ���� !�3�E�W�i�{����� ��ïկ�����/��A�[� �$ENE�TMODE 1p���� + k�k�f������j�OATCFG� q�����Ѵ��C���D�ATA 1rw��Ӱ���*	�*@��'�9�K�]�l�dl���e��ϻ����� ����'ߡϳ�]�o� �ߓߥ߷�1���U��� �#�5�G�Y����ߏ� �����������u�� 1�C�U�g�y������ )�������	-�� ��cu������j�RPOST_L%O��t�[
׶�#5Gi�RROR�_PR� %w�%�L�XTABLE  w�ȟ�����RSEV_N�UM ��  ����  �_A�UTO_ENB � ���X_NON5! uw���"_  *�x �x %�x �x + +w �/x�/�/Q$FLTR=/O&HIS#]�J+_ALM 1vw�� �[x,e�+�/Q?c?u?�?�?�?r�/_"W   w��v!���:j�TCP_VER !w�y!x�?$EXT� o_REQ�&�H)�BCSIZKO=DST�KhIf%�?BT�OL  ]Dz��"�A =D_BWD�0�@�&�A���C;DI�A wķ�x��]�KSTEP�O��Oj�POP_DO��Oh�FDR_GR�P 1xw��!d �	�?�_��yPs��Y�Q'�M"����l��?T� ����VyS��_�]yPA
�A����A��PA�$]A���<�]]@՚�b	dAg��oEo�_Bo�{ofo�o�o�o�o>����>�">���3k M8pKx0a�a]?��^�o�(2�o�oZE~�]@<`�t@S33�u�]�@�q�g��yPF�@ ��|yPG��  @�Fg�fCg�8RL��]?�p�i��~6�X�����875t��5����5`+��~w�:��W���s�� �������]%ݓF�EATURE �y���@���Handling�Tool �]�English� Diction�ary�4D S�t��ard��A�nalog I/�O>�G�gle S�hiftZ�uto� Softwar�e Update��matic B�ackup���g�round Ed�it ��Came�raU�FY�Cnr�RndIm���o�mmon cal�ib UI��n�ˑ�Monito�r$�tr�Rel�iabn��DHC�P �[�ata A�cquis3�\�iagnos��R�v��isplayΑL�icensZ�`�o�cument V�iewe?�^�ua�l Check ?Safety��?hanced����s�Frܐ�xt. DIO /�sfi��@�end�Err>�L��\�4�%s[�rP�K� �@
��FCTN Men�u��vZ���TP ;In��facĵ��GigE־�Đp� Mask Ex�c�g=�HT԰Proxy Sv���igh-Spe�Ski�� Ť�O��mmunic��onsV�ur����q��V�ײconnecwt 2��ncrְ�stru!��ʴ�e�ۡ��J��X�KAR�EL Cmd. �L�ua���Ru�n-Ti<�Env��Ȟ�el +��s��S/W�ƥ����r�Book(Sy�stem)
�MA�CROs,M�/OOffseu�p�HO���o�u�MR8�4����MechStop"+�t����p�im�q����x�R�����od>o�witch���.��4�Optm8F��,�fil䬳��g��p�ulti-�T�Γ�PCM 'fun�Ǽ�o���������Regie�r,q���riݠF����S�Num Sel���/�:� Adju�a�*�W�q�h�tat�u��ߪ�RDM� Robot�s�cove'���ea���<�Freq Awnlyq�Rem���O�n5�����Ser�voO�!��SNPgX b-�v�SN԰�Cliܡ?r�Li#br&�_�� ��q �+oJ�t��ssag��X�@ ����	��@/Iս�MIL�IB��P Fi�rm���P��AcycŐ͛TPTXk��eln���������orquo�i�mula=��|u(�Pa&��ĐX�B�&+�ev.���r�i��TUSB �port �iP�f�aݠ&R EV�NT� nexcept�����%5��VC�rl�c��؁V���"�%q�+S�R SCN�/SGE��/�%UI	�Web Pl��>��A4�3��ۡ��ZDT �Applj�
�{1EOAT����&0?�7Grid�񾡬=.�?iR�".5� F����/גRX-10�iA/L�?Ala�rm Cause�/��ed(�All Smooth5�<��C�scii+�V��Load䠌JUp9l�@w�toS ���rityAvoi+dM(�s7�t�@�ycn������_�CS+���. c��XJo���-T3_�H�.RX��U���Xc?ollabo�����RA�:�.9D��iqn���NRTHI�
�On��e Hel����ֿ�����1�trU�ROS Eth$��A������;�,�G �B�,|HUapV�%�W�t ԰��_iRS�ݐ�64MB DRAM�o�cFRO���L8F� FlD�����2M L�A:�opm�ԕex@�V�
�sh�q��wc�e�u��p��|ty"n�sA�
�%�r����J��^�.v� P)Q/sbS�`���O�N��mai��U����R�q�T1�^FC+Ԍ%̋Fs9�ˌk�̋��Typ߽FC�%�hױV�N Sp�F�orްK��Ԭ�lu�!����cp�PG j��֡�RJ�[L`Sup"}��֐f��3crFP��lu� ��#al�����r��i��
q�4@а�ue�st,IMPLE ׀6*|HZ���c0�BTea(�|����$rtu���V�9H�MI�¤��UIFNc�pono2D�B C�:�L�y�p������� ��ʿܿ	� ��?�6� H�u�l�~ϫϢϴ��� ������;�2�D�q� h�zߧߞ߰������ ��
�7�.�@�m�d�v� ������������ 3�*�<�i�`�r����� ����������/& 8e\n���� ����+"4a Xj������ ��'//0/]/T/f/ �/�/�/�/�/�/�/�/ #??,?Y?P?b?�?�? �?�?�?�?�?�?OO (OUOLO^O�O�O�O�O �O�O�O�O__$_Q_ H_Z_�_~_�_�_�_�_ �_�_oo oMoDoVo �ozo�o�o�o�o�o�o 
I@Rv �������� �E�<�N�{�r����� ��Տ̏ޏ���A� 8�J�w�n�������џ ȟڟ����=�4�F� s�j�|�����ͯį֯ ����9�0�B�o�f� x�����ɿ��ҿ���� �5�,�>�k�b�tφ� ���ϼ��������1� (�:�g�^�p߂ߔ��� �������� �-�$�6� c�Z�l�~������ ������)� �2�_�V� h�z������������� ��%.[Rdv �������! *WN`r�� �����//&/ S/J/\/n/�/�/�/�/ �/�/�/??"?O?F? X?j?|?�?�?�?�?�? �?OOOKOBOTOfO xO�O�O�O�O�O�O_ __G_>_P_b_t_�_ �_�_�_�_�_ooo Co:oLo^opo�o�o�o �o�o�o	 ?6 HZl����� ����;�2�D�V� h�������ˏԏ� ��
�7�.�@�R�d��� ����ǟ��П����� 3�*�<�N�`������� ï��̯����/�&� 8�J�\����������� ȿ�����+�"�4�F� Xυ�|ώϻϲ����� ����'��0�B�T߁� xߊ߷߮��������� #��,�>�P�}�t�� ������������ (�:�L�y�p������� ��������$6 Hul~������  Hg552��21�R7850J�614ATUP�'545'6VwCAMCRIb�UIF'28cN�RE52VR6�3SCHLI�C�DOCV�C�SU869'0^2EIOC�4�R69VESET�?UJ7UR68�MASKPR�XY{7OCOB#(3?+ &3j&[J6%53�H�(�LCHR&OPLGz?0�&MHCRS&]S�'MCS>0.'{552MDSW+7vu'OPu'MPRv&t��(0&PCMz�R0q7+ 2� �'5�1J51�80JP�RS"'69j&FR�DbFREQM�CN93&SN�BA��'SHLB�FM1G�82&H{TC>TMIL��TPA�TPT�XcFELF� �8�J95�T�UTv'95j&UE�V"&UECR&UF]RbVCC
XO�&wVIPnFCSC�F�CSG��IW�EB>HTT>Ra6��H;RVCGiW{IGQWIPGS�V�RCnFDGu'H7.�7R66J5']R�8R51
(6�(%2�(5V�J8�8�6�L=I% �84vg662R64�NVD"&R6�'R[84�g79�(4��S5i'J76j&Du0�gF xRTSF�CR�gCRXv&CsLIZ8ICMS�\Sp>STYnG6)7GCTO>��7�;NNj&ORS�&C �&FCB�FCFv�7CH>FCR"&�FCI�VFC�'JԗPO7GBfM�8OLnaxENDS&LU�&WCPR�7LWS�x�C�STxTE�gS�60FVR�IN�7IHaF�я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{���� ���/AS ew������ �//+/=/O/a/s/ �/�/�/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� �������� %�7�I�[�m�������Ǐُ�  ?H552���21�R78�5�0�J614�AwTUP7�5457��6�VCAM�C�RI��UIF7�2�8��NRE�52�v�R63�SCH��LICƚDOC�V�CSU�86�97�0F�EIOC�Ǜ4�R69v�EgSETW�u�J7u��R68�MASK^�PRXY��7�OCO��3W�����6�3�J65�53�6�H$�LCHƪO�PLGW�0�MH�CRǪS��MCS�V�0��55F�MD�SW���OP��M�PR���6�06�PCM��R0E˓�F�l��6�51f�51���0f�PRS��69��FRD��FRE�Q�MCN�93�6�SNBAכ%�SHLB�ME��ּ�26�HTCV�TMsIL�6�TPAV�oTPTX��EL�ē�6�8%�#��J9�5��TUT��95��UEV��UEC�ƪUFR��VCC�f�O��VIP��C;SC��CSGƚ$��I�WEBV�HTTV�R6՜��S����CG��IG��IP�GS'�RC��DGv��H7��R66f��5�u�R��R51*f�6�2�5v�#�)J׼��6��LU�5��s�v�4��66F�R�64�NVD��R�6��R84�79��4��S5�J7�6�D0uFR�TS&�CR�CR�X��CLI&�e�C�MSV�sV�STY:��6�CTOV�#��V�75�NN�ORqS����6�FCBV��FCF��CHV�F�CR��FCIF�F�C��J#��G
Mv��OL�ENDǪ�LU��CPR��L�u�S�C$�StT�E�S60�FVmRV�IN��IH�� �m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s�������軏͏ߏ�S�TD�LANG���0�B�T�f� x���������ҟ��� ��,�>�P�b�t��� ������ί���� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢϴ��� ������� �2�D�V��h�zߌߞ߰���RB=T
�OPTN���� ��'�9�K�]�o�������������DPN	���)�;�M�_� q��������������� %7I[m �������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu���� �����)�;�M� _�q���������ˏݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+�=� O�a�sυϗϩϻ��� ������'�9�K�]� o߁ߓߥ߷������� ���#�5�G�Y�k�}� ������������� �1�C�U�g�y����� ����������	-?Qc�f�������99���$FEAT_AD�D ?	����  	�#5GYk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ���������DEM�O y   �L�B�T߁� xߊ߷߮��������� ��G�>�P�}�t�� ������������ C�:�L�y�p������� ��������?6 Hul~���� ��;2Dq hz������  /
/7/./@/m/d/v/ �/�/�/�/�/�/�/? 3?*?<?i?`?r?�?�? �?�?�?�?�?O/O&O 8OeO\OnO�O�O�O�O �O�O�O�O+_"_4_a_ X_j_�_�_�_�_�_�_ �_�_'oo0o]oTofo �o�o�o�o�o�o�o�o #,YPb�� �������� (�U�L�^��������� ��ʏ����$�Q� H�Z���~�������Ɵ ����� �M�D�V� ��z�������¯ܯ� �
��I�@�R��v� ��������ؿ��� �E�<�N�{�rτϱ� �Ϻ��������A� 8�J�w�n߀߭ߤ߶� ��������=�4�F� s�j�|�������� ����9�0�B�o�f� x��������������� 5,>kbt� ������1 (:g^p��� ���� /-/$/6/ c/Z/l/�/�/�/�/�/ �/�/�/)? ?2?_?V? h?�?�?�?�?�?�?�? �?%OO.O[OROdO�O �O�O�O�O�O�O�O!_ _*_W_N_`_�_�_�_ �_�_�_�_�_oo&o SoJo\o�o�o�o�o�o �o�o�o"OF X�|����� ����K�B�T��� x�������ۏҏ�� ��G�>�P�}�t��� ����ןΟ����� C�:�L�y�p������� ӯʯܯ	� ��?�6� H�u�l�~�����Ͽƿ ؿ����;�2�D�q� h�zϔϞ�������� ��
�7�.�@�m�d�v� �ߚ��߾�������� 3�*�<�i�`�r��� ����������/�&� 8�e�\�n��������� ��������+"4a Xj������ ��'0]Tf �������� #//,/Y/P/b/|/�/ �/�/�/�/�/�/?? (?U?L?^?x?�?�?�? �?�?�?�?OO$OQO HOZOtO~O�O�O�O�O �O�O__ _M_D_V_ p_z_�_�_�_�_�_�_ o
ooIo@oRolovo �o�o�o�o�o�o E<Nhr�� �������A� 8�J�d�n�������я ȏڏ����=�4�F� `�j�������͟ğ֟ ����9�0�B�\�f� ������ɯ��ү���� �5�,�>�X�b����� ��ſ��ο����1� (�:�T�^ϋςϔ��� �������� �-�$�6� P�Z߇�~ߐ߽ߴ��� ������)� �2�L�V� ��z���������� ��%��.�H�R��v� ��������������! *DN{r�� �����& @Jwn���� ���//"/</F/ s/j/|/�/�/�/�/�/ �/???8?B?o?f? x?�?�?�?�?�?�?O OO4O>OkObOtO�O �O�O�O�O�O__0]  'XF_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX j|������ ���0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ����������
��.�   /�)�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ����� ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�� ������������ &�8�J�\�n������� ����������"4 FXj|���� ���0BT fx������ �//,/>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodo vo�o�o�o�o�o�o�o *<N`r� �������� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$�
4�8�+�N�`�r� �ߖߨߺ�������� �&�8�J�\�n��� ������������"� 4�F�X�j�|������� ��������0B Tfx����� ��,>Pb t������� //(/:/L/^/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�? �?�?�?�?�?O O2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�o�o�o�o�o�o &8J\n�� �������"� 4�F�X�j�|������� ď֏�����0�B� T�f�x���������ҟ �����,�>�P�b� t���������ί�� ��(�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢ� ����������� �2� D�V�h�zߌߞ߰��� ������
��.�@�R� d�v��������� ����*�<�N�`�r� �������������� &8J\n�� ������" 4FXj|��� ����//0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O �O�O�O�O�O�O __�$_6Y�$FEAT�_DEMOIN [ ;T�fP�<P}NTINDEX[[�jQ�NPILEC�OMP z�;���QiRIU��PSETUP2 �{�U�R��  N �Q�S_A�P2BCK 1|~�Y  �)7XDok%�_8o<P�P &oco9U�_�oo�oBo �o�oxo�o1C�o g�o��,�P� ����?��L�u� ���(���Ϗ^�󏂏 �)���M�܏q���� ��6�˟Z�؟���%� ��I�[�������� D�ٯh������3�¯ W��d������@�տ �v�Ϛ�/�A�пe� ���ϛ�*Ͽ�N���r� ��ߨ�=���a�s�� ��&߻���\��߀�� '��K���o���|�� 4���X������#��� G�Y���}������B� ��f�����1�Y�P�P�_ 2�P*�.VR8���*��������l P�C���FR6�:�2�V�T zPz�w�]PG<���*.Fo/"��	�:,�^/�STMi/�/ D/�-M/�/�H�/�?�'?�/�/g?�GIFq?�?�%�?D?V?�?�JPG�?O�%`O�?�?oO�
JSyOĢO��5C�OMO%
�JavaScri3pt�O�?CS�O&_��&_�O %Ca�scading �Style Sh�eetsR_��
A�RGNAME.D)T�_��� \�_S_еA�T�_�_�PDI'SP*�_���To��_�QLaZooCLLB.ZIwo2o$ K:\�a\�o�i�ACollabo�o��o
TPEINS�.XML�_:\�![o�QCusto�m Toolba�rbiPASSW�ORDQo��FR�S:\�dB`Pa�ssword Config���/� �(�e�������� N��r�����=�̏ a������&���J��� 񟀟���9�K�ڟo� ������4�ɯX��|� ��#���G�֯@�}�� ��0�ſ׿f������ 1���U��y��ϯ� >���b���	ߘ�-߼� Q�c��χ�߽߫�L� ��p��ߦ�;���_� ��X��$��H����� ~����7�I���m��� �� �2���V���z��� !��E��i{
� .��d��� �S�wp�< �`�/�+/�O/ a/��//�/8/J/�/ n/?�/�/9?�/]?�/ �?�?"?�?F?�?�?|? O�?5O�?�?kO�?�O O�O�OTO�OxO__ �OC_�Og_y__�_,_ �_P_b_�_�_o�_o Qo�_uoo�o�o:o�o ^o�o�o)�oM�o �o��6��l ��%�7��[��� �� ���D�ُh�z�� ��3�,�i������ ��ßR��v�������$FILE_D�GBCK 1|������� < �)
�SUMMARY.�DG!�͜MD:�U���ِDia�g Summar�y����
CONSLOG��n���ٯ����Consol�e log���	?TPACCN�t��%\�����TP �Accounti�n;���FR6:�IPKDMP.ZIPͿј
�ϥ����Excepti�on"�ӻ��MEMCHECK���������-�Memor?y Data�����@n )��RI�PE�~ϐ�%ߴ��%�� Pack�et L:���L��$�c���STAT���߭� %�A�Status<��^�	FTP�����	��/�mme?nt TBD2�^�� >I)ETHERNEw�
�d�u���﨡Ether�nJ�1�figur�aAϩ��DCSV�RF&���7������ verify� all:��� {4��DIFF/���'���;�Q�dif�f��r�d���CHG01������A����,it�2���27@0���fx3�8��I �p��VTRNDIAG.LSu&8����� Ope���L� ��nost�ic��H�)�VDEV�DAT�������Vi�s�Device�+IMG��,/�>/�/:�i$Ima�gu/+UP E�S/�/FRS:�\?Z=��Upd�ates Lis�tZ?��� FLEXEVEN��/�/��?���1 UIF� EvM�M���-�vZ)CRSEONSPK�/˞�q\!O���CR_TAOR_PEAKbO�ͩPSRBWLD'.CM�O͜E2�O�\?.�PS_ROB�OWELS���:G�IG��@_�?d_���GigE�(O��Nߵ@�)UQHADOW__D_V_�_���Shadow ?Change�����2dt�RRCME�RR�_�_�_oo���4`CFG Err{oro tailo� MA�k�CMSGLIBgoNo`o`�o|R�e��z0ic�oޭa�)�`ZD�0_O�os��ZDf�Pad�l �RNOTI�Rd����Notifi�c����,�AG ��P�ӟt��������� Ώ]�����(���L� ^�폂������G�ܟ k� ����6�şZ�� ~������C�د�y� ���2�D�ӯh����� ���¿Q��u�
�� ��@�Ͽd�v�Ϛ�)� ����_��σ�ߧ�%� N���r�ߖߨ�7��� [�����&��J�\� �߀���3����i� ���"�4���X���|� �����A�����w� ��0��=f��� ��O�s� >�bt�'� K���/�:/L/ �p/��/�/5/�/Y/ �/ ?�/$?�/H?�/U? ~??�?1?�?�?g?�? �? O2O�?VO�?zO�O O�O?O�OcO�O
_�O ._�OR_d_�O�__�_ �_M_�_q_oo�_<o �_`o�_mo�o%o�oIo �o�oo�o8J�o n�o��3�W� {�"��F��j�|� ���/�ď֏e�������0��$FILE�_FRSPRT � �������?�MDONLY 1|S��� 
 �)�MD:_VDA�EXTP.ZZZ�1�⏹�ț6%�NO Back? file ���S�6P�����>� �K�t�����'���ί ]�򯁯�(���L�ۯ p������5�ʿY�׿  Ϗ�$ϳ�H�Z��~� Ϣϴ�C���g���� ��2���V���cߌ�� ��?�����u�
��.�@���d��߈��C�VISBCKq�[���*.VD����S��FR:\��ION\DATA\���v�S�Vision VD��� Y�k����y��B��� ��x���1C��g ���,�P�� ��?�Pu �(��^��/ ��M/�q/�/>/�/ 6/�/Z/�/?�/%?�/ I?[?�/??�?2?D?��?9�LUI_CONFIG }S�����; $ 	�3v�{S�;OMO_O`qO�O�O�I#@|x�? �O�O�O__%\�OH_ Z_l_~_�_'_�_�_�_ �_�_o�_2oDoVoho zo�o#o�o�o�o�o�o 
�o.@Rdv� ������� *�<�N�`�r������ ��̏ޏ�����&�8� J�\�n��������ȟ ڟ쟃���"�4�F�X� j��������į֯� ���0�B�T�f��� ��������ҿ�{�� �,�>�P�b����Ϙ� �ϼ�����w���(� :�L�^��ςߔߦ߸� ����s� ��$�6�H� ��Y�~������]� ����� �2�D���h� z���������Y����� 
.@��dv� ���U�� *<�`r��� �Q��//&/8/ �\/n/�/�/�/;/�/ �/�/�/?"?�/F?X? j?|?�?�?7?�?�?�? �?OO�?BOTOfOxO �O�O3O�O�O�O�O_ _�O>_P_b_t_�_�_ /_�_�_�_�_oo�_�:oLo^opo�o�o$h�  x�o�c�$�FLUI_DAT�A ~���>�a(a�d�RESULT 3��ep ��T�/wiza�rd/guide�d/steps/?Expert�o= Oas���������z�Con�tinue wi�th Gpance�:�L�^�p����������ʏ܏� � �b-�a�e�0� �0`��c�a?��ps������� ��ҟ�����,�>� P��0ow��������� ѯ�����+�=�O��a�?�1�C�U�e�cllbs�ֿ���� �0�B�T�f�xϊϜ� [�����������,� >�P�b�t߆ߘߪ�i��{��ߟ�]�e�rip(pſ-�?�Q�c�u� ������������ �)�;�M�_�q����� �����������������`�e�#pTi�meUS/DST 	��������!3E�Enabl(�y��� ����	//-/?/
Q/�b�)�/M_q24|�/�/? ?)?;?M?_?q?�?�? Tf�?�?�?OO%O 7OIO[OmOO�O�Ob/�t/�/�/Z�"qRegion�O5_G_Y_ k_}_�_�_�_�_�_�_��America!�#o5oGoYoko}o �o�o�o�o�o�o��A�y�O�O3�O_qEditor�o�� �������+��=� � Touch Panel rs� (recommenp�)K������� Ə؏���� �2�D�|�%��I[qaccesoܟ�  ��$�6�H�Z�l�~������Conne�ct to Network��֯� ����0�B�T�f�x�(����x��@��}�䏟�,!��s Int?roduct!_4� F�X�j�|ώϠϲ��� �������0�B�T� f�xߊߜ߮��������� ɿ��" �i�{�������� ������/�A� �e� w��������������� +=�H�3��+�O��� �� 2DVh z�K������ 
//./@/R/d/v/�/ �/Yk}�/�?? *?<?N?`?r?�?�?�? �?�?�?��?O&O8O JO\OnO�O�O�O�O�O �O�O�/_�/1_�/X_ j_|_�_�_�_�_�_�_ �_oo0oBoS_foxo �o�o�o�o�o�o�o ,>�O_!_�E_ �������(� :�L�^�p�����So�� ʏ܏� ��$�6�H� Z�l�~���O��s՟ ���� �2�D�V�h� z�������¯ԯ毥� 
��.�@�R�d�v��� ������п⿡��ş '�9���`�rτϖϨ� ����������&�8� ��\�n߀ߒߤ߶��� �������"�4��=� �a��Mϲ������� ����0�B�T�f�x� ��I߮��������� ,>Pbt�E� ��i����( :L^p���� ���� //$/6/H/ Z/l/~/�/�/�/�/�/ ����/?�V?h? z?�?�?�?�?�?�?�? 
OO.O�ROdOvO�O �O�O�O�O�O�O__ *_<_�/??�_C?�_ �_�_�_�_oo&o8o Jo\ono�o?O�o�o�o �o�o�o"4FX j|�M___q_��_ ���0�B�T�f�x� ��������ҏ�o�� �,�>�P�b�t����� ����Ο�����%� �L�^�p��������� ʯܯ� ��$�6�G� Z�l�~�������ƿؿ ���� �2��S�� w�9��ϰ��������� 
��.�@�R�d�v߈� G��߾��������� *�<�N�`�r��Cϥ� g���ύ���&�8� J�\�n����������� ������"4FX j|������� ���-��Tfx �������/ /,/��P/b/t/�/�/ �/�/�/�/�/??(? �1U??A�?�? �?�?�? OO$O6OHO ZOlO~O=/�O�O�O�O �O�O_ _2_D_V_h_ z_9?�?]?�_�_�?�_ 
oo.o@oRodovo�o �o�o�o�o�O�o *<N`r��� ���_�_�_�_#��_ J�\�n���������ȏ ڏ����"��oF�X� j�|�������ğ֟� ����0����u� 7�������ү���� �,�>�P�b�t�3��� ����ο����(� :�L�^�pς�A�S�e� �ω��� ��$�6�H� Z�l�~ߐߢߴ��߅� ����� �2�D�V�h� z����������� �����@�R�d�v��� ������������ *;�N`r��� ����&�� G	�k-����� ���/"/4/F/X/ j/|/;�/�/�/�/�/ �/??0?B?T?f?x? 7�?[�?�?�?O O,O>OPObOtO�O�O �O�O�O�/�O__(_ :_L_^_p_�_�_�_�_ �_�?�_�?o!o�OHo Zolo~o�o�o�o�o�o �o�o �ODVh z������� 
���_%o�_I�s�5o ������Џ���� *�<�N�`�r�1���� ��̟ޟ���&�8� J�\�n�-�w�Q���ů ������"�4�F�X� j�|�������Ŀ��� ����0�B�T�f�x� �ϜϮ���������� �ٯ>�P�b�t߆ߘ� �߼���������տ :�L�^�p����� ������ ��$����� �i�+ߐ��������� ���� 2DVh '������� 
.@Rdv5� G�Y��}���// */</N/`/r/�/�/�/ �/y�/�/??&?8? J?\?n?�?�?�?�?�? ��?�O�4OFOXO jO|O�O�O�O�O�O�O �O__/OB_T_f_x_ �_�_�_�_�_�_�_o o�?;o�?_o!O�o�o �o�o�o�o�o( :L^p/_��� ��� ��$�6�H� Z�l�+o��Oo��sou� ���� �2�D�V�h� z����������� 
��.�@�R�d�v��� ������}�߯���� ٟ<�N�`�r������� ��̿޿���ӟ8� J�\�nπϒϤ϶��� �������ϯ��=� g�)��ߠ߲������� ����0�B�T�f�%� ������������� �,�>�P�b�!�k�E� ����{�����( :L^p���� w��� $6H Zl~���s��� ����/��2/D/V/h/ z/�/�/�/�/�/�/�/ 
?�.?@?R?d?v?�? �?�?�?�?�?�?OO ���]O/�O�O�O �O�O�O�O__&_8_ J_\_?�_�_�_�_�_ �_�_�_o"o4oFoXo jo)O;OMO�oqO�o�o �o0BTfx ���m_���� �,�>�P�b�t����� ����{oݏ�o��o(� :�L�^�p��������� ʟܟ� ��#�6�H� Z�l�~�������Ưد ����͏/��S�� z�������¿Կ��� 
��.�@�R�d�#��� �ϬϾ��������� *�<�N�`����C��� g�i�������&�8� J�\�n�����u� �������"�4�F�X� j�|�������q����� ��	��0BTfx ������� ��,>Pbt�� �����/�� ��1/[/�/�/�/�/ �/�/�/ ??$?6?H? Z?~?�?�?�?�?�? �?�?O O2ODOVO/ _/9/�O�Oo/�O�O�O 
__._@_R_d_v_�_ �_�_k?�_�_�_oo *o<oNo`oro�o�o�o gOyO�O�O�o�O&8 J\n����� ����_"�4�F�X� j�|�������ď֏� ����o�o�oQ�x� ��������ҟ���� �,�>�P��t����� ����ί����(� :�L�^��/�A���e� ʿܿ� ��$�6�H� Z�l�~ϐϢ�a����� ����� �2�D�V�h� zߌߞ߰�o��ߓ��� ���.�@�R�d�v�� ������������ *�<�N�`�r������� ����������#�� G	�n����� ���"4FX �|������ �//0/B/T/u/ 7�/[]/�/�/�/? ?,?>?P?b?t?�?�? �?i�?�?�?OO(O :OLO^OpO�O�O�Oe/ �O�/�O�O�?$_6_H_ Z_l_~_�_�_�_�_�_ �_�_�? o2oDoVoho zo�o�o�o�o�o�o�o �O_�O%O_v� �������� *�<�N�or������� ��̏ޏ����&�8� J�	S-w���cȟ ڟ����"�4�F�X� j�|�����_�į֯� ����0�B�T�f�x� ����[�m����󿵟 �,�>�P�b�tφϘ� �ϼ������ϱ��(� :�L�^�p߂ߔߦ߸� ������ ￿ѿ�E� �l�~�������� ����� �2�D��h� z��������������� 
.@R�#�5� �Y���� *<N`r��U� ����//&/8/ J/\/n/�/�/�/c�/ ��/�?"?4?F?X? j?|?�?�?�?�?�?�? �??O0OBOTOfOxO �O�O�O�O�O�O�O�/ _�/;_�/b_t_�_�_ �_�_�_�_�_oo(o :oLoOpo�o�o�o�o �o�o�o $6H _i+_�O_Q�� ��� �2�D�V�h� z�����]oԏ��� 
��.�@�R�d�v��� ��Y��}ߟ񟵏� *�<�N�`�r������� ��̯ޯ𯯏�&�8� J�\�n���������ȿ ڿ쿫���ϟ�C�� j�|ώϠϲ������� ����0�B��f�x� �ߜ߮���������� �,�>���G�!�k�� Wϼ���������(� :�L�^�p�����S߸� ������ $6H Zl~�O�a�s�� ��� 2DVh z�������� 
//./@/R/d/v/�/ �/�/�/�/�/�/�� �9?�`?r?�?�?�? �?�?�?�?OO&O8O �\OnO�O�O�O�O�O �O�O�O_"_4_F_? ?)?�_M?�_�_�_�_ �_oo0oBoTofoxo �oIO�o�o�o�o�o ,>Pbt�� W_�{_��_��(� :�L�^�p��������� ʏ܏���$�6�H� Z�l�~�������Ɵ؟ ꟩��/��V�h� z�������¯ԯ��� 
��.�@���d�v��� ������п����� *�<���]����C�E� ����������&�8� J�\�n߀ߒ�Q����� �������"�4�F�X� j�|��Mϯ�q����� ����0�B�T�f�x� �������������� ,>Pbt�� ���������� 7��^p���� ��� //$/6/�� Z/l/~/�/�/�/�/�/ �/�/? ?2?�; _?�?K�?�?�?�?�? 
OO.O@OROdOvO�O G/�O�O�O�O�O__ *_<_N_`_r_�_C?U? g?y?�_�?oo&o8o Jo\ono�o�o�o�o�o �o�O�o"4FX j|������ �_�_�_-��_T�f�x� ��������ҏ���� �,��oP�b�t����� ����Ο�����(� :�����A����� ʯܯ� ��$�6�H� Z�l�~�=�����ƿؿ ���� �2�D�V�h� zό�K���o��ϓ��� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� �����������#��� J�\�n����������� ������"4��X j|������ �0��Q�u 7�9�����/ /,/>/P/b/t/�/E �/�/�/�/�/??(? :?L?^?p?�?A�?e �?�?�/ OO$O6OHO ZOlO~O�O�O�O�O�O �/�O_ _2_D_V_h_ z_�_�_�_�_�_�?�? �?o+o�?Rodovo�o �o�o�o�o�o�o *�ON`r��� ������&��_ /o	oS�}�?o����ȏ ڏ����"�4�F�X� j�|�;����ğ֟� ����0�B�T�f�x� 7�I�[�m�ϯ����� �,�>�P�b�t����� ����ο�����(� :�L�^�pςϔϦϸ� ���ϛ�����!��H� Z�l�~ߐߢߴ����� ����� �߿D�V�h� z������������ 
��.������s�5� ������������ *<N`r1�� ����&8 J\n�?��c�� ����/"/4/F/X/ j/|/�/�/�/�/�/� �/??0?B?T?f?x? �?�?�?�?�?��?� O�>OPObOtO�O�O �O�O�O�O�O__(_ �/L_^_p_�_�_�_�_ �_�_�_ oo$o�?Eo Oio+O-o�o�o�o�o �o�o 2DVh z9_������ 
��.�@�R�d�v�5o ��Yo��͏���� *�<�N�`�r������� ��̟����&�8� J�\�n���������ȯ ��я������F�X� j�|�������Ŀֿ� ����ݟB�T�f�x� �ϜϮ���������� �ٯ#���G�q�3��� �߼���������(� :�L�^�p�/ϔ��� ������ ��$�6�H� Z�l�+�=�O�a����� ���� 2DVh z�������� 
.@Rdv� ����������/ ��</N/`/r/�/�/�/ �/�/�/�/??�8? J?\?n?�?�?�?�?�? �?�?�?O"O��/ gO)/�O�O�O�O�O�O �O__0_B_T_f_%? w_�_�_�_�_�_�_o o,o>oPoboto3O�o WO�o{O�o�o( :L^p���� ��o� ��$�6�H� Z�l�~�������Ə�o 珩o��o2�D�V�h� z�������ԟ��� 
���@�R�d�v��� ������Я����� ׏9���]��!����� ��̿޿���&�8� J�\�n�-��Ϥ϶��� �������"�4�F�X� j�)���M����߅��� ����0�B�T�f�x� ������������ �,�>�P�b�t����� ����{��ߟ����� :L^p���� ��� ��6H Zl~����� ��/����;/e/ '�/�/�/�/�/�/�/ 
??.?@?R?d?#�? �?�?�?�?�?�?OO *O<ONO`O/1/C/U/ �Oy/�O�O__&_8_ J_\_n_�_�_�_�_u? �_�_�_o"o4oFoXo jo|o�o�o�o�o�O�O �O	�O0BTfx �������� �_,�>�P�b�t����� ����Ώ������o �o�o[��������� ʟܟ� ��$�6�H� Z��k�������Ưد ���� �2�D�V�h� '���K���o�Կ��� 
��.�@�R�d�vψ� �ϬϾ�Ͽ������ *�<�N�`�r߄ߖߨ� ��y��ߝ�����&�8� J�\�n������� ���������4�F�X� j�|������������� ����-��Q� ������� ,>Pb!��� �����//(/ :/L/^//A�/�/ y�/�/ ??$?6?H? Z?l?~?�?�?�?s�? �?�?O O2ODOVOhO zO�O�O�Oo/�/�/�O _�/._@_R_d_v_�_ �_�_�_�_�_�_o�? *o<oNo`oro�o�o�o �o�o�o�o�O_�O /Y_����� ����"�4�F�X� o|�������ď֏� ����0�B�T�% 7I��mҟ���� �,�>�P�b�t����� ��i�ί����(� :�L�^�p��������� w���������$�6�H� Z�l�~ϐϢϴ����� ���ϻ� �2�D�V�h� zߌߞ߰��������� 
�ɿۿ�O��v�� ������������ *�<�N��_������� ��������&8 J\�}?�c�� ���"4FX j|������ �//0/B/T/f/x/ �/�/�/m�/��/� ?,?>?P?b?t?�?�? �?�?�?�?�?O�(O :OLO^OpO�O�O�O�O �O�O�O _�/!_�/E_ ?	_~_�_�_�_�_�_ �_�_o o2oDoVoO zo�o�o�o�o�o�o�o 
.@R_s5_ ��mo����� *�<�N�`�r������� gȍޏ����&�8� J�\�n�������c� �џ���"�4�F�X� j�|�������į֯� �����0�B�T�f�x� ��������ҿ����� ��ٟ#�M��tφϘ� �ϼ���������(� :�L��p߂ߔߦ߸� ������ ��$�6�H� ��+�=ϟ�a����� ����� �2�D�V�h� z�����]��������� 
.@Rdv����k�}������$FMR2_GR�P 1���� �C4�  B��	 ��9K6F@� a@�6G� � �Fg�fC��8R�y?�  x��66�X����875t��5���5`+�y�A�  /+BHx�w-%@S339%B�5[/l-6@6! �/xl/�/�/�/�/? �/&??J?5?G?�?k?��?��_CFG �TK�?�? O|O�9NO /
F0FA K@�<�RM_CHKTYP  ��$&�� ROMa@_MsINg@�����@u�R XSSB�3��� 7�O���C�O�O�5�TP_DEF_O/W  ��$W�IRCOMf@_��$GENOVRD�_DO�F��E]TYH��D dbUdKTo_ENB7_ KP�RAVC��G�@ �Y�O�_�?�oyo&oI* ��QOU��NAIRI< �@��oGo�o�o�o��C�p3��O:��B�+sL�i\�O�PSMT��Y�(�@
t�$HOS�TC�21��@s�5 MC���R{��� _ 27.00�1�  e�]�o��� ����K�ď֏���������	anonymous!�O�a�s�D���� �4���� ����D�!�3�E�W� i���������ï柀� .���/�A�S���� ��П����Ŀ��� �+�r�O�a�sυϗ� ����������'� n��������ϓ�ڿ�� ��������F�#�5�G� Y�k���υ������ ����B�T�f�C�z�g� �ߋ������������ 	-P�����u� �����(�:�< )p�M_q���� ����/$Zl I/[/m//�/��� �//�/D!?3?E?W? /?�?�?�?�?�/�? ./OO/OAOSO�/�/ �/�/�?�O?�O�O_ _+_r?O_a_s_�_�_ �O�?O�_�_oo'o��t�qENT 1��hk P!�_no  �p\o�o�o�o �o�o�o�o�o: _"�F�j�� ���%��I��m� 0���T�f�Ǐ��돮� �ҏ3���,�i�X��� P���t�՟��៼�
� /��S��w�:���^� �����������ܯ=�� �QUICC0�J�&�!192.�168.1.10c�X�1��v�8��\��2�ƿؿ9�!R�OUTER:��!���a��PCJ�OG��e�!*� ��0��U�CAMgPRT�϶�!�����RTS���x�� !Softw�are Oper�ator Pan�elU߇���7kNA�ME !Kj!�ROBO����S_�CFG 1�Ki� �Au�to-start{ed�DFTP�Oa�O�_���O���� ������E_�.�@�R� u�c�	����������� cN:�L�^�;r���R �������� %H�[m� ��jO|O�O�O4!/ hE/W/i/{/�/T�/ �/�/�/�//�//?A? S?e?w?�?����? ?�?</O+O=OOO? sO�O�O�O�O�?`O�O __'_9_K_�?�?�? �?�O�_�?�_�_�_o #o�OGoYoko}o�o�_ 4o�o�o�o�of_ x_�_g�o��_�� ���o��-�?�Q� tu��������Ϗ� (:L^`�2��q� ����������ݟ�� �%�H�ʟ[�m���� ������� �ί4�!� h�E�W�i�{���T��� ÿտ�
�Ϟ�/�A��S�e�w����_ER�R ��ڇϗ�P�DUSIZ  j�^6����>��?WRD ?(�����  guest���+��=�O�a���SCD_�GROUP 3��(� ,�"�IF�T��$PA��OM�P�� ��_S�H��ED�� $C��COM��TTP�_AUTH 1���� <!iPendanm�x�#��+!KAREL�:*x���KC������VISION SET��@(����?�-�W�R� ��v������������������G�CTRL K���a�
��FFF9E3���FRS:D�EFAULT��FANUC W�eb Server�
tdG����/�� 2DV��W�R_CONFIGw ���������IDL_C_PU_PC� �sB���� BH��MIN����GNR_IO���������HMI_EDI�T ���
 ($/C/��2/k/V/�/ z/�/�/�/�/�/?�/ 1??U?@?y?d?�?�? ./�?�?�?�?OO?O QO<OuO`O�O�O�O�O��O�O�O__;_�N�PT_SIM_D�O�*NSTA�L_SCRN� ��\UQTPMOD�NTOL�Wl[�R�TYbX�qV�K�E�NB�W�ӭOL_NK 1����� o%o7oIo[omoo�R_MASTE��Y�%OSLAVE ���ϮeRAMCOACHE�o�ROM�O_CFG�o�S�c�UO'��bCMT�_OP�  "��5sY�CL�ou� _AS�G 1����
 �o������ �"�4�F�X�j�|���\�kwrNUM�����
�bIP�o�gRTRY_CN@uQO_UPD��a���1 �bp�b��n��hM��аP}T?��k ��._������ ɟ۟퟈S���)�;� M�_�q� �������˯ ݯ�~��%�7�I�[� m��������ǿٿ� ����!�3�E�W�i�{� 
ϟϱ��������ψ� ��/�A�S�e�w߉�� �߿���������+� =�O�a�s���&�� ����������9�K� ]�o�����"������� ��������GYk }��0���� �CUgy� �,>���	// -/�Q/c/u/�/�/�/ :/�/�/�/??)?�/ �/_?q?�?�?�?�?H? �?�?OO%O7O�?[O mOO�O�O�ODOVO�O �O_!_3_E_�Oi_{_ �_�_�_�_R_�_�_o o/oAo�_�_wo�o�o �o�o�o`o�o+ =O�os���� �\n��'�9�K� ]����������ɏۏ�i�c�_MEMBE�RS 2�:�   $:� ���v����1���RCA_AC�C 2���   [~�� c�v ��p .4 6��l�l�l����� ����  ��� a�BUF0�01 2�n�= ���u0  uW0�����������"�"��@�@������[����u�0��R�R�$�R�2u0m����BR�OR�]R�l�u0�]H�y�u0G�-`��V�����������U���ʢ�ע�梤R!������U'�4�C�P⤀��䢑�䢙�䢡��U�⤤⤱���U��������U��!�.�U;�K�X�g�Ut�������	��ߙ2����� �����!��(� -�1�-�9�:�@��H� M�Q�c�]�y���]� ]¡�]©�]±�]¹� ]���]�ɠ]�Ѡ]�٠ ]�*����������� ���	��������� ��(��¢�8���A��� I���Q���Y���a��� i���q���y��� ����¡�� ��±�¹����� ɰ�Ѱ�ٰ���ߙ3�������� �!�/�6�1�?�l�@� O�N�Z�l�a�f�j�f� i�f�q�f��f��f� !���f�1���f⩢�� f⹢��f�ɢ��f�٢ ��l����������� 	�����'����0� ?���A�O���Q�_��� a�o���q��⁲�� ⑲��⡲��Ⱳ ��������Ѳ�������CFG 2�n� 4l��
l�J��<l�47���HIS钜n� ��� 2025�-11-3�l��    #� &f  '� "珪�  PTl�7 X�`�hl�z�pl�$  x��� 8 ��;  ��   7 9���
 2F$�6[}�Rq29 }	7v����������  � % � � � -�R  *$� l��B��aN/ `/r/�/�/�/�/�/�/ �/'/9/&?8?J?\?n? �?�?�?�?�?�/?�? O"O4OFOXOjO|O�O �O�?�?�O�O�O__ 0_B_T_f_x_�O�O�O �_�_�_�_oo,o>o�Po�O��[m
8
 c� 8���o�o�6d� �b� �b� _+  X�  �X�  d��!qc
	,: J!r���b �oWEW���� �����:�a �2�a ,*q 1  \�_�_m���� ����Ǐُ�����_ X�E�W�i�{������� ß՟��0���/�A� S�e�w����������� ����+�=�O�a� s���������߿� ��'�9�K�]�oρ� J�Ѐo�o

eq� ��������� �� � ��� ��� eq� �Geq	$">� 	�x�fx�� ����������,���� �� Z� �� ��п���������� ��&�8�o��n��� �������������� G�Y�FXj|�� ����1�0 BTfx���� �	//,/>/P/�b/t/�/�/�Ϙ�I_�CFG 2���� H
Cycl�e Time��Busy�Idyl�"�min�+=1Up�&��Read�'�Dow8?�` 1��#Count�	ONum �"����<��b�qaPROmG�"�������)/softp�art/genl�ink?curr�ent=menu�page,1133,1�/OO/OAO�3b5leSDT_ISOLC  ����p�/J23_DSP_ENBL��vK0�@INC �M�ӄ@A   �?&p=���<#��
�A�I:�o����N_���O<_�GOB�0C�CF�1�FVQ�G_GROUP �1�vK	r<A��C�٢_D_?���?�_��Q�_o.o�@o�_dovo�o�o���,_NYG_IN_A�UTODԫMPOS�RE^_pVKANJ?I_MASK v�H�qRELMON #��˔?��y_ox������.6r�3��7�C���u�o�D�KCL_L�`NU�ML��EYLOGOGINGDЫ���Q��E�0LANGUA_GE ��~���DEFAUgLT ����LG�!���:2�?��W�80H  ����'��  � 
���ћ��GOUF �;��
��(U�T1:\��   �-�?�Q�h�u�����@����ϟ�����(g�4�8i�N_DISP ��O8�_�_~��LOCTOL�����Dz`�A�A��GBOOK ���Ad�1
�
�۠#� ����#�5�G�Y�i�0��3{�W�	��쉠�QQJ¿Կ1��_BUFF 2�vK' ���25
��ڢVB&�7 Co�llaborativ�=�OΗώϠ� ����������'��0߀]�T�fߓߊߜ��DCS ��9�B�A x���Rh�%�-�?�Q���IO 2���c ���Q�� ������������ *�<�N�b�r������� ��������&:~e�ER_ITMsNd�o������ �#5GYk} ���������NhSEV�`�MdTYPsN�c/u/8�/
-�aRST5����SCRN_FL +2�s��0����/�??1?C?U?g?�/T�PK�sOR"��NG�NAM�D��~�N�U?PS_ACR� ^�4DIGI�8+)�U_LOAD[PG� %�:%T_?NOVICEt?���MAXUALRMX2��a���E
ZB&�1_P�5�` ��y�Z@CY��˭�O+����ۡ�D|PP 2�.˫ �Uf	R/_ 
_C_._g_y_\_�_�_ �_�_�_�_�_oo?o Qo4ouo`o�o|o�o�o �o�o�o)M8 qTf����� ��%��I�,�>�� j�����Ǐُ����� !���W�B�{�f��� ����՟����ܟ�/� �S�>�w���l����� ѯ��Ư��+��O��a�D���p���RHDBGDEF ��E��ѱO��_LDXD�ISA�0�;c�ME�MO_AP�0E {?�;
 ױ ��3�E�W�i�{ύϟ����Z@FRQ_CF�G ��G۳AM ��@��Ô�<�ԃd%�� ������B��K���*i�/k� **: tҔ�g�y�ߔ��߱� ���������J �Es�J d�����,(H���[����� @�'�Q�v�]������� ��������*N~PJISC 1��9Z� ������ܿ������	Zl_M?STR �#-,�SCD 1�"͠ {������ ��//A/,/e/P/ �/t/�/�/�/�/�/? �/+??O?:?L?�?p? �?�?�?�?�?�?O'O OKO6OoOZO�O~O�O �O�O�O�O_�O5_ _ Y_D_i_�_z_�_�_�_ �_�_�_o
ooUo@o yodo�o�o�o�o�o�o �o?*cN�6MK���;���$MLTARM����N��r ���հ��İME�TPU��zr���CNDSP_AD�COL%�ٰ0�CM�NTF� 9�FN�b�f�7�FSTLI8��x�4 �;ڎ��s����9�POS�CF��q�PRP�Me��STD�1��; 4�#�
 v��qv�����r����� ���̟ޟ ���V� 8�J���n���¯��������9�SING_�CHK  ��$oMODA���t��{�~2�DEV }	�	MC:f��HSIZE��zp��2�TASK %��%$123456789 ӿ�0�TRIG 1�; lĵ�2ϻ�!�bϻ�YP����H��1�EM_INF� 1�N�`)�AT&FV0E�0g���)��E0�V1&A3&B1�&D2&S0&C�1S0=��)A#TZ��2��H6�^���Rφ��A�߶�q�������� ��5��� ���ߏ�B߳����� ������1�C�*�g� �,��P�b�t����� ��R�?���u0 ����������� ����M q��� Z���/�%/� �[/ 2�/�/h �//�/�/�3?�/W? >?{?�?@/�?d/v/�/ �/O�//OAOx?eO?��ODO�O�O�O�O_�N�ITORÀG ?�z�   	EOXEC1~s&R2,X3,X4,X5,X��.VU7,X8,X9~s'R �2�T+R�T7R�TCR�T OR�T[R�TgR�TsR�TPR�T�R�S2�X2�XU2�X2�X2�X2�XU2�X2�X2�X2h�3�X3�X37R2�R�_GRP_SV �1��� (�>��:8>�s����=Z�׿2n?��a�ƽ�_D�B���cIO/N_DB<��@�zq  �����1tk�$��>w�zp�zp Y��@Nep7U�rp�>{ Mp Qu? -ud1������8�PG_JOOG �ʏ�{
�}2�:�o�?=���?�����0�B��~\�n���������H�?��C�@�Qqȏڏ���  ������qL_NA_ME !ĵ8���!Defau�lt Perso�nality (�from FD)�eq1�RMK_EN�ONLY�_�R2��a 1�L�X�L�8�gpl d����şן��� ��1�C�U�g�y��� ������ӯ���	�� ��
�<�N�`�r�����ਿ��̿޿�  :��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+��<�S ew����������A�a���B�Bw��P f������/ !/3/E/W/i/{/�/�/ �/���/�/??/? A?S?e?w?�?�?�?�? �?�?�?�/�/+O=OOO aOsO�O�O�O�O�O�O �O__'_9_&O�SB���`z_�[7rdtS ���_�]�_�_�W������S"oe_oXoa ��qogoyo�o�o�o��o�ouP�p"|����	`[oUgy8q�K�A\����s� �A��y@h�Q�Qʿ�"���Tk\~$��  ��P��PE�xC�  �I�@oa�<o��p� ������ߏ
f�Q*��҈��0��PCr� � 3r �.�� @D�  A�?��G�-�?.I�.@�I�A����  �;�	lY�	 ��X  ������� �, � ������uPK�o������]K��K]��K	�.���w�r_	����@
��)�b�1�����I��Y�����T�;fY�{S���'3����I�>J����;Î?v�>��==@�����E��RѯעZ���wp��u��� D!�3���7pg  � � �9�͏W���	�'� � u��I� �  y��u��:�È��?È=��ͱ���@��ǰ�3��D\�3�E�&���N�pC�  'Y�&�Z��i�b�@f�i�n�C�����I�C����&b��r�� p����B�p�Ŕq���}ر�.DzƏ<ߛ��`�K�pߖ���������А� 4P����.z���d  �Pؠ?�ff�_��	� 2p>�P���8.f�t�>L���U���(.��P�����ð��
ĉ��� x��;�e�m��KZ;��=g;�4�<�<����%�G���3����p?fff�?ذ?&S���@{=0e�?��q� +�rN�Z���I���G� ��7���(�����! E0iT����+��F�p��� #��D��w� ������// =/(/a/L/�/p/��/ �p�6�/Z#?�/ ? Y?k?}?��?�?>?�?��?�?�?�?1O�����KD�y^KCO�OO�O���ذO�O�O�Oai���J��}�D#D1���.�D��@�A�mQa��9N,ȴA�;�^@��T@�|j@$�?��V�>�z������=#�
>�\)?��
=��G�-]�{�=���,��C+��Bp���P���6��C98R����?N@���(��5-]G��p�Gsb�F��}�G�>.E�VD�Kn����I�� F��W�E��'E���D��;n����I��`E��G��cE�vmD���-_ �oQ_�o�o�o �o$ H3X~i�� �������D� /�h�S���w������� �я
���.��R�=� v�a�s�����П���� ߟ��(�N�9�r�]� ��������ޯɯۯ� ��8�#�\�G���k��� ����ڿſ���"�� F�1�C�|�gϠϋ���@����������P(�Q�34�] ������Q�	�9�Oߵ53~�qmm��aҀ5Q����aғ����ߵ1�������1��U�C�y�g��%P�P���!�/��'���
�x��.������4� ;�t�_����������� ����:%��/0�/d����� ���7%[@Im���027�  B�S@J@�KCH#PzS@�0@ZO /1/C/U/g/y/�-�#��/�/�/�/�/�3�?�3�� @�3J��0�0�13��5
 ?f?x? �?�?�?�?�?�?�?O�O,O>OPO�Z@1 ����ۯ�c/�$�MR_CABLE� 2ƕ� ��TT�����ڰO ���O�)�@���C_�� ��_O_u_7_I__�_ �_�_�_�_o�_�_o Koqo3oEo{o�o�o�o �o�o�o�o�oGm /�K!�"���O� ���ذ�$�6���w*Y�** �C�OM ȖI����œ � c��%% 2345?678901����! ��Ï��� � !5� �!
���M�not segnt b��W���TESTFE�CSALGR  eg�*!d[�41�Y
k�������$�pB���������� 9�UD1:\ma�intenanc?es.xmlğ��  C:�D?EFAULT�,�B�GRP 2�z� � �� ��% � �%!1st �cleaning� of cont�. v�ilat�ion 56���B��!0�����+B���*�����+��"%���mech��c�al check^1�  �k�0u�|��ԯ����Ϳ�߿�@���rollCerS�e�w�ū���m�ϑϣϵ�@�B�asic qua?rterly�*�<�ƪ,\�)�;�M�_ߌq�8�MJ��ߓ "�8��� ���ߕ� �����+�=��C �g�ߋ�ʦ�߹���������@�Ov�erhau�ߔ��?� x� I�P����}���������� $n�������)l�A Sew������  �+=O� s������� /R�9/�(/��/ �/�/�/�//�/�/N/ #?r/G?Y?k?}?�?�/ �???�?8?OO1O COUO�?yO�?�?�O�? �O�O�O	__jO?_�O �Ou_�O�_�_�_�_�_ 0_oT_f_;o�__oqo �o�o�o�_�oo,o Po%7I[m�o� �o�o����!� 3��W�������� ÏՏ�6����l�� ��e�w���������џ �2��V�+�=�O�a� s������ͯ�� ��'�9���]����� ��⯷�ɿۿ���N� #�r���YϨ�}Ϗϡ� �������8�J��n� C�U�g�yߋ��ϯ��� ���4�	��-�?�Q� ��u������ߞ����� ����f�;����� ������������� P���t�I[m� �����:! 3EW�{���  ���//lA/ ��w/��/�/�/�/8�/X*�"	 X�/?.?@?�)B a/o?m/ o%w?�?�?}?�?�?O O�?�?OOaOsO1OCO �O�O�O�O�O__'_ �O�O]_o_�_?_Q_�_��_�_�_�_�\ о�!?�  @�! M?HoZolo�&4op�o�o�o�(*�o** F�@ �Q �V�`o'9�o]8o�����/^& �o�����/�A� S�e���#�����я �����+�q����� 7�������k�͟ߟ� �I�[���K�]�o����C�����ɯ��o$��!�$MR_HI_ST 2��U#��� 
 \7"$ �23456789C013�;���b2�90/����[���./� ���ǿٿF�X�j�!� 3ρϲ���{��ϟ�� ���B���f�x�/ߜ� S����߉��߭��,� ��P��t��=��$��SKCFMAPw  �U&�)�b
�� �����ONREL  ��$#������EXC/FENB�
�����&�FNC-��JO�GOVLIM�d�#�v���KEY�zy���_PAN�������RUNi��y���SFSPD�TYPM����SI�GN��T1MO�Tk����_CE_GRP 1��U��+�0�ow�# d����� �&�6\�7 y�m���/� 4/F/-/j/!/t/�/�/ �/{/�/�/�/?�+��QZ_EDIT
�����TCOM_C_FG 1���0��}?�?�? 
^1SI' �N����?��?���?$O�����?XO78T_ARC�_*�X�T_M�N_MODE
=�U:_SPL{O;�UAP_CPL�O�<�NOCHECK� ?�� �� _#_5_G_Y_k_ }_�_�_�_�_�_�_�_�oo��NO_WA�IT_L	S7> N�Tf1����%���qa_ERRH2�������?o�o�o�oB��OGj�@O�c}Ӧm| c�vGA�A���Aԫ���g2�@C�0����B�J�2��<���?����)��n�bPARAuM�b����t�GO�8
�.�@� = n�]�o�w�Q��� ��������Ϗ�)��7�[�m� ���~��ODRDSP�C�8�OFFSET�_CARI0�OǖDsISԟœS_A�@�ARK
T9OPE?N_FILE���1T6�0OPTIO�N_IO����K�M_PRG %���%$*����'�WO���Ns8�ǥ�� ��ur����	 �����Ӧ�����RG�_DSBL  �����jN���RI_ENTTO���C�����A ��U^�@IM_DS����r��V��LCT �{mP2ڢ�3̹��ydҩ��_PEX�@����RAT�G d�8��̐UP )װ�:����S�e�XKωϗ��$�r2G��L�XLȚ�l㰂��� ����'�9�K�]�o� �ߓߥ߷��������� �#�5�G���2��v� �������������e�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?�q 1�~?�?�?�?�?�?�?��?O O2ODO�yA�a�tn?~M��~O�O�P�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�O�Oo$o6o HoZolo~o�o�o�o�o �o�o�o �_oV hz������ �
��.�@�R�d�QO�ES������B�d�ӏ�ʏ����@����Y�D�}�0�� r���������ԟڟ��@�p���=�M��q��	`��������c�:�o�¯ԯ���>�A�  �k�TC�C�ڰ"ڰ����O��  ����-���)�C�  �t�k��� g�����Կ��ѿ
�5����_:�ĳ�OU����3��3�H���n�� �� ^�\� @oD�  p�?�v�b\�?:px�:qC4r��p�(��  ;�	�l��	 �X  ������� �,� � �������H�ʪ����H����Hw�zH���ϝ�8�<B���B�  Xѐ�x`�o�*��3����t�>u���fC{ߍ���:pB\�
�Ѵ=9:qK�t�� ����$���*���� DP�^���b�g  � � �h�����)�	�'� � ���I� �  y��'�=�������t�@����!�b��^;b�t�U�(�yN��r�  '��"E�C�И�t�C�И�`�ߗ���jA�@�����%�B�� ��,0���H:qDz�k��ߏz���݀������ 4P���:u�z:���	f��?�ff'�&8�� ]�m�8:p��>L�����$�(:p�P��	��`����:� x��;e�m"�KZ�;�=g;�4�<<���E/Tv���b���?ff�f?�?&� )�@�=0�%?�� �%_9��}!��$�x��/ v��/f'��W,??P? ;?t?_?�?�?�?�?�? �?O�?(OOLO�/�/ �/EO�OAO�O�O�O�O _�O_H_3_l_W_�_ {_�_�_1��_A���eO +o�ORooOo�o�o�o K/�o�omo�o*'`+�,�zt����CL�H��}?Ƀ����
�������u����D1��/n�t��p�q��@�I�h~,ȴA�;�^@��T@�|j@$�?��V�n�z������=#�
>�\)?��
=��G����{�=��,��C+��Bp�����6��C98R����?}p���(��5��G��p�Gsb�F��}�G�>.E�VD�KL�����I�� F��W�E��'E���D��;L�����I��`E��G��cE�vmD���\� ՟��ҟ���/��S� >�w�b�������ѯ�� �����=�(�:�s� ^���������߿ʿ� � �9�$�]�Hρ�l� �ϐϢ���������#� �G�2�W�}�hߡߌ� �߰��������
�C� .�g�R��v���� ����	���-��Q�<� u�`�r�����������@��'M�(��34�]O!����8h~�%3~�qm����5Q�������!���  `N��r��	eP@"P��Q�_/V/9/x$/]/H)����c/ j/�/�/�/�/�/�/�/ !??E?0?i?T?"&�_0�_�?�?�8��?�? O�?OBO0OfOTO�O@xO�O�O�O�O2f?_  B��pyp$QKCHR�z�p@� N_`_r_�_�_�_�]c�O�_�_oo+o�?�Bc� @Jd4�QJc�D
 2o�o�o �o�o�o�o%7�I[m��oa ������c/�$�PARAM_ME�NU ? ��  �DEFPULS�E��	WAIT�TMOUT�{R�CV� SH�ELL_WRK.�$CUR_STY�L�p"�OPT�8Q8�PTBM�G�C��R_DECSN �p������������ ��-�(�:�L�u�p���������qSSREL_ID  ���̕USE_P�ROG %�z%8���͓CCR�pޒ���s1�_HOST7 !�z!6�s��+�T�=���V�h����˯*�_TIME��rޖF��pGDE�BUGܐ�{͓GI�NP_FLMSK���#�TR2�#�PG�AP� ��_b�CyH1�"�TYPE�|�P������� �0�Y�T�f�xϡϜ� �����������1�,� >�P�y�t߆ߘ��߼� ����	���(�Q�L��^�p��%�WORD� ?	�{
 	�PR�p#MA9I��q"SUd���cTE��p#��	1���COLn%��!����L�� !���F�d�TRACE�CTL 1� ��q � #����_�_DT Q� ���z�D � ��ba��_`�� ����������1`CUgy�z t����� ,>Pbt��� ����//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�U��oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�.�o P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv���� ���*<N `r������ �//&/8/J/\/n/ Dϒ/�/�/�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z�����������$PGTR�ACELEN  ���  ������Ά_U�P ����2������΁_CFG ���S烸�
���*��:�D�O���O� � �O��DEF�SPD ��췁���΀H_C�ONFIG �\��� ����5dĔ�݂ ��ǑaP^�a�㑹��΀�IN�TRL ���=�8^���PEv��೗���p*�ÑO�΀LID����	T�LLB �1ⳙ ���BӐB4��O�� 䘼����Q�� << ��?�������M�3� U���i���������ӿ ��	�7�T�Ϣk� b�tϡ�诚���������S�GRP 1�������@A!�ߚ�4I���A ��Cu�C��OCjVF�/��Ȕa�zي�ÑÐ��t��ޯs������ӿߨ�B������������A�S�&�B34�_�������j������ ���	�B�-���Q����M�������  Dz ����.�����&L 7p[���� ���6!Zh�)w
V7.1�0beta1*��Ɛ@�*�@��) @�+A �Ē?��
?f�ff>����B_33A�Q�0��B(��A���AK��h���@�//'/9/P�p*��W�ӑ�n/�/�%����R�fh����*���P2�L R��/�/�/�/�/H?�Ĕ�I�u�&:�� �?��x?�?A���P!6\3 Bu�B��?�5SBH�3[4��o�L�4��[45��/B
\3x3Dx�?YO�?aOkO}O�<<�R@��O �C�O�O�O�O�DA�X��KNOW_M  �Z�%�X�SV 賚ڒ���_ �_�_?�_�_�_o��Ԃ�W�M+�鳛 ���	@�3#����_�o�\A��o
]bV4�@u���u��e�o�l,�X�MR+��JmT3?��W��1C{�OADBA�NFWDL_V�ST^+�1 1����P4C���[��i/ �����?�1�C� ��g�y��������ӏ �*�	��`�?�Q�c�w2�|Va�up�<ʟ���p3��Ɵ؟Ꟃw4��+�=��wA5Z�l�~����w6����ѯ㯂w7 ��$�6��w8S�e�w����w+MAmp������OVLD  ���yo߄rPARNUM  �{+þ��?υqSCH�� ��
��X���{s��U�PDX�)ź��Ϧ�_CMP_@`���p|P�'yu�ER_C;HK���yqbb3��.�RSpp?Q'_MOm��_}ߥ��_RES_G�p���
�e�����0�#� T�G�x�k�}��������������׳��� ������:�Y�^��� Y�y������Ӭ����� ����������R� 6UZ�ӥ�u����V 1�FvpVa�@k�p��THR_INRp��(bzyudMASS� Z)MNGM�ON_QUEUE� �uyvup\!*��N�UZ�NW���END��߶EcXE����BE�|��OPTIO���ۚPROGRAoM %z%���~ϘTASK_�I��.OCFG ��z+�n/� DAkTACc�+�0�;�up! 2 �??/?A?S?]51 s?�?�?�?�? �6p1�?�?�?O"O,F^�!INFOCc��-��bdlO~O�O�O�O �O�O�O�O_ _2_D_ V_h_z_�_�_�_�_�_h�/A@FD��, 	�l�!��K_�!�)fN!fENB��0m���Pf2YokhG�!2��0k X,		�d�=��·o���e�a$�pd��i�i��g_EDIT ���/%7����*SYSTEM*up�V9.40107� cr7/23/2�021 A���Pw��PRGA�DJ_p  h �$X[�p +$Y�xZ�xW�x���tZқtSPEED�_�p�p$NEXT_CYCLE�pg���q�FG�p� ��pALG�O_V �pNY�Q_FREQ�W�IN_TYP�q�)�SIZ1�O�LCAP�r!�[��M+�����qCREATE9D�r�IFY�r@!�NAM�p%h�_}GJ�STATU�оJ�DEBUG�rM_AILTI�����EVEU��LAS�T�����tELEM�� � $E�NAB�rN�EASyI򁼁AXIS�p$P߄�����q?ROT_RA" �rGMAX ��qE��-LC�AB
���C �D_LVՁ`�BAAS��`�1�{���_� κ�$x���RMr� RB�;�DIS����X_SPo�΁��� �u�P� |� 	� 2 m\�AN�� ��;�����Ӓ�� ��0�PAYLOx��3�V�_DOU�q�S���p�tPREF�� ( $GWRID�E
���iR���Y�  �p�OTOƀ�q  �p��!�p��k��OXY� � w$L��_POp|�נVa�SRV���)���DIREC�T_1� �2(�3�(�4(�5(�6(�7R(�8��qF��A�}� $VALu>�GROUP������F�� !"��@!��������RAN泲���Rx��/���TOTAX��F��PW�I=!>%�REGEN#�8� ������/���ڶnaTzЉ���#�_S����8�(�V[�'���4����GRE��w���Hp��D�����V_H���DAY3�V��S_�Y�Œ;�SUMM�AR��2 $�CONFIG_S�Eȃ���ʅ_RU�N�m�C�С�$CM�PR��P�DEVh���_�I�ZP��*Ӥ���ENHAN�CE�	�
�8��1���INT��q!M)b�q�2K�����OVRo�PGu�IqX��;���OVCT������v�
 4 �����a˟��PSL�G"�� \ @�;��?�1���SƁϕc�U������Ò�4�U�q]�Tp� (`�-��r�J<�O� CK�IL_MJ���VN�+�頓TQn{�N5���C��ULȀD�V(�CF6�P_�຀@�MW�[V1V�V1d�2s�U2d�3s�3d�4s�4d��'�	�������p	�IN	VIB1qp1� 2!pq/�,3 3,4 4 ,�p?��;��A���`N�������PL��TORr3�	���[�SAV���d�MC_FOL�D 	$SLP�����M,�I��L� �pL�b���KEEP_HNA�DD	!Ke�UC7COMc�k��
�lOP��p�pl��lREM��k��΢���U���ekHPW� �KSBM��ŠCOLLAB|�Ӱn��n�+�IT�O���$NOL�FCsALX� �DON�rx���� ,���FL���$SY�Ny,M�C=��~��UP_DLY�q=s"DELA� ��ڗ�Y(�AD��$TABTP_R�#��QSKIPj%g ����OR� �E�� P_��� �) ���p7��%9��%9 A�$:N�$:[�$:h�$:�u�$:��$:9�q�R=A�� X������MB�NFLIC]��0"�U!�o���NO_H� �\�< _SWITCHk��RA_PARAM=G� ��p��U��WJ��:Cӣ�_NGRLT� OO��U�����X�<A��T_�Ja1F�rAPS�W�EIGH]�J4CH�aDOR��aD��COO��)�2�_FJװ����sA�AV��C�HO1B.�.�l�J2�0�q-$�EX��T$�'QIT��'Q�pG'Q-�G��RDC�m"� � ��<��
R�]��
H���RGE�A��4��U�FLG0`g��H��ER	��SPC6R�rUM_|'P��2TH2No���@Q 1 �@ED���� � D �وIi�2+_P�25cS�ᰁ�+�L10_CI�8�pe� �pk� ���UՖD��zaxT�p�Q(�;a��c ��޲+�i���e��`� P`DESI�GRb$�VL1:i1�Gf�c�g10�_D�S��D��w�POS;11�q l�pr0��x1C/#AT�B���U
WusIND ��}�mqCp�mq`B	�oHOME�r 	a
Bq2GrM_q�P���!@s3Gr���� ��$�`!@s4GrG�Y�k�}�����
6�5Grď֏���(����6GrA�S��e�w�����6�7Gr���П�������8Gr;�M�_�q������S �q    �@sM��P�!�K@��! T`M��&M�IO��m�I��2�OK _OPy��� ¼�Q6�POWEG" 7�x EQ�1�E � #s%Ȳ$wDSBo�GNA�b�� C�P2�BS2;32S�$ �iP��9xc�ICE<@%�cPE`2� @IT���P�OPB7 1�FLOW�TRa@2���U$�CUN��`�AU�XT��2Ѷ�ERF�AC3İUU�v�CH��% t<�_9�EЎA$FREEFROM�¦�A�PX q�UP1D"YbA�PT.�pE�EX0����!�FqA%b�/��RV�a�G� &  j��E�" 1�AL� � �+�jc'��D�  2& �S\P~cP(
  �$7PB�%�R�2� ��T�`sAXU���DSP�ր�@�W���:`$��RN�P�%�@����K��_�MIR�����MT��AP���P"�qD�QSYz������Q{PG7�BRKH����ƅ AXI�  ^��i���1 �՞��BSOC���N���DUMMY16ށ1$SV�DE���I�FSPD_OKVR79� D��&��OR��֠N"`��F_����@OV��S�F�RUN��"F�0�����UF"@G�T�Od�LCH�"�%R�ECOV��9@�@W��`&�ӂH��:`_�0��  @�RTI�NVE��8AOFSr��CK�KbFWD��������1B��TR2�a�B �FD� �h�1= B1pBL�  �6� A1L�V��Kb�����#��@+<�A�M:��0��j��_�M@ ~�@h���T$�X`x ��T$HBAK���F��A�����PPA�
��	�������DVC_DB�3@pA�A�"��X1`�X3�`��S�@�`�0��U8ꣳ�h�CABPP
R �S #��c�B�@��>�GUBCPU�"��S�P�`R��11)�ARŲ�!$HW_CGpl�11� F&A1�Ԡ@8p�$UN�ITr�l e AT�TRIr@y"��CY�C5B�CA��F�LTR_2_FI�������2bP��CwHK_��SCT��F_e'F_o,�"�*�FS�Jj"CHA��Q�'91Is�82RS�D����1���_�Tg�`� i�EM�NPMf�T&2 8p�&2- �6DIAG~pERAILACNTBMw�LO@�Q��M7��PS��� � ,��PRBSZ`�`�BC4&�	��F�UN5s��RIN��PZaߠ�07Dh�RAH@���`� `C�@��`C�Q�CBLCU	RuH�DA�K�!�H�H�DAp�aA�H�C�EL�D������C��jA�1�CTIBUu�8p�$CE_RIA��QJ�AF P��X>S�`DUT2�0C���};OI0DF�_LC�H���k�LM�LF�aHRDYO,���RG�@HZ0���ߠ�@�UMULSE�P�'3iB$J���J����FAN�_ALM�dbWR=NeHARD�����P��k@2aN�r�J�_}�AUJ R�+4�TO_SBR ��~b�Іje 6?A�c_MPINF��{!��d�A�cREG�NQV��ɣZ�D��NsFLW%6r$M�@ � ��f� �0 h'u�CM4NF�!�ON	 e!e#�(b*r3F��3 �	 ���q)v5�$�$Y�r���Zu�_��p*7$ �/�EGE��ӌ��qAR��i���2p�3�u�@<�AXE��wROB��RED�֓WR��c�_���S�Y`��q� ?�SI�WcRI���vE STհP�ӭ d���Eg!�"�t8��^a��B����r��9�3� OTO�a9���ARY��ǂ0�1����FIE��ӿ$LINK�QGkTH��T_�������30���X�YZ���!*�OFIF�����ˀ	B��,Bl������m�FI� ��C@Iû�,B��_J$�F�����S`����3-!A$1�w0���R��C��&,�DU���3�P�3TUR`XS.�Ձb�bXX�� ݗFL��d���pL�0���34����� 1)�K��M�5�5%B'��ORQ�6��fC㘴��0B�O;�D�,�������a�OVE��rM�����s2��s 2��r1���0���0�g /�AN=!�2�DQ�q ���q�}R�*��6�`���s��V���ER��
jA	�2E��.�C��	A���0��XE�2Ӈ�A��AAX��F��A �N!�SŴ1_��Q_� ��^ʬ�^ʴ�^��0^���^ʷ�^�1&�^ƒP [ɒPkɒP{ɒP�ɒP �ɒP�ɒP�ɒP�ɒP������ɪ �R>�DEBU=#$8ADc�2����
�AB�7���r�V� <" 
�� i�q��-!��%��׆� �׬��״����1�י���׷�JT��DR�m�L�AB��ݥ9 FG�RO� ݒ=l� B_�1�u���}��`�����ޥ��qa��AND �����qa� �Eq��1��A@�� ��NT$`��c�VEL�1��m��1u���QP���m�NA[w�(�C�N1� ��3줙�  ?�SERVEc�p�+ $@@d@��M!��PO
�� _�0T !�򗱬p,  $TRQ�b
(� -DR2,+"P�0?_ . l"@!N�&ERR��"I� 8q���~TOQ����AL�p]�e���0G���%�����RE>�@ / ,��/�I -��RA� O2. d�&���_! 0�p$`&��2tPM��OC�A�8 1  pC�OUNT�� ��F�ZN_CFG2# 4B �f�"T�:# ��Ӝ� � `^�s3 ���M:0��R�qC@��/�:0�F!A1P��?V�X�� ���r���� �9P:b��HELpe�4 5��B�_BAS�cRSR�f @�S�!QY �1�Y 2|*3|*4�|*5|*6|*7|*8�L!RO�����3NL�q �AB���0nZ ACK��INT_uUS`�Pta9�_PU�>b%ROU��PH@�h9#�u`w��9�TPFWD_KcAR��ar RE���PP��A]@QUE��i&��	�f�>`QaI `��9#�j3r��f��SEME��6��PAn�STY4SO�0�DI'1�`���18��rQ_TM�cMANsRQXF�END��$KEYSWI�TCHj31:A�4H}E	�BEATM�3PE�pLE��1��J�HU~3F�42S?D�DO_HOMBPOl:a0EF��PRr�P�*�v�uC�@O�Q<o �OV_Mϒ��Eq�OCM���7���p8%HK�q5 �D��g�Uj�2M��p�4R��FORC��cWAR��NYOM>�p 6 @�Ԣ�*v`U|�P�p1�V'p��T3�V4��OR#Oʏ0L�R7��hUN�LOE0hdED>Va  �S�@dG8 <pAQ9�l1�MSUPG�UaC�ALC_PLAN�cc1��AYS1�1|:b�9 � X`��P �q;a�թ�w��2��j�M$P�㣒��fyt$��rSC�M �pm�q ���aq��0�jtYzZzEU�Q�b�� T!�Hr�pPv~	NPX_ASfw: 0g ADD���$SIZ%a�$VA��MUL�TIP�"ns�PA��Q; � $ T9op�B���rS��j!yC~ �vFRIF�2�S�0�YT�pNF[DODBUX�B��u&�!���CMtA�Е���������+Z >��< � �p��TEg�����$SG%L��T��X�&{��x�㰀��STMTe��ЃPSEG�2��ByW���SHOW؅n�1BAN�`TPO�@��gᣥ��������mV�_G�= ���$PC���O�F�B�QP\�SP�0A�&0^�� VDG���>� �cA00�����P���P���P����P��5��6��7*��8��9��A��b`����P��w᧖��F����h���1��v�h��י1�1�1��1��1�1%�12�1�?�1L�1Y�1f�2���2��2��2ʙ2�י2�2�2��2��2�2%�22�2�?�2L�2Y�2f�3���3��3��3ʙ3
י3�3�����U3�3%�32�3߹U3L�3Y�3f�4��U4��4��4ʙ4יU4�4�4��4�U4�4%�42�4߹U4L�4Y�4f�5��U5��5��5ʙ5יU5�5�5��5�U5�5%�52�5߹U5L�5Y�5f�6��U6��6��6ʙ6יU6��6�6��6�U6(�6%�62�6߹U6L�6Y�6f�7��U7��7��7ʙ7יU7��7�7��7�U7(�7%�72�7߹�7L�7Y�7f�[V��`_UPD��? y�c 
ZB�����@ x $gTOR�1T�  �caOP �, ZQ_7�RE^��� J��S�sC�A��_Ux�p��YSLOA"A � �u$�v���w�@���@��bVALUv10�6�=F�ID_L[C:�HI5I�R$FI�LE_X3eu4$��C7 �SAV��B� hM �E_BL�CK�3�ȁ�D_CPU��p��p5�hz��@S2R C � PW���� 	�!LAށS�R�#.!'$RUN�`G@%$D!'$�@G%e!$e!'%HR03$� �'$7aT2Pa_LI��RD  � G�_O�2�0P_EsDI�R�"SPD�#E�"i0ȁ�p�Q��DCS9@G)�F � 
$JPQC71��� S:C;}C9$MDL73$5P>9TC�`@7�UF�@?8S� ?8COBu �@�"|�L�G�P;;� 9�:;�qTABU�I_�!L�HGb�% �FB3G$��3A�sR�LLB_AVAI�B���3�!I $� SEL� NẼ�@RG_rD N��Ta���4{SC�PJ �1�/AB�PT�R?�w@_9M]`L�K \M f&/QL_��FMj��P�Gi�U9R�6��P+S_�P\� �p�E}E7B�TBC2�e�L ���``�`b$�!FT�P'T�`TDCg�� BPLp��sNU;WTH��qhhTgtWR�2$�pERVE.S�T;S�T�w�R_ACkP ?MX -$�Q�`@.S�T;S�PU@�`ICn�`LOW�GF1�QR2g�`��p�S�ERTIA�d^0i�P�PEkDEUe�LoACEMzCC#c�V�BrpTf�edg�a�TCV�l�adgTRQ�l�e�j|�Scu��e�dcu�J7_ 4JH!��Se@qde�Q�2�0���1�PRcuPJKlvVK<�~qcQ~q�w�spJ0��q�sJJv�sJJ�sAAL�s@�p�s�p�v���r5sS�`N1�l�p�k�`5d�XA_́� PCF�BN `M GRO�U ��bh�NPC�0sD�REQUIR�R� EBU�C�Q�6=g0 2Mz��P�d�QSGUO�@^�)APPR0C7@֍ 
$� N��CL	O� ǉS^U܉Se>@�BC�@A�"P �$PM]P�`�`sR�_MGa!�C���+���0�@,�BRK*�N�OLD*�SHOR�TMO�!m�Z��JWA�SP�tp`�sp`�s�p`�sp`�sp`�A��7:��8sQIR_�RTQ� m��R.Q��cQ�PATH �*� �*��X&���-P�NT|@A�"p�l�� �IN�RUC4`�a��C�`UM��Y
`�)p��>�Q���cP���p��PAYL�OAh�J2L& R_Am@�L ������+�R_F2LgSHR�T/�LO����0���>���ACR@L0z�p�y�ޤsRH�5b$H+���FL�EX��#�JVR P��_._�_�_�QJ�US : �_�Vd`0�G��_tQd`�_�_lF1G��ũǀo0oBoTofoxo��E �o�o�o�o�o�o�o  ����wz3lt���� 3EWF�^zT!��X���ju��uu~� W؁���p�u�u�u`�u����UM��(�T �P5�G�Y��' AT��l�pE�L0�_B��s�J�Svz�JEW�CTR7B�`NA��d�HAN/D_VB�����TUO@`+�`T�SW8F�A�V� $$M��e  G�AV�Qs�De�o�AA��@�	$�A(5�G�AU�Ad�� �6��G�DU�Dd�P2D�G/ -STI�54V�5Ng�DYF �� +�x����P&�G�&��A��lw�o�Q�k�P ������ʕӕܕ��sDX�TW 7 �� ��3%�?!OASYMT�(�m��T�V*�o�A�t�_SH�~������$����Ưد�J񬢐�p#39"���_VI���`8�q0V_UN!IrS�4��.�Jmu�2 ��2A��4X��4�6a��pt�������&E_�h����RE��CH( ?X ̱����TOc�PP�VPsSvD�US�RU�P��@���z@�D�A}@_5��U��P�EyAa��RPR�OG_NA��$>�$LAST����CANs�ISz@XYZ_SPu�DW]�R@Ͱ,VSV@�E1QE9Nc��DCUR�H#�ޜ�HR_T��Y�tQ9S�d��O��T 
Z�tQ?�SZ ��I�!A�D ���Q���#�S���� ��3�vP [ � -ME�O��R4#B�!T�PPT0F@1�a-�1�̰� h�1a%iT0� $DUMMY1���$PS_��RF���!�$lfװFLA*�YP�bc$GLB_TI ��U�e`ձ��LIF�(!\����g`OqW�P��eVOL#q�b �a_2��[d2 �[`����b�P�cZ`�TC��$BAUYDv��cST��B�2�g`ARITY0sD�_WAItAIyC,J2�OU6�ZqyyTLANS�`�{S��SZc��BUF_��r�fиx�PyyCH�K_�@CES��V� JO`E�aA<�x�bUBYT��� ��r�.�.� ��aA���M�������Q]c Xʰ����ST�����SBR@M2�1_@��T$SV�_ER�b����CL��`��A1�O�BpPG�Lh0EW(!^ 4� $a$Uq$�q$W�9�At�@R����Ӄ�Uم_ "��Dw$GI��}$ف� ^��(!`� L�.��"}$Fz�"E6�NEAR�N�B$F}��TQ�L���J�@R� �amP$JOIN�Ta�)�&ՁMSE]T(!b  +�Ec�2�^�ST��H�_�(!_c�  ��U��?���LOCK_�FO@� �PBGLmV��GL'�TE�@sXM���EMP�����K��b�$U�؂a�2_���q��`<� �q�^��C�E/�?��� $KA�Rb�M�STPDRqA܀����VECX������IUq�av�H=E�TOOL����V��REǠIS3d��6��ACH̐�m b^QONe[d3����IdB�`@$R�AIL_BOXE:a���ROB�@D��?���HOWWA�R0Aa�i`-�ROLMtb��$�*���T��`ܱ���O_FU�!>��HTML58QS��� e�"Հ�(!dF����@�(!e󲈁�����І}p(!f t��m�^a��t��B�PO��AIPE�N���O�����q��AORDED0�m �z�XT`��A�) ��P�O�P �g D �`OB�����ǯ�Uc�`���� ��SYS��A�DR��pP`U@^  �h ,"��f$�A��E��EтV�WVA�Qi �c �@ق�UPR�B>�$EDI�Ad�_VSHWRU�z�ƀ�IS�Uq�pND��P7���G�HEAD��! @���!i�KE�UqO`CP)P��JM�P��L�U�TR�ACE�Tj����IL�S��C��N�E���TICKt!M4�_N��{HNr�k @���HWC��P�FF��`gSTYeB+�LO�a�9�' ��[�C�l3�
L�@�F%$A��D=��S�!$�1�p aȌe�q�ePv �FSQ�U��#LO�b_1TGERC`!oPS?�m 5���R�m@3���ܡ�O`	c #IZ�d�A�eha�q�tb}�hA}pP~r��_SDO�B�X�pSSQN�SAXI�q��v��bS�U�@TL���RgEQ_ܠ��ET���`�CY%�P��Z&��A,f\!\d9x�P� MBSR$$nl-�w �����c
�uV
Qh(�AA���dC`�A�@�	�Y��D���p�E"�	CC�C���/�/�/	4IS}C�` o h��cDSmడ[`SP�@&�AT� 
R��L��XbADDR�s�$Hp� IF�Ch�_'2CH���pO����- �TUk�Ir p�CUCp�V��I�Rq�4���c��
K�
��^ ��N�Pr \z�D����|,K� P�"CN���*CƮ��!�TXS/CREE��s�Pp@�INA˃<�4�D�������`t T ᫀ�b����O Y6��0�º�U4h�RR��������R1�T  �;UE��u �j �qrz`Ś��RSML����U����V�1tPS_��6\��1�9G\����C��2@4 2��0Ov�R��&F~�AMTN_FL*��`Q��W� ��BB�L_/�WB`�Pw �����BO ��BL�E"�Cg�R"�DRI�GHtRD��!C'KGRB`�ET���G>�AWIDTHs����RB��a�r�UI溰EYհRx d��ʰ�����`y�B�ACK��tb>U����PFO��QWLAB��?(�PI��$URm�~P�P�P�Hy1 y 8 $�PT_��,"�R�PRUp�s5�da��R�QO%!t�zV�ȇ��pU�@�SR ���L�UM�S�� ERV�J��SP��T{ � " GE�Rh� L�¯�LPAeE���)^g�lh�lh�*ki5ik6ik7ikp�P`�Z�x����$u1x��p�Q zQ�USRل| <�z��PU2�a#2�FO\O 2�PRI*m9��[�@pTRIPK��m�UNDO��})���Yp��y�����h����p ~��Rp�qG ��T0���-!�rOS2��vAR��2�s�CA⏐����ro���Pi�UIaCA����3Ibn�N�sOFFA�D@��%�Ob�r���L�,t��GU��Ps���p�����+QSUBo�� ��E_EXE���VeуsWO� ��#��w��WA�l�p΁fP
 V�_DB���pT��pO�V░���3O9R/�5�RAU@6��TK���__���� |j �OWN|j�34$SRC�0�`���DA���_MP�FI����ESP ��T�$0��c��g�pY�q�z�E!� `%��ۂ34J���COP&��$���p_���0/�+�6���CT�Cہ��ہ�D �DCuS��P4�gCOMp�@�;��Oo�=���XK�^�/�VT�q'���Y٤Z��2��0�@p�w#SB����(2�\0˰_��M��%!�]�DIC#��AY\�3G�PEE�@T�QFS�VR1���eQL�� a��P�D ��f� z��f�> ���6�FPq�A�t�b# �L2?SHADOW��#~ʱ_UNSCAd��׳OWD�˰DGD}E#LEGAC)�^q'�VC\ C��� v�������m�RF07���7d`yC2`7�DRIVo�	��ϠC�A]�(�` ����MY_UBY �d?Ĳ��s��1��$0�����_ఆ���mL��BM�A$�7DEY	�EXp@C�/�MU��X��,��0cUS��.�;p_R"1��0p#�2�GP�ACIN*���RG ��c�y�:�y��sy�C�/�RE�R"!�q��8�y�D@� L !��G�P�"�г��R�pD@�&P�Px1Q���	.���RE��SW&q�_Ar��+�{��Oq�AA/�3�hErZ�U���� PV�HK���PJ���_/�Q0{�EAN���ۀ2�2��P�MR�CVCA� �:`O#RG��Q�dR	��L�����REFoG���� ��!�+`	�p���@�����<���q�_����r��� S�`C���p��G�@D� ��0��!��#q�š�OUx����?� ����2�J@0� 1�*p�����0 UmL�@��CO�0f)��� NT� [��Z�Qf�af% L飏��Q��a��VIAچ� ̈́�@HD7 6P$�JO�`oB�$�Z_UPo��2Z_LOW��$�QiB<n��1$EP�s��y�� 1!f m�� 1¦4� 5��PA�A �C7ACH&�LO�w@�ВQB���Cn�%I#F^��Tm��N��$HO2�32{��Uÿ2O�@���R`o��=a��ƐVP��<X@A"_SIZ&�K$�Z$�F(�G'���CM]Pk*FAIo�G���AD�)/�MR1E���"P'GP�0����9�ASYNBUFǧRTD�%�$P!��COLE_2D_D4�5W�sw�~�U��QO��%ECCU��VEM��v]2�VIRC�!5�#�2��!_>�*&�pWp��AuG	9R�XYZ@�3�W���8��4+Q2z0T"��IM�16��2P�GRABB��q��;�LERD�C ;�F_D��F�fC50MH�PE�R�[���� ��KQLAqS�@��[_GEb� �H൑~23�E�T����"���b��I��D�ҙ6m�BG_L3EVnQ{�PK|Л6,\q��GI�@N\P4�An��A��!g�drҍS� �NRT�VLʁc�Ų��#ah��c"!D�qDE�@���Xа�X����(�1��d��pzZ����d�c���D4q�Բ�2pT��U&�� -$�ITPr9p[Q8��ՓV�VSF$�d��  fp/�f�U�R&ҿ�SMZu�dr��ADJ`C�� ;ZDVf� D�X�AL� � 4 PE�RIKB$MSG_Q3$Q!o%[���p'��dr:g�q�Q� �XVR\t�̆B�pT_\��R��/ZABC"����Sr䚣�
W��aACT�VS' � �� $|u�0�cCT3IV�Q!IOu¥s�&D�IT�x�DVFϐ
x�P���!����pPS���� ��#��!���q!LS�TD�!�  �_S�T���aq�CHx�� L-�@��u��Ɛ*���P GNA�#�C�!q�_FUiN�� uqIPu�3�HR�$L���}XZMPCF"���`bƀ�rX�ف��LNK��
Ł�0#�?� $ !��^ބCMCMk�C8��C"����P{q O$J8�2�D6! >�O�H���T���2������M���UX�1݅UXE1Ѡ��1C���Y����������˗7�FT�FG>�������Z���� �k�� ���YD'@ �� 8n�R� U�ӱ$HEIGH�d�:h?(! 'v�������� � Gd��qp$B% � E���SHIF��hR�Vn�F�`�HpC � 3�(�8H`O�ѡ�ȭC��+%D	�"�CE�pV���SPHE}Rs� � ,! �M�c�u��$PO?WERFL �R|�e���|�p�RG�`ް�������A�  ���?`��`d��NS�b ����?�  Bz�|� l�  <@�|��%����������ŵ�� 2�ӷ�� 	H��l�&���>��w�A |��t$���*��/�� **:��`�ϥ��͘���������ɘ��|�����5����� ��%ߟ�I�[߉�� ������������w� !�3�a�W�i����� ������O����9�/� A���e�w�������' �����=O }s������ �k'UK]� �����C/�� -/#/5/�/Y/k/�/�/ �/?�/�/?�/?�? 1?C?q?g?y?�?�?�? �?�?�?_O	OOIO?O<QO�� 	 �O�O �O_�E��3_���O`_��O�_�_÷PREF� Ӻ``
���IORITY �`|���`����pSaPL`z����WUT�V�qÈ�ODU~��e���_?�OG���Gx��R��,fHIB�qOy�|kTOEN�T 1��yP(!AF_b�`�o�g?!tcp�o}�!ud�o)~!icm�0b�XY̳�k �|�)� ����������u��� ���N�5�r�Y���@����̏�����*/c̳ӹ���E�W�|��>��A�F��/���4���|��,�7�A~��,  ��P�����%�|�'���Z��h�z�����|���ENHANCE 	#�7�s�7��d�����  �D,f�T
�_�S����OPORTe�rb����U��_CAR�TREP�Pr|brS�KSTAg�kSL�GS�`�k������Unothing�������Ϳ>�P�b�To��TEMP ?isϨE�/�_a_seibanm_��i_��� ��0��T�?�x�cߜ� �ߙ��߽������� >�)�N�t�_���� ����������:�%� ^�I���m��������� �� ��$H3l Wi������ �D/hS��w���uϪ�VE�RSI�P=g  �disabl�e��SAVE �?j	267_0H705���k/!�m//*�/ !	�(%b�O�+�/�S�e?6?H?Z?l?z:�%<�/�?4�*'_j` +1�kX �0ub�uE�?OqG�PURG�E��Bp`�ncqWF <@�a�TӒ*fW�`]D�aa�WRUP_DELAY z��f�B_HOT �%?e'b��OnER_?NORMAL�HGbx�O%_�GSEMI_�*_i_�QQSKIP�3.��3x��_� �_�_�_�]?eo+go Ko]ooo5o�o�o�o�o �o�o�o�o5GY i�}���� ���1�C�U��y� g���������я�����-�?�7%�$RA?CFG �[ќ��3�]�_PAR�AM�Q3y��S �@И@`�G�42�C۠��2��C�bFB�B]�BTI�F���J]�CVTMkOU�����]��DCR�3�Y ���Q@%x��B!huA��?�1�>�a�9����]�'����"�+��g�y�-�1���@�1ϱ�_��o� ;e�m����KZ;�=g;�?4�<<���f@8����� �5� G�Y�k�}�������ſ�׿���xURDIO_TYPE  �V��5��EDPRO�T_a�&,>��4BHbCEސS�v�Q2c� ��B�ꐪϸ���ϐ� ���&�ݹ�W�V_~� o����߱������� ��A�O�m�r���9� ������������� �=�_�d������� ����������'I� Nm����� ����#EJi +k����� �//4/F//g// �/y/�/�/�/�/�/	? +/0?O/?c?Q?�?u? �?�?�?�?�??;?,O���S�INT 2��I���l�G;� �jO|K��鯤O�f�0 �O�K�?�O�?_ __N_<_r_X_�_�_ �_�_�_�_�_�_&oo Jo8ono�ofo�o�o�o �o�o�o�o"F4 j|b����������B�O�EFPOS1 1"�?  xO�� o×O����ݏ鈃��� Ϗ0��T��x���� 7���ҟm�������� >�P����7������� W��{�����:�կ ^����������S�e� �� ��$Ͽ�H��l� �iϢ�=���a��υ� � ߻����h�Sߌ� '߰�K���o���
�� .���R���v��#�5� o����������<� ��9�r����1���U� ����������8#\ ����?��u ��"�FX� ?���_��/ �	/B/�f//�/%/ �/�/[/m/�/?�/,? �/P?�/t??q?�?E? �?i?�?�?O(O�?�? OpO[O�O/O�OSO�O wO�O_�O6_�OZ_�O ~_�_+_=_w_�_�_�_ �_ o�_Do�_Aozocf�2 1r�o.o ho�o�o
o.�oR �oO�#�G�k �����N�9�r� ���1���U������� ���8�ӏ\���	�� U�����ڟu�����"� ���X��|����;� į_�q������	�B� ݯf����%�����[� ��ϣ�,�ǿٿ� %φ�qϪ�E���i��� ����(���L���p�� ��/�A�Sߍ������ ��6���Z���W��+� ��O���s������ ��V�A�z����9��� ]���������@�� d��#]��� }�*�'`� ��C�gy� �&//J/�n/	/�/ -/�/�/c/�/�/?�/ 4?�/�/�/-?�?y?�? M?�?q?�?�?�?0O�?�TO�?xOO�O�o�d3 1�oIO[O�O_ �O7_=O[_�O__|_ �_P_�_t_�_�_!o�_ �_�_o{ofo�o:o�o ^o�o�o�o�oA�o e �$6H�� ���+��O��L� �� ���D�͏h�񏌏 �����K�6�o�
��� .���R���퟈���� 5�ПY�����R��� ��ׯr��������� U��y����8���\� n�������?�ڿc� ����"τϽ�X���|� ߠ�)�������"߃� nߧ�B���f��ߊ��� %���I���m���,� >�P���������3� ��W���T���(���L� ��p�����������S >w�6�Z� ���=�a�  Z���z/ �'/�$/]/��//�/@/�/�O�D4 1�Ov/�/�/@?+?d? j/�?#?�?G?�?�?}? O�?*O�?NO�?�?O GO�O�O�OgO�O�O_ �O_J_�On_	_�_-_ �_Q_c_u_�_o�_4o �_Xo�_|ooyo�oMo �oqo�o�o�o�o�o xc�7�[� ���>��b�� ��!�3�E����ˏ� ��(�ÏL��I���� ��A�ʟe������ �H�3�l����+��� O���ꯅ����2�ͯ V����O�����Կ o�����Ϸ��R�� v�Ϛ�5Ͼ�Y�k�}� ����<���`��τ� ߁ߺ�U���y��� &���������k�� ?���c������"��� F���j����)�;�M� ��������0��T ��Q�%�I�mx��/�$5 1�/ ���mX��� P�t�/�3/� W/�{//(/:/t/�/ �/�/�/?�/A?�/>? w??�?6?�?Z?�?~? �?�?�?=O(OaO�?�O  O�ODO�O�OzO_�O '_�OK_�O�O
_D_�_ �_�_d_�_�_o�_o Go�_koo�o*o�oNo `oro�o�o1�oU �oyv�J�n �������u� `���4���X��|�ޏ ���;�֏_������ 0�B�|�ݟȟ���%� ��I��F�����>� ǯb�믆������E� 0�i����(���L��� 翂�Ϧ�/�ʿS��  ��LϭϘ���l��� ��ߴ��O���s�� ��2߻�V�h�zߴ��  �9���]��߁��~� ��R���v����#�	6 1&���� �����������}� ��<��`��� �CUg��& �J�n	k�? �c��/��� 	/j/U/�/)/�/M/�/ q/�/?�/0?�/T?�/ x??%?7?q?�?�?�? �?O�?>O�?;OtOO �O3O�OWO�O{O�O�O �O:_%_^_�O�__�_ A_�_�_w_ o�_$o�_ Ho�_�_oAo�o�o�o ao�o�o�oD�o h�'�K]o �
��.��R��v� �s���G�Џk�􏏏 ���ŏ׏�r�]��� 1���U�ޟy�۟��� 8�ӟ\������-�?� y�گů����"���F� �C�|����;�Ŀ_� 迃������B�-�f� ϊ�%Ϯ�Iϫ���πߣ�,���P�6�H�7 1S����I��� ��������3���0� i���(��L���p� �����/��S���w� ���6�����l����� ��=������6� ��V�z�  9�]���@ Rd���#/�G/ �k//h/�/</�/`/ �/�/?�/�/�/?g? R?�?&?�?J?�?n?�? 	O�?-O�?QO�?uOO "O4OnO�O�O�O�O_ �O;_�O8_q__�_0_ �_T_�_x_�_�_�_7o "o[o�_oo�o>o�o �oto�o�o!�oE�o �o>���^� ����A��e� � ��$���H�Z�l���� �+�ƏO��s��p� ��D�͟h�񟌟��� ԟ�o�Z���.��� R�ۯv�د���5�Я�Y���}�c�u�8 1��*�<�v���߿� �<�׿`���]ϖ�1� ��U���y�ߝϯ��� ��\�G߀�ߤ�?��� c����ߙ�"��F��� j���)�c������ �����0���-�f�� ��%���I���m���� ��,P��t� 3��i��� :���3�� S�w /��6/� Z/�~//�/=/O/a/ �/�/�/ ?�/D?�/h? ?e?�?9?�?]?�?�? 
O�?�?�?OdOOO�O #O�OGO�OkO�O_�O *_�ON_�Or___1_ k_�_�_�_�_o�_8o �_5ono	o�o-o�oQo �ouo�o�o�o4X �o|�;��q ����B���� ;�������[���� ���>�ُb�����!��������MASK +1 �������~ΗXNO  ݟ����MOTE  ����S�_CFG !Z���N�����PL_RANGV��N������OWER� "��Ϡ��S�M_DRYPRG7 %���%W���եTART #�Ǯ�UME_PR�O���q���_EX�EC_ENB  y����GSPDJ�쌰����TDB̯���RMп��IA_OPTION��֋����NGoVERS���`�řI_AIR7PUR�� R�+�\��ÛMT_֐T �X���ΐOBOT�_ISOLC����������NAM�E8��H�ĚOB_CATEG�ϣ,���S�[�.�ORD_NUM ?Ǩ���H705  N��ߨߺ��ΐPC_TIME�OUT�� xΐS7232s�1$���� LTEA�CH PENDAaN��o���)���V�T�Main�tenance /ConsN�&�M��"B�P�No Use6�r�8����p����̒��NPO$���Ҏ�"���CH�_LM�Q���	�a�,�!UD1:��.�RՐVAIL�w��粥*�SRW  t� ����5�R_INTVAL���� ����V_DATA_G�RP 2'����/ D��P��� ����	����� �B0RTf ������/� />/,/b/P/�/t/�/ �/�/�/�/?�/(?? L?:?p?^?�?�?�?�? �?�?�?O O"O$O6O lOZO�O~O�O�O�O�O �O_�O2_ _V_D_z_ h_�_�_�_�_�_�_�_ o
o@o.oPovodo�o���$SAF_D?O_PULSW�[�xS���i�SCAN�Ҳ�����SCà(�3�4о��S�S�
������q�q�qN� �L^p� ��5��� ���$��+��r2M�qqdY�P�`�J�9	t/� @���� ����ʋ|��� r ք��_ @N��T ��'�9�K�X�T D��X����� ����ɟ۟����#� 5�G�Y�k�}�������<䅎������Ǧ  "�;�#oR� ���p"��
�u��Di���q$q�  � ���uq%�\��� ����ҿ�����,� >�P�b�tφϘϪϼ� ��������(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z����珈�������� ����g�;�D�V�h� z���������������(�Ӣ0�r�i�y��� $�7I[m�� �����!3 EWi{���� ���////A/S/ e/w/�/�/�/�/�/�/ �/?r�+?=?O?a?s? �?�?�?�?�?8��?O O'O9OKO]OoO�O�� $�r�O�O�O�O	_ _-_?_Q_c_u_�_�Y �_�_�_�_�_oo&o 8oJo\ono�o�o�o�o �o�o�o�o"4F Xj|�c�路g� ������0�B� T�f�x���������ҏ������:�Ҧ���y�3�	�	�1234567�8��h!B�!�� \��p0����Ο��� ��(�:�@��c�u� ��������ϯ��� �)�;�M�_�q����� R���ɿۿ����#� 5�G�Y�k�}Ϗϡϳ� ���ϖ�����1�C� U�g�yߋߝ߯����� ����	��-���Q�c� u����������� ��)�;�M�_�q��� B���������� %7I[m�� ������!3 EWi{���� ���////�S/ e/w/�/�/�/�/�/�/ �/??+?=?O?a?s? �?D/�?�?�?�?�?O O'O9OKO]OoO�O�O �O�O�O�O*����O�	_�E�?5_G_Y_�y�Cz  A��z �  ��x2�r� }��)�
�W�  	�*�2�O�_�_ oo"l�#\��_hozo �o�o�o�o�o�o�o
 .@Rdv�� ��Mo����*� <�N�`�r��������� ̏ޏ����&�8�J�B�X #P$P�Q�R<u�� k��Q  ������S�P��|�Q�Qt  �PhÙ۟�P(� `,b�����]�PFl�$�SCR_GRP �1*4+4�4 � �,a� �U	 �v�� ~������d���%���pɯ���h]��P~�D1� D7n�3��Fl
CR�X-10iA/L� 2345678+90�Pd� r��P�d�L ��,a
�1o��������[ ¶~�+fm�ͣm��Fcg�p�����ӹ	�Ĳ�.�@�R�d�t���H�~�Ă�m��ϴ������ϼ��,a��1���U�[��G�imXhuP,[~��u��B�  B!ƠߞҷԚ�A�P���  @1`�՚�@������ ?���H����ښ�F@ F�`A�I�@�m�X� ��|���������� �������:�%�7�I�[�B�i�������� ��������-Q< u`��En�ٯ����W�P�"+f@@_�5��1`b���x����ͣ�O�,dAA�������Fa�,a �#!"/4/E-!Z(f/x/NG/ (�P�!(�  �/�/�/��/�/?#9Ab����S7س�M��ECLVL  �,a��ݲ�Q@�f1L_DEFAU�LTn4b1��1`�3HOTS�TR�=��2MIP_OWERFm0pUz�5�4WFDO�6� �5L�ERVENT 1+u1u1�3� L!DUM�_EIP#?5H�j�!AF_INEx�0SO,d!FT)O��NIO�O!���O ���O�O!RP?C_MAIN�O�Hq��O>_SVIS_��I�-_�_!OPcCUf�_�Wy_��_!TP�PPU��_<Id�_"o!
P�MON_PROX	Y#o?Feono�R<o�8Mf]o�o!RD�M_SRV�o<Ig�o!R��"=HYh�oR!
PM�o�9LiA�!RL�SYNC��y8|��!ROS(O���4�6�!
C}E�PMTCOM7��?Fk%���!	K�C'ONS��>Glq�Ώ�!K�WASRCd�o?Fm���!K�'USB�=Hn	�f�!STM�0��;JoU����O֟�c�����CICE_KL �?%K (%SVCPRG1��DG�1�2G�L�6�3o�Dt�6�4����6�5��Dį6�6��6�7� �6���W�R�9_�d�3���6�9���6� a�ܿ6����6���,� 6�ٯT�6��|�6�)� ��6�Q���6�y���^� ���^�ʿD�^��l� ^�ϔ�^�Bϼ�^�j� ��^����^���4�^� ��\�^�
߄2�� �6��/����V�� <�'�`�K���o����� ��������&J 5nY����� ���4F1j U�y����� /�0//T/?/x/c/ �/�/�/�/�/�/�/? ?>?)?P?t?_?�?
�_DEV I��MC:�84����4GRP �2/E�0+�bx� 	� 
 ,
@�0�?OD8O JO1OnOUO�O�O�O�O �O�O�O�O"_	_F_-_ j_|_c_�_�[O�_�_ �_o�_,ooPo7oIo �omo�o�o�o�o�o��o(:!^�_  �1i@���� ��� �=�$�a�s� Z���~��������؏ �l
�K���qp�W� �Q���	�Ο���� �(��L�3�E���i� ����ʯܯ�_ ��ɯ 6��Z�A�~���w��� ��ؿ�ѿ���2�D� +�h�Oό�s�9���]� ���ϳ��ߙ�'�� v�]ߚ߁߾��߷��� ���*��N��r�� ;������������ &�8��\�C���g�y� ����������g�4 -jQ�u�� ���B) fx_����) ��/,//P/7/t/ [/m/�/�/�/�/�/? �/(??L?^?E?�?�7�d �[~
�6� s 	 A�;*=� 6?��=���D�>����g�:��0��ī���|@�-�@�5�_�eA5��-�=BG+h�&����6)AB��m����`�x��=�?7O%T�ELEOP8OcN�[~y��5�o��ʾTF������������|��ҝ�����E�1�E@��*�A`�~��n�!��$�A����M�Y<T��������C=�J����Gc��McO��I�JO/_�[~���6r _�1<��׻��y;���	A`�ʛ1bP���N	V�A�&�@в@����@)E�]�1������0ד� �x���Q��?U?�Q��O�_ _ _oDS�I�I2o o�VoDozoho�o�o%� o�o�_�o�o0 TBx�o��oh� d���,��P�� w��@�����Ώ��ޏ ��(�j�O������ p�����ʟ��ڟ �B� '�f��Z�H�~�l��� ��Ư������د��  �V�D�z�h����ſ �������
��R� @�vϸ���ܿf��Ͼ� �������Nߐ�u� ��>ߨߖ��ߺ�����  �V�|�M��&��n� ��������.��R� ��F���V�|�j����� �����*���B 0Rxf���� ���>,N t���d��� �//:/|a/s/*/ L/&/�/�/�/�/�/? T/9?x/?l?Z?|?~? �?�?�?�?,?OP?�? DO2OhOVOxOzO�O�O O�O(O�O_
_@_._ d_R_t_�O�O�_ _�_ �_�_oo<o*o`o�_ �o�_Po�oLo�o�o�o 8zo_�o(� �������R 7�v �j�X���|��� ���*��N�؏B� 0�f�T���x�����՟ 矞������>�,�b� P���ȟ���v��ί ���:�(�^����� įN�����ܿʿ��  �6�x�]Ϝ�&ϐ�~� �Ϣ�������>�d�5� t��h�Vߌ�z߰ߞ� �����:���.���>� d�R��v������� �����*��:�`�N� �������t����� ��&6\����� L������" dI[4|� ����<!/`� T/B/d/f/x/�/�/�/ /�/8/�/,??P?>? `?b?t?�?�/�??�? O�?(OOLO:O\O�? �?�O�?�O�O�O _�O $__H_�Oo_�O8_�_ 4_�_�_�_�_�_ ob_ Go�_ozoho�o�o�o �o�o�o:o^o�oR @vd���� �6�*��N�<�r� `������Ϗ������ ��&��J�8�n����� ԏ^�ȟ��؟ڟ�"� �F���m���6����� į��ԯ֯��`�E� ���x�f��������� п&�L��\���P�>� t�bϘφϼ�����"� ��ߨ�&�L�:�p�^� ���ϻ��τ������  �"�H�6�l�ߓ��� \������������ D���k���4������� ������
L�1C�� ��d����� $	H�<*LN `����� � //8/&/H/J/\/�/ ��/��/�/�/?�/ 4?"?D?�/�/�?�/j? �?�?�?�?O�?0Or? WO�? O�OO�O�O�O �O�O_JO/_nO�Ob_ P_�_t_�_�_�_�_"_ oF_�_:o(o^oLo�o po�o�o�_�oo�o  6$ZH~�o� �n�j���2�  �V��}��F����� ��ԏ
���.�p�U� �����v��������� П�H�-�l���`�N� ��r��������4�� D�ޯ8�&�\�J���n� ���˿
�������� 4�"�X�F�|Ͼ���� l���������
�0�� Tߖ�{ߺ�D߮ߜ��� �������,�n�S�� ��t�������� 4��+������L��� p����������0��� $46H~l� ������  02Dz���j ����/
/,/� �y/�R/�/�/�/�/ �/�/?Z/??~/?r? ?�?�?�?�?�?�?2? OV?�?JO8OnO\O~O �O�O�O
O�O.O�O"_ _F_4_j_X_z_�_�O �__�_�_�_ooBo 0ofo�_�o�oVoxoRo �o�o�o>�oe �o.������ ��X=�|�p�^� �����������0�� T�ޏH�6�l�Z���~� ������,�Ɵ �� D�2�h�V���Ο��� |��x����
�@�.� d�����ʯT������ п���<�~�cϢ� ,ϖτϺϨ������� �V�;�z��n�\ߒ� �߶ߤ�������� ����4�j�X��|�� ����������� 0�f�T��������z� ������,b �����R���� �j�a�: ������ /B '/f�Z/�j/�/~/ �/�/�//�/>/�/2?  ?V?D?f?�?z?�?�/ �??�?
O�?.OORO @ObO�O�?�O�?xO�O �O_�O*__N_�Ou_ �_>_`_:_�_�_�_o��_&oh_Mo�_�P��$SERV_MA_IL  �U�`���QvdOUTPU}T�h�P}@vdRV 20f;  �` (a\o<�ovdSAVE�l�i�TOP10 21��i d 6� s�P6r _ �a2oXj|��� ������0�B� T�f�x���������ҏ �����,�>�P�b� t���������Ο������(�:�guYP��cFZN_CF�G 2e��c�T�a�e|�GRP� 23��q ,�B   AƠ�QD�;� BǠ� � B4�SRB{21�fHELL�C4ev�`�o��|/�>�%RSR>� ?�Q���u�����ҿ�� ����,��P�;�t�h_Ϙϩ����s`��¼����Ϸͻ�b�P�&�'�ސW
��2�Pd��g���HK 15�� ,ߡ߫ߥ������� ��@�;�M�_�������������OMM 6��?���FTOV_ENB��d�au�OW_R�EG_UI_��bIMIOFWDL*��7.�ɥ��WAIT�\�`ٞ����`����d��TIM�������VA�`����_�UNIT[�*yL]Cy�TRY��u-v`ME�8���a�w֑d ��9� ������<���X�Pڠ6p`?�  ��o+=�`VL��l�fMON_AL�IAS ?e.��`heGo���� ��/)/;/M/�q/ �/�/�/�/d/�/�/? ?%?�/I?[?m??�? <?�?�?�?�?�?�?!O 3OEOWOO{O�O�O�O �OnO�O�O__/_�O S_e_w_�_�_F_�_�_ �_�_�_o+o=oOoao o�o�o�o�o�oxo�o '9�o]o� �>������ #�5�G�Y�k������ ��ŏ׏������1� C��g�y�����H��� ӟ���	���-�?�Q� c�u� �������ϯ� ����)�;��L�q� ������R�˿ݿ�� Ͼ�7�I�[�m��*� �ϵ������ϖ��!� 3�E���i�{ߍߟ߱� \�����������A� S�e�w��4����� ������+�=�O��� s���������f����� '��K]o� �>����� #5GY}�����l�$SMO�N_DEFPRO�G &����� &�*SYSTEM*����RECAL�L ?}� (� �}
xyzr�ate 11 >�192.168.�56.1:227�12 *=V/2 `f!�/�/�/�,}K' k/g/y/
??.?�&J/ �/X? ?�?�?�?�/Z? �?~?O!O3OF?�?�?��?�O�O�O�?lK15124iO{O__0_��Dtpdisc 0�O�@�O�O�_�_��_�Etpconn 0ULb_t_oo�)o�K8copy �frs:orde�rfil.dat� virt:\tmpback\S_��@�o�o�o�M/Kbm?db:*.*`oro`{o0�D3xKd:\�oUp�o�@�o�(���@4KuaSe �E��#�5�HK�� ��������E�O]D880�`j�|���1��CK_߇����� �����_ULb�t��� )�<�NE֟�������8���O�O716�^z�`��/�B_֯6 � ��������T�f�x� 	��-�@�R������ �ϩϼ�ί�r��� '�:oLo^o��67ߔ� �߹o�of���{��� 0�C��h����ߐ�� ���X�j������#� 5�H������������<Ə�Y4772h�z� /B��� ���� �����ULbt)��7K�]�So���}.��f�� z////B�2K�^� ����/�/�/F���d/ ��/?"?4?GY� ��?�?�?�`?�{? OO0OC/�?�/y/�O �O�O�/�/dO�/__ ,_??Q?�?u?�_�_�_ �?�?j_�?oo(o7k��$SNPX_A�SG 2:����Va� 7 0D�%�7o~o�  ?�GfPAR�AM ;Ve^`a �	lkP>��D�>��d�� ��I`OFT_�KB_CFG  �C�\eFcOPIN_SIM  Vk�b+=OYsI`�RVNORDY_�DO  �eu�krQSTP_DS�B~�b�>kSR� <Vi � =&c`ELEO�e��>�>�W`I`TOP_ON_ERRx�Gb�PTN zVeP��D:��RING_PRM�'��rVCNT_GOP 2=Ve�ac`x 	���DИ�яؼ���BgVD�RP' 1>�i�`�Vq ؏0�B�T�f�x����� ����ҟ�����,� >�e�b�t��������� ί���+�(�:�L� ^�p���������ʿ� � ��$�6�H�Z�l� ~ϐϷϴ��������� � �2�D�V�}�zߌ� �߰���������
�� C�@�R�d�v���� ������	���*�<� N�`�r����������� ����&8J\ n������� �"4[Xj| �������!/ /0/B/T/f/x/�/�/ �/�/�/�/�/??,? >?P?b?t?�?�?�?�?��?�?�?O�PRG�_COUNT�f9�P�)IENBe�+E�MUC�dbO_UPD� 1?�{T  
ODR�O�O�O�O�O __A_<_N_`_�_�_ �_�_�_�_�_�_oo &o8oao\ono�o�o�o �o�o�o�o�o94 FX�|���� �����0�Y�T� f�x����������� ���1�,�>�P�y�t� ��������Ο��	�� �(�Q�L�^�p����� �����ܯ� �)�$� 6�H�q�l�~������� ƿؿ���� �I�D��V�"L_INFO {1@�E�@��	 yϽϨ�����ɽվU>?>��=>�����A����Aԫ���g2�@C�0���B�J��ϟ  >@O�i�=���� D��@BQs�A���*C2�/?�?�kB��p߂��-@YSDEBUG�:@�@�o�d�I��S�P_PASS:E�B?��LOG uA���A  o�9i�v�  �Ao�UD1:\��<}���_MPC�ݚEHk�}�A&�� �A~K�SAV B��`IA���*�i�1��SVB�TEM_T�IME 1C����@ 0��n�ŧi�d��*���ME?MBK  �EA��������X�|�@� V�������������h�,9
�� ��@�` r�������� �@R dv�����
Le�//(/:/L/^/ p/�/�/�/�/�/�/�/� ??$?6?H?Z?��SKV�[�EAj��?�?�?V��+�@]2��|�?i�  0`o� ^
:O.@R�O�O�O}N�o�� ��OB�P�O_'_9_-L2�Y_�_�_�_�_�_o�$�_�_� o'o9oKo]ooo�o�o �o�o�o�o�o�o#�5GYk_?T1SVGUNSPD��� '����p2M�ODE_LIM #D��Ҋt2�p�q�E�݉uABUI_DCS H}5B���0�G�n��D���|-�X�>���*���� 
��e����E��r�i������uEDIT I���xSCRN �J���rS�G �K�.�(�0߅SK_OPTION�и^����_DI��ENB  -�����BC2_GRP 2L���MP�C�ʓ�|BCCF2/�N���� =����C8���\�G� ��k�������گů�� �"��F�1�C�|�g� ����Ŀ���ӿ�� 	�B�-�f�QϊϜ�ʂ �϶�������v��
� /�U�@�yߧ��`�i� ���߰�����
���.� �>�@�R��v��� ��������*��N� <�r�`����������� ����̀4FX ��|j����� ��B0fT vx�����/ �,//</b/P/�/t/ �/�/�/�/�/�/�/(? ?L?d?v?�?�?�? 6?�?�?�?O O6OHO ZO(O~OlO�O�O�O�O �O�O�O __D_2_h_ V_�_z_�_�_�_�_�_ 
o�_.oo>o@oRo�o vo�ob?�o�o�o �o<*Lr`�� ������&�� 6�8�J���n�����ȏ ���ڏ��"��F�4� j�X���|�������� ֟��o$�6�T�f�x� ��������ү����� ��>�,�b�P���t� �������ο��(� �L�:�\ς�pϦϔ� �ϸ������� ��H� 6�l�"��ߖߴ����� V������2� �V�h� z�H���������� ����
�@�.�d�R��� v������������� *N<^`r� ������&8 �\Jl���� ����"//F/4/ V/X/j/�/�/�/�/�/ �/?�/?B?0?f?T? �?x?�?�?�?�?�?O �?,O�DOVOtO�O�O O�O�O�O�O�O_ V�4P�$TBCSG_GRP 2O U��  ��4Q 
 ?�  __q_[_�__�_ �_�_�_�_o%k8R?S�QF\d�H�Ta?4Q	 HA����#e>���>�$a�\#eAT��A WR�o�hdjma��G�?Lfg�bpܚo�n�ffhf�̑ͼb4P|j��o*}@���Rhf�ff>G�33pa#e<qB�o�+=xrRp�qUy�rt~��H�y rIpTv�pBȺt~	xf 	x(�;���f���N��`���ˏڋ����	�V3.00WR	�crxlڃ	�*��3R~t��H�H��� \�.�]�  cC.�����V8QJ2?SRF]��~��CFG T U�PQ SPܚ���r�ܟ1��1�W�e�	Pe���v� ����ӯ������� �Q�<�u�`������� ��Ϳ�޿��;�&� _�Jσ�nπϹϤ��� ����WRq@�0�B� ��u�`߅߫ߖ��ߺ� �����)�;�M��q� \������4Q _�� �O ���J�8�n�\� �������������� ��4"XFhj| ������ .TBxf��nO ����//>/,/ b/P/�/t/�/�/�/�/ �/�/�/?:?(?^?p? �?�?N?�?�?�?�?�? �? O6O$OZOHO~OlO �O�O�O�O�O�O�O _ _D_2_T_V_h_�_�_ �_�_�_�_
o�_o@o �Xojo|o&o�o�o�o �o�o�o*N` r�B����� ��&��6�\�J��� n�����ȏ��؏ڏ� "��F�4�j�X���|� ��ğ���֟���0� �@�B�T���x����� ү䯎o���̯ʯP� >�t�b����������� ���Կ&�L�:�p� ^ϔϦϸ��τ����� � �"�H�6�l�Zߐ� ~ߴߢ���������� 2� �V�D�z�h��� �����������
�,� .�@�v�������\� ������<*` N����x�� �8J\( �������� /4/"/X/F/|/j/�/ �/�/�/�/�/�/?? B?0?f?T?v?�?�?�? �?�?�?OO��2ODO �� O�OtO�O�O�O�O �O_�O(_:_L_
__ �_p_�_�_�_�_�_ o �_$oo4o6oHo~olo �o�o�o�o�o�o�o  D2hV�z� ����
��.�� R�@�b���v���&OXO ֏菒�����N�<� r�`�������̟ޟ� ����$�&�8�n��� ����^�ȯ���گ� �� �"�4�j�X���|� ����ֿĿ����0� �T�B�x�fψϊϜ� ����������>�P� ��h�zߌ�6߼ߪ��� �������:�(�^�p� ���R������� ����  &�*� �*�>�*��$TB�JOP_GRP �2U����  ?���KC*�	V�]�Wd������X  *���� �, � ���*� �@&�?��	 �A������C�  �DD�����>v�>�\? ��a�G�:�o��;ߴAT������A�<��MX�����>��\)?;���8Q�����L��>�0 &�;�iG.��Ap�< � F�A�ff��v��� ):VM�.�� S>�o*�@��R�Cр	��������ff�:�6�/�?�33�B   ��/������>):�S����� �/�/@��H�%&/�/�z�=� <#�
*���v�;/�ڪ!?���4B�3?'? 2	��2?hZ?D?R?�? �?�?F?�?�?�?�?O AOO�?`OzOdOrO�O,�O*�C�*���A��	V3.00{��crxl��*�P��%�%c5Z �F� JZH� F6� F^� F�� F�f� F� G�� G5 G<
� G^] G�� G���G�*��G�S G�;o G��ERDu��\E[� E�� F( F-�� FU` F} � F�N F�� F�� Fͺ� F� F�V� G� Gz� Ga 9ѷI�Q�LHefJ4�o,b*�0c1����OH�ED_TCH� Xd�+X2S�2&�&�d$'X�o��o*�1F�TES�TPARS  ���cV�HRpAB�LE 1Yd� AN`*�����g$j
�g�h�h)�1��g	�h
�h�hHu*�U�h�h�h%v'RDI0n�GY k}��u	�O�#�@-�?�Q�c�u�)rS�l� �z6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z���I� ��m�Fwͩ��ȏڏ 쏘�����x)r~��NUM  ��n���2� �Ep�)r_CFG �Z��I���@V�IMEBF_TTqtD��e޶VER������޳R 1[�8{ 8�o*�d%�Q� ��د  9� K�]�oρϓϥϷ��� �������#�5�G�Y� k�}��ߡ߳������� ����1���E�W�i� {������������ ��/�A�S�e�w��� �������������+=O�_���@���`LIF M\��D`�����DR�(FP
�:!p�!p� d� ��MI_CHAN�� � DBGL�VL��fET�HERAD ?u��0`1�_}��ROUT��!�j!��SNMASKY�j255.%S/�//A/S�`OOLO_FS_DIp��CORQCTRL� ]8{��1o�-T �/�/�/??+?=?O? a?s?�?�?�?�?�?�? �?OL�/6O%OZOc�PE_DETAI�7�*PGL_CONFIG c�������/cel�l/$CID$/grp1^O�O�O�O
__|���G_Y_k_ }_�_�_0_�_�_�_�_ oo�_CoUogoyo�o �o,o>o�o�o�o	 -�oQcu��� :�����)�� �_�q���������׮}N����%�7�I�a�KOq�P��M����� ʟܟ� �G�$�6�H� Z�l�~������Ưد ������2�D�V�h� z������¿Կ��� 
ϙ�.�@�R�d�vψ� ��)Ͼ��������� ��<�N�`�r߄ߖ�%� ����������&�� J�\�n����3��� �������"���F�X��j�|��������@��User Vi�ew �I}}12�34567890 ����+=Ex ,�e����2��B� �����`r��3�Oas����x4>//�'/9/K/]/�~/x5 ��/�/�/�/�/?p/2?x6�/k?}?�?�? �?�?$?�?x7Z?O 1OCOUOgOyO�?�Ox8O�O�O�O	__-_��ON_TR lCamera�� �O�_�_�_�_�_�_˂E�_o)o;n��Uogo`yo�o�o�o�)  mV �	�_�o#5GY  o}���o������F_�mV=� k�}�������ŏl� ���X�1�C�U�g�y� ��2�D��"�ן��� ��1�؏U�g�y�ğ ������ӯ�����D� �k��E�W�i�{����� F�ÿտ�2���/� A�S�e��nUY9���� ��������	߰�-�?� Qߜ�u߇ߙ߽߫��� v�D�If��-�?�Q� c�u�ߙ������ ����)�;���D��I ��������������� )t�M_q���N�`�93�� 0B��Sx� 1�����//
�J	oU0�U/g/y/ �/�/�/V�/�/�/� ?-???Q?c?u?/./ tPv[?�?�?�?OO (O�/LO^OpO�?�O�O �O�O�O�O�?oU�k�O :_L_^_p_�_�_;O�_ �_�_'_ oo$o6oHo Zo_;%N��_�o�o�o �o�o �_$6H�o l~����moe ��]�$�6�H�Z�l� �������؏��� � �2��e&�ɏ~� ������Ɵ؟����  �k�D�V�h�z����� E�e��5����� � 2�D��h�z���ׯ���¿Կ���
ϱ�  ��9�K�]�oρπ�ϥϷ���������   ��5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u����� ����������)�;M_q�  
���(  �-�( 	 ���� ���#35G@}k����
� �Y�
//./�� R/d/v/�/�/�/��� �/�/�/A/?0?B?T? f?x?�/�?�?�??�? �?OO,O>O�?bOtO �O�?�O�O�O�O�O_ KO]O:_L_^_�O�_�_ �_�_�_�_#_ oo$o k_HoZolo~o�o�o�_ �o�o�o1o 2D Vh�o�o���	 ��
��.�@��d� v��������Џ�� �M�*�<�N���r��� ������̟�%��� &�m�J�\�n������� �ȯگ�3��"�4� F�X�j����������� ֿ�����0�w��� f�xϊ�ѿ�������� ���O�,�>�Pߗ�t� �ߘߪ߼������� �]�:�L�^�p����߻@ ������������ ��"�frh:\tpg�l\robots�\crx!�10ia_l.xml�� D�V�h�z�������������������0 BTfx���� �����,>P bt������ ��/(/:/L/^/p/ �/�/�/�/�/�/��/ ?$?6?H?Z?l?~?�? �?�?�?�?�/�?O O 2ODOVOhOzO�O�O�O �O�O�?�O
__._@_ R_d_v_�_�_�_�_�_ �O�_oo*o<oNo`o ro�o�o�o�o�o�n ��6� ���<�< 	� ?� �k!�o;iOq �������� �%�S�9�k���o���裏я����(�$�TPGL_OUT?PUT f����w�� � &�8�J�\�n������� ��ȟڟ����"�4� F�X�j�|�������į��p�ր2345?678901��� ��1�C�K����r� ��������̿d�п� �&�8�J��}T�|� �Ϡϲ���\�n���� �0�B�T���bߊߜ� ������j�����,� >�P����߆���� ����x����(�:�L� ^���l����������� t���$6HZl z������ � 2DVh  �������/ ./@/R/d/v//�/�/��/�/�/�/�/ۂ $$��ί<7*? \?N?�?r?�?�?�?�? �?�?OO4O&OXOJO |OnO�O�O�O�O�O�O _�O0_"_T_}�an_@�_�_�_�_�_�]@��_o	z ( 	 V_Do2ohoVo�o zo�o�o�o�o�o
�o .R@vd�� �������(��*�<�r�`���ܦ� ? <<I_ˏ ݏ�������:�L� ֪��}���)���ş�� �����k��C�ݟ/� y���e���������� ���-�?��c�u�ӯ ]�����W���Ϳ�� )χ���_�q��yϧ� �ϓ�����M��%߿� �[�5�Gߑߣ�߫� ��s����!���E�W� ��?���9������ ���i���A�S���w� ��c�u����/��� ��=)s��� ��U���' 9�!o	[�� ���K�#/5/� Y/k/E/w/�/�/�/ �/�/�/?�/?U?g? �/�?�?7?�?�?�?�?�	OO��)WGL�1.XML�_PM��$TPOFF_L�IM ���P����^FN_SV�f@  �TxJP_MON g��SzD�P�P2ZI�STRTCHK �h��xFk_aBVTCOMPAT�H�Q|FVWVAR �i�M:X�D ��O R_�P�B�bA_DEFPRO�G %�I%?TELEOPi_�O�_DISPLAY�m@�N�RINST_�MSK  �\ ��ZINUSER�_�TLCKl�[QUICKMEN:o��TSCREY`���Rtpsc@�Tat`yixB�`_�i�STZxIRACE_CFG j�I�:T�@	[T
?���hHNL 2k�Z���aA[ gR-? Qcu����z�eITEM 2l{� �%$1234567890 ��  =<
�0�B�J�  !P�X�dP���[S���"�� �X�
�|���W���r� ֏����.��0�B�\� f�����6�\�n�ҟ�� ������>���"� ��.�����ίR���� Ŀֿ:��^�p�9ϔ� Tϸ�xϊ���d� ��H��l��>�Pߴ� \�������v� ����� �h�(�ߞ߰�4�L� �ߦ�����@�R�� v�6���Z�l������ ���*���N��� �� ����������X� ��J
n�� �b����"4 F�/|</N/�Z/ ���//�/0/�/? f/?�/�/e?�/�?�/ �?�?�?,?�?P?b?t? �?�?DOjO|O�?�OO O(O�O�O^O_0_�O <_�O�O�_�O�__�_��_H_�_l_~_Go�dS��bm�oLj�  �rLj �a�o�Y
 �o�o�o�o{j�UD1:\|���^aR_GRP �1n�{� 	 @�PRd{N� r����~��p����q+��O�:�?�  j�|�f����� �����ҏ����>� ,�b�P���t����������	e���\cS�CB 2ohk U�R�d�v��������Я�RlUTOR?IAL phk�o�-�WgV_CONFIG qhm�a�o��o��<�OUTPU�T rhi}�����ܿ� ��$� 6�H�Z�l�~ϐϢϴ� z�ɿ���� ��$�6� H�Z�l�~ߐߢߴ��� ������� �2�D�V� h�z���������� ��
��.�@�R�d�v� �������������� *<N`r�� ������& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/� �/�/??0?B?T?f? x?�?�?�?�?�/�?�? OO,O>OPObOtO�O �O�O�O�?�O�O__ (_:_L_^_p_�_�_�_ �_�_f�x�ǿoo,o >oPoboto�o�o�o�o �o�o�O(:L ^p������ �o ��$�6�H�Z�l� ~�������Ə؏�� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я����*�<� N�`�r���������̿ ޿���&�8�J�\� nπϒϤ϶������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ������������,� >�P�b�t�����������������X���#��N�_r ������� &8J��n�� ������/"/ 4/F/X/i|/�/�/�/ �/�/�/�/??0?B? T?e/x?�?�?�?�?�? �?�?OO,O>OPOa? tO�O�O�O�O�O�O�O __(_:_L_^_oO�_ �_�_�_�_�_�_ oo $o6oHoZok_~o�o�o �o�o�o�o�o 2 DVgoz���� ���
��.�@�R� d�u��������Џ� ���*�<�N�`�q� ��������̟ޟ����&�8�J�\�k��$�TX_SCREE�N 1s%; �}�k��� ��ӯ���	���Z ��I�[�m������� ,�ٿ����!�3Ϫ� W�ο{ύϟϱ����� L���p��/�A�S�e� w��� ߭߿������� �~�+��O�a�s�� ��� ���D����� '�9�K���������� ������R���v�#5�GYk}����$�UALRM_MS�G ?����� �n���	: -^Qc������� /�SEV � �2&�E�CFG u�����  n�@��  Ab!   B�n�
 /u��� �/�/�/�/�/�/??�%?7?I?W7>!GRPw 2vH+ 0n��	 /�?� I_�BBL_NOTE� wH*T���lu���w��T �2DEFPROz� %� (%� Ow�	OBO-OfOQO�O uO�O�O�O�O�O_�O�,_�<FKEYDA�TA 1x���0�p W'n�  U?�_�_�0_�_�_�U,(7_on��_7oo [oBoo�oxo�o�o�o �o�o�o3E,i P�������`���A�p^��Q� x���������ҏu�f� ����1�C�U��y� ��������ӟb���	� �-�?�Q�c�򟇯�� ����ϯ�p���)� ;�M�_�������� ˿ݿ�~��%�7�I� [�m����ϣϵ����� ��z��!�3�E�W�i� {�
ߟ߱��������� ���/�A�S�e�w�� ������������� +�=�O�a�s���\��� ��������
�'9 K]o��"�� ����5GY k}����� �//�C/U/g/y/ �/�/,/�/�/�/�/	? ?�/??Q?c?u?�?�? �?:?�?�?�?OO)O �?MO_OqO�O�O�O6O �O�O�O__%_7_�O [_m__�_�_�_D_�_ �_�_o!o3o�_Woio@{o�o�o�o�o���k���������o}�o8J$v, 6�{.������ ���/��S�:�w� ��p�����я�ʏ� �+��O�a�H���l� ������ߟ���'� 9�Ho]�o��������� ɯX�����#�5�G� ֯k�}�������ſT� �����1�C�U�� yϋϝϯ�����b��� 	��-�?�Q���u߇� �߽߫�����p��� )�;�M�_��߃��� ������l���%�7� I�[�m���������� ����z�!3EW i�������� �П/ASew ~������/ �+/=/O/a/s/�// �/�/�/�/�/?�/'? 9?K?]?o?�?�?"?�? �?�?�?�?O�?5OGO YOkO}O�OO�O�O�O �O�O__�OC_U_g_ y_�_�_,_�_�_�_�_ 	oo�_?oQocouo�o �o�o:o�o�o�o )�oM_q��� 6�����%�7��9�����b�t���^�������,��돞���� 3�E�,�i�P������� ß���������A� S�:�w�^�������ѯ ����ܯ�+�
O�a� s��������Ϳ߿� ��'�9�ȿ]�oρ� �ϥϷ�F�������� #�5���Y�k�}ߏߡ� ����T�������1� C���g�y������ P�����	��-�?�Q� ��u�����������^� ��);M��q ������l %7I[�� ����h�/!/ 3/E/W/i/@��/�/�/ �/�/�/�??/?A? S?e?w??�?�?�?�? �?�?�?O+O=OOOaO sOO�O�O�O�O�O�O _�O'_9_K_]_o_�_ _�_�_�_�_�_�_�_ #o5oGoYoko}o�oo �o�o�o�o�o�o1 CUgy��� ���	���?�Q� c�u�����(���Ϗ� �����;�M�_�q�Ѓ�����~ ���>~ ���ҟ� ��Ο�*��,�[� ��f�������ٯ�� �����3��W�i�P� ��t���ÿ���ο� �/�A�(�e�Lωϛ� z/����������(� =�O�a�s߅ߗߩ�8� ��������'��K� ]�o����4����� �����#�5���Y�k� }�������B������� 1��Ugy� ���P��	 -?�cu��� �L��//)/;/ M/�q/�/�/�/�/�/ Z/�/??%?7?I?�/ m??�?�?�?�?�?�� �?O!O3OEOWO^?{O �O�O�O�O�O�OvO_ _/_A_S_e_�O�_�_ �_�_�_�_r_oo+o =oOoaosoo�o�o�o �o�o�o�o'9K ]o�o����� ���#�5�G�Y�k� }������ŏ׏��� ���1�C�U�g�y��� �����ӟ���	��� -�?�Q�c�u���������ϯ�����0����0���B�T�f�>�����t�,��˿~��ֿ�%� �I�0�m��fϣϊ� ����������!�3�� W�>�{�bߟ߱ߘ��� ������?/�A�S�e� w���������� ����=�O�a�s��� ��&��������� ��9K]o��� 4����#� GYk}��0� ���//1/�U/ g/y/�/�/�/>/�/�/ �/	??-?�/Q?c?u? �?�?�?�?L?�?�?O O)O;O�?_OqO�O�O �O�OHO�O�O__%_ 7_I_ �m__�_�_�_ �_�O�_�_o!o3oEo Wo�_{o�o�o�o�o�o do�o/AS�o w������r ��+�=�O�a���� ������͏ߏn��� '�9�K�]�o������� ��ɟ۟�|��#�5� G�Y�k���������ů ׯ������1�C�U� g�y��������ӿ� �����-�?�Q�c�uϴ��^P���^P��������ͮ���
���,��;���_� F߃ߕ�|߹ߠ����� �����7�I�0�m�T� ������������ !��E�,�i�{�Z_�� �����������/ ASew��� ����+=O as����� �//�9/K/]/o/ �/�/"/�/�/�/�/�/ ?�/5?G?Y?k?}?�? �?0?�?�?�?�?OO �?COUOgOyO�O�O,O �O�O�O�O	__-_�O Q_c_u_�_�_�_:_�_ �_�_oo)o�_Mo_o qo�o�o�o�o���o�o %7>o[m ����V��� !�3�E��i�{����� ��ÏR������/� A�S��w��������� џ`�����+�=�O� ޟs���������ͯ߯ n���'�9�K�]�� ��������ɿۿj��� �#�5�G�Y�k����� �ϳ�������x��� 1�C�U�g��ϋߝ߯ߠ���������`��}��`���"�@4�F��h�z�T�,f� ��^���������)� �M�_�F���j����� ��������7 [B�x��� ��o!3EWi xߍ������ �///A/S/e/w// �/�/�/�/�/�/�/? +?=?O?a?s?�??�? �?�?�?�?O�?'O9O KO]OoO�OO�O�O�O �O�O�O_�O5_G_Y_ k_}_�__�_�_�_�_ �_o�_1oCoUogoyo �o�o,o�o�o�o�o	 �o?Qcu�� (������)�  M�_�q�������� ˏݏ���%�7�Ə [�m��������D�ٟ ����!�3�W�i� {�������ïR���� ��/�A�Яe�w��� ������N������ +�=�O�޿sυϗϩ� ����\�����'�9� K���o߁ߓߥ߷��� ��j����#�5�G�Y� ��}��������f� ����1�C�U�g�>��i��>������������������,��?&c u\������ �)M4q� j�����/� %//I/[/:�/�/�/ �/�/�/���/?!?3? E?W?i?�/�?�?�?�? �?�?v?OO/OAOSO eO�?�O�O�O�O�O�O �O�O_+_=_O_a_s_ _�_�_�_�_�_�_�_ o'o9oKo]ooo�oo �o�o�o�o�o�o�o# 5GYk}�� ������1�C� U�g�y��������ӏ ���	���-�?�Q�c� u�����p/��ϟ�� ���;�M�_�q��� ����6�˯ݯ��� %���I�[�m������ 2�ǿٿ����!�3� ¿W�i�{ύϟϱ�@� ��������/߾�S� e�w߉ߛ߭߿�N��� ����+�=���a�s� �����J������ �'�9�K���o����� ������X�����# 5G��k}���h�����������&�HZ4,F/�>/ �����	/�-/ ?/&/c/J/�/�/�/�/ �/�/�/�/?�/;?"? _?q?X?�?|?�?�?�� �?OO%O7OIOXmO O�O�O�O�O�OhO�O _!_3_E_W_�O{_�_ �_�_�_�_d_�_oo /oAoSoeo�_�o�o�o �o�o�oro+= Oa�o����� ����'�9�K�]� o��������ɏۏ� |��#�5�G�Y�k�}� �����şן����� �1�C�U�g�y���� ����ӯ���	��?-� ?�Q�c�u��������� Ͽ���Ϧ�;�M� _�qσϕ�$Ϲ����� ���ߢ�7�I�[�m� ߑߣ�2��������� �!��E�W�i�{�� ��.����������� /���S�e�w������� <�������+�� Oas����J ��'9�] o����F����/#/5/G/�$U�I_INUSER  ���h!��  �H/L/_MENH�IST 1yh%�  (�w  �(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1�/�/??f0?�)�/�/13�/ |?�?�?�?�'E?W>2k?�?O"O4O��/>�?148,29O�O�O�O�O���O�O�O __*_<_�O`_r_�_ �_�_�_I_�_�_oo &o8o�_Iono�o�o�o�o�o��\a�!\o�o /ASVow� ����`��� +�=�O��������� ��͏ߏn���'�9� K�]�쏁�������ɟ ۟j�|��#�5�G�Y� k���������ůׯ� �o�o�1�C�U�g�y� |�������ӿ����� �-�?�Q�c�uχ�� �Ͻ�������ߔ�)� ;�M�_�q߃�ߧ߹� ���������7�I� [�m��� ������ ��������E�W�i� {��������������� ��ASew� ��<��� +�Oas��� 8���//'/9/ �]/o/�/�/�/�/F/ �/�/�/?#?5? �2� k?}?�?�?�?�?�/�? �?OO1OCO�?�?yO �O�O�O�O�ObO�O	_ _-_?_Q_�Ou_�_�_ �_�_�_^_p_oo)o ;oMo_o�_�o�o�o�o �o�olo%7I�[F?��$UI_�PANEDATA 1{����q�  	��}  frh/�cgtp/fle�xdev.stm�?_width=�0&_heigh�t=10�p�pic�e=TP&_li�nes=15&_�columns=�4�pfont=2�4&_page=whole�pmI6?)  rim�9�  �pP�b�t����� �������Ǐ��(� :�!�^�E�����{������ܟ�՟�I6� X14�G�L�^�p� ��������ʯ=�ܯ � �$�6�H�Z���~�e� ������ؿ����� � 2��V�=�zό�sϰ�#��Ɠs����� )�;�Mߠ�q�䯕ߧ� ��������V��%�� I�0�m��f����� ��������!��E�W� ���ύ����������� :�~�/ASew ������  =$asZ� ~����d�v�'/ 9/K/]/o/�/��/�/ *�/�/�/?#?5?�/ Y?@?}?�?v?�?�?�? �?�?O�?1OCO*OgO NO�O�/�/�O�O�O 	__-_�OQ_�/u_�_ �_�_�_�_6_�_o�_ )ooMo_oFo�ojo�o �o�o�o�o�o%7 �O�Om���� �^_�!�3�E�W� i�{������Ï��� ������A�S�:�w� ^�������џDV� �+�=�O�a������� 
���ͯ߯���|� 9� �]�o�V���z��� ɿ���Կ�#�
�G�0.�k�ޟ�}�|ϵ� ���������)��4� ��#�`�r߄ߖߨߺ� !����������8�� \�C���y������������������$�UI_POSTY�PE  ��� 	 ��s�B�QUICKM_EN  Q�`��v�D�RESTOR�E 1|��  ��B����������m ASew�,�� ����+=O an���� �//�9/K/]/o/ �/�/6/�/�/�/�/�/ �??0?�/k?}?�? �?�?V?�?�?�?OO �?COUOgOyO�O6?@O �O�O.O�O	__-_?_ Q_�Ou_�_�_�_�_`_ �_�_oo)o�O6oHo Zo�_�o�o�o�o�o�o %7I[�o�������SCR�E��?���u1sc��u2��3�4�5�6��7�8��sTATM�� ����:��USER�p��rTL�p�ks���4��U5��6��7��8���B�NDO_CFG� }Q�����B�P�DE����None��v�_I�NFO 2~��)���0%�D��� 2�s�V�������͟ߟ ��'�9��]�o��R���z��OFFS�ET �Q�-� ��hs��p����� G�>�P�}�t���Я�� ׿ο����C�:πL�^Ϩ����͘���
����av��WOR/K �!������.�@ߢ�u�UFRAME  ����RTOL_ABRqT�����ENB��~��GRP 1������Cz  A� �����*�<�N� `�r��֐�U���~��MSK  մ)���N��%!���%z����_EVNı����+�ׂ3��«
 h�U�EV��!td:�\event_u�ser\�u�C7�z���jpF��n�SP�s�x�spotw�eld��!C6 ��������!��� G|'��5kY� ����>�� �1�Ug�� �/��	/^/M/�/ -/?/�/c/�/�/�/�/@$?�/H?�/:J�W�33�����8C?�?�? �?�?�?�?O+O OOOaO<O�O�OrO�O �O�O�O_�O'_9__�]_o_J_�_�_�_�$�VALD_CPC� 2�« 8�_�_� w��q�d�R�*o_oqo��hsNbd�j�`��i�da{ �oav�_�ooo3Bo Wi{�o�o�o�o� �o�PA�0�e� w�������� ��(�=�L�a�s�
� ������ʏ����� $�ޟH�:�o������� ��ڟ؟����� �2� G�V�k�}�������¯ ԯ�����.��R� S�yϋϚ�������� ��	��*�<�Q�`�u� �ߖϨϺ�������� �&�8�M�\�q��� �߶���n������"� 4�F�[�j������� ���������!0�B� Wf�{�������� ���,>te T������� /+/:La/p�/ �/./�����// '?6/H/?l/^?�?�? �/�/�/�/�/?#O�? D?V?kOz?�O�O�?�? �?�?�?_O1_@ORO 9_vOw_�_�_�O�O�O _�__-o<_N_`_uo �_�o�o�_�_�_�_o &o;Jo\oq�o� ���o�o�o� �" 7�FXj������ �����!�0�E� T�f�{�������ßҏ ����
�,�A�P�b� ����x�����Ο��� ��(�*�O�^�p��� ������R�ܯ� �� Ϳ6�K�Z�l�&ϐ��� ����ؿ���"� �2� G���h�zϏߞϳ��� ������
��1�@�U� d�v�]�ߛ������� ���,��<�Q�`�r� ������������� �&�;J�_n���� ���������� $F[j|��� ����0E/ Ti/x��/��/�/ �/�//,/.?P/e? t/�/�/�?�?�?�?�/ ??(?:?L?NOsO�? �?�O�?�O�OvO OO $O6O�OZOo_~O�OJ_ �O�_�_�_�O_ _F_�D_V[�$VARS�_CONFIG ���Pxa�  FP]S��\lCMR_GR�P 2�xk� ha	`�`  %�1: SC13?0EF2 *�o�`�]T�VU�P�h`��5_Pa?�  �A@%pp*`�Vn No9xCVXd�v��a��<uA)�%p�q�_R���_R B��� #�_Q'��H��l�;� ��{�����؏ÏՏ� e��D�/�A�z�-������ddIA_WOR�K �xeܐ<�Pf,		�Qxe|���G�P ����YǑRTSYNC�SET  xi��xa-�WINURLg ?=�`������������ȯگSIONTMOU9��]Sd� ��_�CFG �S����S۵P~�` FR:\���\DATA\� �� MC3��LOG@�   7UD13�EXd�_Q�' B@ ����x�e_ſx�ɿ��VW � n6  ���VV�l�q  =����?�]T<�y�>Y�TRAIN���6N� 
gp?�C�D���TK���b�xk (g�����_��� ������U�C�y�g߀�ߋߝ߯������_�GE��xk�`�_P�
�P�RꋰR�E��xe*�`hLE�X�xl`1-e��VMPHASE'  xec�ec�RTD_FILT�ER 2�xk �u�0����0� B�T�f�x�����VW�� ������ $6H�Zl_iSHIFTMENU 1�xk/
 <�\%���������� =&sJ\��������'/��	LIVE/SN�A�c%vsflsiv��9/���� 7�U�`\"menur/w//�/�/������]��MO���y��5`h`ZD4��V�_Q<��0��$W�AITDINEN�D��a2p6OK C �i�<���?S�?�9TIM�����<Gw?M�?*K�?
J��?
J�?�8RELE���:G6p3���r1_�ACTO 9Hܑ�8_n<� �ԙ�%�/x:_af�BRDIS�`~�N�$XVR���y��$ZAB�C�b1�S; ,��j�I�2B_ZmI1��@VSPT ��y��eG�
�*��/o�*!o7o�WDCSCHG �ԛ�(��P\g@�PI-PL2�S?i��o��o�o�ZMPCF_OG 1��ii�0'� �S;Ms�S��i���p'��g��e2���g0���?�蕼�Ĕ?�啼�m<���i<��J����V��RD��@BQs�A���*I�?�q>�:�8>�s����=Z�׿2n?�����0����?�Z�~����Ï�>�C2��/?��kB��ڏ�ӈ������*�@�N�x��/�	�?����K����/$E;��^�;�!������UB���j��c�A��8I�0��?��)��M8���=EvϾ>Z ?d��glp����o�_CYLI�ND�� { ���� ,(  * =�N�G�:�w�^����� ��ѯ���7�� ��<�#�5�r������� ����޿y�_����8�@ύ�nπ�㜻ã wQ �5�����S �����(�ٻ�X���r�A��SPH�ERE 2��� ҿ��"ϧ������P� c�>�P�̿t���ߪ� �����'���]�o� L���p�W�i�������������PZZ�F � 6