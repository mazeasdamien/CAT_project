��   K�A��*SYST�EM*��V9.4�0107 7/�23/2021 A 	  ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_���$$�CLASS  O�����D���DVERSIO�N  �XK/IRTU�AL-9LOO�R G��DD<x$?�������k,  1 <DwX< y�����D@����	/��Z�Zm//��/_/�/�/�/$ ��/�/	?';�$M�NU>A\"�  <�?/o?��[?}? �?�?�?�?�?�?O�? O1O_OEOgO�O{O�O �O�O�O�O_�O_I_��;5NUM  ������92TOO=LC?\ 
Y?[_ �_3_�_o�_�_;o!o 3oUo�oio�o�o�o�o �o�o�o	7?m Se�����oZ �Q�Vy�Wy