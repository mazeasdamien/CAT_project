��   ��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����CCSCB2�_GRP_T � h $CO�MPMATEXP_1  :2F	�RIXU   d?$OFFSEAFGAGEsm;f�z� z_OKRGf � ��P��H FS_TYTS�BFRAMEe�$INIT_TO�L�RANGE2�_Ff�T�F�TRATIOe|� �H_LIMU��LFSOF�ST_S�mUP�S_����	e� O�L_{UDUMM�Y2U�3�����$$CLA�SS  �������I��I�V�ERSION��  XK~�IRTUAL�ܻ' 3 �I�/ ���d"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B?�T?f?x?�?�?�� �?�  �?�7:׃o�0���@o  'Bd����0@��0 �?F xA1E-AC�  AE��0�0�0W@�BpGO�;tO��FP��