��   �c�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����DCSS_C�PC_T 4 �$COMMEN�T $EN�ABLE  �$MODJGRP�_NUMKL\�  $UFR�M\] _VTX �M �   $�Y�Z1K $Z�2�STOP_T�YPKDSBIO�IDXKENBL_CALMD��USE_PRED�IC? �ELAY�_TIMJSPEED_CTRLKOVR_LIM? *p D� �L�0�UT�OOi��O���&S. ǰ 8J\TC �u
!���\�� jY0 � � �CHG�_SIZ�$A�P!�E�DIS"�]$!�C_+{#�s%O#J�p 	]$J d#� �&s"�"{#�)�$��'�_SEEX�PAN#N�iG�STAT/ D�FP_BASE_ $0K$4�!� .6_V7>H�73hJ- � q}�\AXS\3UP�LW�7����a7r � < w?�?�?��?�?�x//	7ELEM/ T �&B.2�NO�G]@%CNHA��DF#� $DAT�A)he0  �PJ�@ 2� 
&P5 �� 1U*n   �_VSiSZbRj0jR(��VyT(�R%S{TR/OBOT�X�SAR�o�U�V$CUR�_��R &SET�U4"	 $�d P_MGN�I?NP_ASSe#� PB!� `CiH�77`e��.fXc1�CONFIG_CHK`E�_PO* }dSHR�ST�gM^#/eOT�HERRBT�j_G]�R�dTv �ku>�dVALD_7h�e,�4hT1r
0R HpLHt� 0  lt<8NerRFYhH~tD�5�1� ��W��_A$R�jSPH/ (G%QПQ�Q3?wBOX/ 8�@F!��F!�G �r��zTU�IRi@  ,��F�pER%@2� $�p �l�_Sf�A�ZN>/ 0 IF1(@�p��Z_�0��_�0?wu0  @��QWyv	*��~����$$CL`  O���!���Q���Q�VERSIO�N�  �XK2�IRTU�AL�0�' 2 �?�Q  ((�����&@^����P����ϟ��������d<�9�Cz  P�8���a��� ������ׯ���� �.�@�R�d�f����� �������Կ	��*� <�N�`�r����ϫϺ� ̿����߮�8�J� \�n�)ߒϧ߶��ς� �����%�4�F�X�~� |ߎߣ�.��������� �!�0�B�T�f�x�� ������������ />�P�b���v��� �������+: L^p����� �� /'/9/HZ l/�/��/��� �//#?5?D/V/h/z/ �/�?�/�?�/�/�?
? O1OCOR?d?v?�?�O �?�O�?�?O	_�O-_ ?_NO`OrO�O�O�O�_ �_�O�Oo_)o;o�_ \_n_�_�_Mo�_�o�_ �_�oo7IXojo |o�o�o�o�R�o�o �3�E�Tfx� ����Տ��ݏ� �A�S�b�t������� ��џ�����(�=� O�^�p���������ʟ ߯� ��$�9�K�]� l�~���6���Ưۿ� ���#�2�G�Y�h�z� ��������Կ����
� �.�C�U�g�vψϚ� �Ϯ��������<�-� �Q�c�r߄ߖߨߺ� ��������)�8�M� _�������q��� �������4�&[m |������������v 3BWix� ������ />?/e/w/��� ��/��///(/=? L/a?s?�/�/�/�/�/ �?�/O?$?9OH?]O oO�O�?�?�?ZO�O�? �OO O2OG_VOk_}_ �O�O�O�O�O�_�Oo _._CoR_goyo�o�_ �_�_�_�o�_	o*o `oQ@u��o�o�o �o�o�o��&8M� \q�������� ����"�4��X�J� �������ď������$DCSS_C?SC 25���Q  P�;���Z���~�A� ����w�د������ � �D�V��z�=���a� ¿��濩����߿@� �d�'ψ�KϬϾρ� �ϥ����*���N�� r߄�Gߨ�k��ߏ��� ���&���J��n�1� ��U��y������~�GRP 2�' ����	�s� ^��������������� '��7]H�l ������� 5 2kV�z� �����/
/// U/@/y/d/�/�/�/�/ �/�/	?�/-??*?c? N?�?r?�?�?�?�?�? �?OO'OMO8OqO\O �O�O�O�O�O�O_�O %__"_[_F__�_�_ n_�_�_�_�_o�_o�Eo0oio�_GST�AT 2�E�ߜ< 6�?5����3|X=��x��2�.�6��C��6C=����6u�~��`C� �B�?��C���X`�<�fc>>���K��74����?�  �a��`4��Z����e�����$�[�?��b_����ޗ����y�\4���x�!D0�P y>/��S=��?{�.����T�`����9�^�#���U[>E���Pbth�>T_?z�"�p%�p�R�p�>�oh��b�=2wC�ϢCWmD��� y?aW�>�x�=���߾�oi?�p�2�v������w�[?�a���`�Dc�z�o�o �l��\�n��P��� ����Џ����jp�� ����z!�O�5�G�i� k�}���͟��՟�� ����ŏ{������� ï��������O�5� c�-�k�Q�c������� ���Ͽ����9� g�i����ۯ������ ���'��/�]��E� �ߥ�?����ߵ���� ����G�Y�3�}��i� {����������1� C��/�y�o߁߯��� [���������-? cuO����� ��)5_9 K������w� /%/�I/[/5/c/�/ k/}/�/�/�/�/?�/ ?E??1?{?�?g?�? �?�?�?�?��?/OAO �?eOwOQOcO�O�O�O �O�O�O_+___a_ ;_M_�_�_�_�_�_�_ �_oOOKo]o�_io �omoo�o�o�o�o �oG!3}�i �������1� C�9oG�y��e����� �����я��-��� c�u�O���������� ��͟�)��M�_�9� g���O�}�˯ݯw�� ����I�#�5���� k���ǿ������׿� 3�E��i�{�U�gϱ� �������ϓ��/�	� �e�w�Qߛ߭߇߹� �߽����+��O�a� ;�m��q�������� ������K�]�7��� ��m����������� ��5G!O}Wi ������1 ��gy��� ����/-//Q/ c/=/O/�/s/�/�/�/ �/??�/?M?CU �?�?/?�?�?�?�?O O�?7OIO#OUOOYO kO�O�O�O�O�O�O	_ 3___i_{_q?_�_ K_�_�_�_�_o/o	o 7oeo?oQo�o�o�o�o �o�o�o�oOa ;��q���_� ���9�K�%�7��� [�m���ɏ�����ُ �5��!�k�}�W��� ����������1� ˟=�g�A�S������� ӯ寿������Q� c�=�����s���Ͽ�� ������M��9� �ϕ�oϹ��ϥ���� ����7�I�#�m��Y� �ߵߏߡ�������!� 3��;�i�#�Q��� K������������	� S�e�?�����u����� ������=O) ;�{���g� ��9K%o� [������� #/5//A/k/E/W/�/ �/��/�/�/�/?1? ?U?g?A?o?�?w?�? �?�?�?	OO�?#OQO +O=O�O�OsO�O�O�O �O_�/�O;_M_�Oq_ �_]_o_�_�_�_�_o �_%o7oo#omoGoYo �o�o�o�o�o�o�o! _)_Wiu�y �������)� S�-�?�����u���я ��ݏ���=�O�E S����q���͟��� �ݟ�9��%�o��� [����������ǯٯ�#�5��Y�k�a��$�DCSS_JPC� 2`�Q? ( DQ�����ʴԿذ����ʿ ܿ1� ��$�y�Hχ� l��ϐ��ϴ�	����� ,�Q� �2߇�V�h�z� �ߞ��������;�
� _�.�@��d�v���� ������%���I��m� <�N������������� ����3W&{J �n������ �AO4�X� |����/�� O//0/B/�/f/�/�/ �/�/?�/'?�/?]? ,?>?P?�?t?�?�?�? �?O�?5OOOXO}O LO^O�O�O�O�O�O�O _�OC__g_6_�_Z_ l_�_�_�_�_	o�_oT4c��S����Louo&o�o�`ddo�o�o �o�o	�o-�oQ u<�`r��� ���;��_�&��� J���n�ˏ��ُ��� ڏ����m�4���X� ��|�ٟ����ğ!�� E���0�y���f�ï ��篮��ү/���S� �w�>���b������� ������=��a�(� ��Lϩ�p��ϔ��ϸ� ����%�K��o�6ߓ� Z߷�~��ߢ�����#� ��1��k�2�D�V�h� ���������1��� U��y�@���d�v��� ��������?c *�N�r��� ���q8 �\����/��%/�FdMODELw 2Skx��o(
 <o$c (/  o&�(�/ �/�/�/�/�/�/�/? ?d?;?M?�?q?�?�? �?�?�?O�?ONO%O 7OIO[OmOO�_�Oy/ �O�O&_�O_\_3_E_ W_�_{_�_�_�_�_o �_�_oXo/oAo�oeo wo�o�o�o�o�o�o �O�O�O/�� �������P� '�9�K�]�o���Ώ�� ���ۏ����#�5� ��Y�k���Se���� �������1�C��� g�y�Ư������ӯ� ��D��-�z�Q�c�u� ��������Ͽ�.�ɟ ۟	�ψ��qσ��� �Ϲ������<��%� 7߄�[�mߺߑߣ��� ������8��!�n�E� W��?�Q�cϑ��y� ����F��/�|�S�e� w�������������0 +=Oa�� �������>�� �]o��� �����/#/p/ G/Y/�/}/�/�/�/�/ �/$?�/?Z?1?C?U? +�?O}?�?�?�?�? 2O	OOhO?OQOcO�O �O�O�O�O�O_�O_ _d_;_M_�_q_�_�_ �_�_�_�?*o�?�_o roIo[o�oo�o�o�o �o�o&�o\3E Wi{����� ����/�A�o�� ;oi�{�菿�я��� ��+�=�O���s��� ҟ����͟ߟ��P� '�9���]�o������� �������߯�^�5� G���k�}���ܿ��ſ ����H��1�Cϐ� g�y��ϝϯ������� ��D��-���'�U� g���O߽�������� R�)�;��_�q��� ��������<��%� 7�I�[�m��������� �ߝ�����J��3E Wi{����� ��/|Se �������0/ //f/A/S/�/ ;/�/�/?�/�/>?? '?t?K?]?o?�?�?�? �?�?�?(O�?O#OpO GOYO�O}O�O�Ow/�/ �/�O�O�O_1_~_U_ g_�_�_�_�_�_�_�_ 2o	ooho?oQocouo �o�o�o�o�o�o �Ov_?Q'� ����*���%� 7�I�[������ޏ�� Ǐُ����\�3�E����i�{���Җ�$D�CSS_PSTA�T �����Q   g �� �� (&�K�2�o���� ������$�˟į֯���� ������'��SETUPw 	�Bȶ���X�r����������ۿ�g��T1�SC 2
K����Cz�#�5�G� ��CP R�D$�Dl�Ϥ�^���� �ϻ��"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x�� ������������� ,�>�P�b�t������� ��������(: L^p����~� �����-�Q cu������ �//)/;/M/_/q/ �/�/�/�/�/�/�/? ?%?7?I?[?m??�? �?�?�?�?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�__/_B S_e_w_F_�_�_�_�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9K]o� �������� #�5�G�Y�k�}����� ��ŏ׏�����1�  _U�g�y��_������ �����	��-�?�Q� c�u���������ϯ� ���)�;�M�_�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�W�i�{�J��߱� ğ���������/�A� S�e�w������� ������+�=�O�a� s��������������� '9K]o� ������� #5GYk}�� �������/1/ C//g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_�!o 3oEoX/io{o�o\o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�ok�}��o^� ��ů�������1� C�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m�����$DCSS_T�CPMAP  �������Q @ ��J���������U������	��U
��������u��W�  ��U�������������⡋��������������� ��!��"���#��$��%��&���'��(��)��*���+��,��-��.���/��0��1��2���3��4��5��6���7��8��9��:���;��<��=��>��?��@��UIR�O 2�����������0 BTfx��������,1 ��U��y���� ���	//-/?/Q/ c/u/�/�/�/6�/Z �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7O�/[O�/O�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_�_��_NO�_��UIZNw 2��	 �����(o:oLoR�%ozo �o�oao�o�o�o�o
 .�oRdvE� �������*� <�N�`�#�����e��� ̏ޏ�����&�8�� \�n���C�����ȟ�� ����ӟ4�F�X�'� |�����c�u�֯请����0��_��UFRwM R����� ��w���������ѿ� ����+�=�O�a�s� �ϗϩϻ����������'�9�K�\�r�� \߄ߖ�qߺ��ߧ��� ���&�8��\�n�I� ������������ ��4�F�]�o�|���-� ������������0 TfA��w� ����>P g�t�%���� ��/(//L/^/9/ o/�/�/�/�/�/�/ ? ?�/6?H?_l?~?? �?�?�?�?�?�?�? O 2OOVOhOCO�O�OyO �O�O�O�O
_�O._@_ W?d_v__�_�_�_�_ �_�_�_o*ooNo`o ;o�o�oqo�o�o�o�o �o&8O_!n� ������� "��F�X�3�|���i� ��ď�����Տ�0� B�Yf�x�������� ҟ䟿�����>�P� +�t���a�����ί�� ��߯(�:�@�