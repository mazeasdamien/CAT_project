��   ��A��*SYST�EM*��V9.4�0107 7/�23/2021 A 
  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41p� d =R��&�J_  4 �$(F3IDX؞�_ICI��?�MIX_BG�-y
_NAM�c MODc_U�Sd�IFY_T�I� ��MK�R-  $�LINc   "_SIZcg��� �. h $USE_FL�C 3!�:&iF*SIAMA7#QC#QBn'oSCAN�AX�+�IN�*I��_COUNrRO( ��!_TMR_VA�g#h>�i a �'` ����1n�+WAR�$�iH�!�#N3CH��PE�$O�!PR"�'Ioq7iOqf�OoATH- �P $ENABL+�0BT�f�$$CLAS�S  ����A��5��5�0VE�RS�G�  XKAIRTU� O@'/ @E_5�������-@{FA@A�E��%A�O���O�O�����QEI2\K �O;_M___q_�_ �_�_�_�_�_�_oo�%o7oIo�O)W?<"Hg@ ���j�@�o�o�i�� � �2\I  4%Xo��}A�A�o ;_qP������@�A���� 8��)�n�M�A@�c$"P+ �k�K-@��ń�AЄX�A@A-@�N ��
��.�@�R�d�v� ��������П���F�A 偍A��(�:�L�^� p���������ʯܯ�dDxMsW� 2���h�O�a�s��� ������Ϳ߿��� '��A�Z�l�~ϐϢ� ����������� �2� =�V�h�zߌߞ߰��� ������
��.�@�K� d�v��������� ����*�<�G�Y�r� �������������� &8JU�n�� ������" 4FXc|��� ����//0/B/ T/_q�/�/�/�/�/ �/�/??,?>?P?b? ah�4�0���?�p