��   g�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����BIN_CF�G_TX 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG���DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST��NSS�* 8�D�FACE_NUM? �$DBG_LE�VEL�OM_N�AM� !� FTޒ @� LOsG_8	,CMO>�$DNLD_F�ILTER�SUBDIRCAPCp��8 . 4� �H{ADDRT�YP�H NGT1H�� �z +�LSq D $ROBOTIG ��PEER�� MwASK�MRU~�OMGDEV�.�TP�PINFO~�  $�$$TI ���RCM+�T A$( /�Q�SIZ�!S� T�ATUS_%$MAILSERV� $PLAN� �<$LIN<$�CLU��<$T�O�P$CC�&F�R�&YJEC|!�Z%ENB � A�LAR:!B�TP�,�#,V8 S���$VAR�)M�O�N�&���&APPL��&PA� �%��'P�OR�Y#_�!�"A�LERT�&i2UR�L }Z3AT�TAC��0ERR�_THROU3US0�9H!�8� CH- c%�4MAX?WS_�|1��1MOD��1I�  �1o }(�1PWD  � cLA��0�ND�1�TRYFDELA�-C�0G'AERSI���1Q'ROBICL�K_HM 0Q'� XM�L+ 3SGFRM2U3T� !OUU3 3G_�-COP1�F�33�AQ'C[2�%�B_AU�� 9 R�!�UPDb&PCOU�{!�CFO 2 
$V*W�@c%�ACC_HYQSNA��UMMY1oW2�"$DM*  �$DIS��S=M	 l5��o!�"%Q7�IZP�%H� �VR�0�UP� �_DLVSPAR���QN,#
3 ��_�R!_WI�CT?Z_INDE�3^`gOFF� ~URmi�D�)c�  � t Z!`MO�N��cD��bHOUU#E%A�f�a�f�a��fLOCA� #{$NS0H_HE����@I�/  �d8`ARPH&�_7IPF�W_* O2�F``QFAsD90�VHO_� 5R42�PSWq?�TEL�� P��\�90WORAXQ�E� LV�[R2��ICE��p� ��$cs  ��)��q��
��
�p�PyS�A�w# kXK	�Iz0AL���' �
���F�����!�p�i��]$� 2Q��P ��������� Q���!�q����$� _?FLTR  �\�W �������!���$Q�2��7r{SH`D 1Q�E P㏙�f��� ş��韬��П1��� =��f���N���r�ӯ �������ޯ�Q�� u�8���\�������� ���ڿ;���_�"�X� �τϹ�|��Ϡ���� ���6�[���Bߣ� f��ߊ��߮���!��� E��i�,��P�b��� ��������/���(��e�T���L�����z _�LUA1�x!�1.��0��p���1|��p�255.0L��r��n���2�����d %7I[3 e��� ����[4���T'9[5U���{���[6���D �/�/)/s��Qȁ�a��a�P������ OQ� ��u.<�/ ?&?�/J?\?n?A?�?�?m�P�?�?�?�?�? O.O@OROOvO�O�O�u.kOl�q��O�L�
ZDT StatusZO�O5_G_Y_�n�}iRCon�nect: ir�c{T//alert^�_�_�_�_mW#_�oo,o>oPobot�2^�P~2g���go�o �o�o�o�o�o	-�?Qcul�$$c�962b37a-�1ac0-eb2�a-f1c7-8�c6eb5138?a8c  (�_�@_���"�p�1!
W��(��"S��JE�`� X��C� ��,$� ��W���ˏ���֏ ��%��I�0�m��f� ����ǟ�������!�4�u�R����� 7DM_�!�����SMTP_CTR�L 	����% ����DF���ۯt�ʯ ��'��Lz�N��!�
j��y�q�u�����Ԙ��#L�USTOM j�2�����  ���$_TCPIPd�j�a�H�%�"�EL������!���H!�T�b<�n�rj_3_tpd7� ��~i�!KCLG��L�i���5�!CR�T�ϔ����"u�!�CONS��M��[�ib_smon����