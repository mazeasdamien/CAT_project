��   g�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����BIN_CF�G_TX 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG���DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST��NSS�* 8�D�FACE_NUM? �$DBG_LE�VEL�OM_N�AM� !� FTޒ @� LOsG_8	,CMO>�$DNLD_F�ILTER�SUBDIRCAPCp��8 . 4� �H{ADDRT�YP�H NGT1H����z +�LSq D $ROBOTIG ��PEER�� MwASK�MRU~;OMGDEV���PINFO. �  $$$�TI ��R�CM+T �A$( /�QSI�Z�!S� TAT�US_%$MAI�LSERV $�PLAN� <$�LIN<$CLyU��<$TO�oP$CC�&FR�&�YJEC|!Z%E�NB � ALA5R:!B�TP,�#�,V8 S��$VkAR�)M�ON�&����&APPL�&P�A� �%��'POR��Y#_�!�"ALE�RT�&i2URL �}Z3ATTA�C��0ERR_T7HROU3US�9H!��8� CH- c%�4M�AX?WS_|1;��1MOD��1AI�  �1o (�1�PWD  � LAط�0�ND�1TR=YFDELA-C�0<G'AERSI��1vQ'ROBICLK_HqM 0Q'� XML+ �3SGFRMU3T̑ !OUU3 G_�-COP1�F33�A�Q'C[2�%�B_AU��� 9 R�!UP=Db&PCOU{!�C�FO 3 
�$V*W�@c%AC�C_HYQSNA�U�MMY1oW2"$D�M*  $gDIS��SM	 l5�o!�"!%Q7�IZP�%� ��VR�0�UP� _D�LVSPAR��?�SN,
�3 �_�R!_WI��CTZ_INDE��3^`OFF� ~U�RmiD�)c�  ? t Z!`'MON��cD��bHOUU#E%A�f�ax�f�a�fLOCA� �#$NS0H_H-E���@I�/ w d8`ARPH&��_IPF�W_�* O�F``QFApsD90�VHO_� �5R42PSWq?�T;EL� P��r�90WORA5XQE� LV�[:R2�ICE��p�� �$cs  �����q��
��
��p�PS�A�w�# XK	�Iz0A�L��' �
�
��F����!�p�i�w�$� 2Q��P��������� �Q���!�q����$�� _FLTR  \�\� �����������$Q�2���7rSH`D 1Q� P㏙�f���ş��韬��П 1���=��f���N��� r�ӯ�������ޯ� Q��u�8���\����� ��󿶿�ڿ;���_� "�XϕτϹ�|��Ϡ� ������6�[��� Bߣ�f��ߊ��߮��� !���E��i�,��P� b����������/� ��(�e�T���L������z _LUA1�x/!1.��0��p����1��p�2551.0��r��n���2����d %7I[3e��� ����[4���T'9[5U���{���[6���D  �//)/s��Qȁ�MA��MA��P����?� Q� ��u.<�/?&?�/J?\?n?A?�?�?m�P�?�?�? �?�?O.O@OROOvO�O�Ou.kOl�q��O��L
ZDT StatusZO�O5_�G_Y_n�}iRC�onnect: �irc{T//alert^�_�_�_�_ mW#_oo,o>oPobo�t�^�P~2g��� go�o�o�o�o�o�o	�-?Qcul�$�$c962b37�a-1ac0-e�b2a-f1c7�-8c6eb56�401a8  ( �_�_���"�p�)1!W��(��"S�`�JE�� X��tQ���,$���W���ˏ ���֏��%��I�0� m��f�����ǟ��������!��u�R������ DM_�!�����SMTP_CTRL 	����%����DF��� ۯt�ʯ��'��Lz�N�� 
j��y��q�u���������#L�USTOM' j������ � ���$TCPIPd�j��H�%�"��EL�����!���H!T�b<�n��rj3_tp�d7� ��i�!KCLG�L�i���5�!CRT�ϔ�����"u�!CON�S��M�[�ib_Osmon����