��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1CES0�2eG ��  QA> �1
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1�TU4QQ_M�AR�x1R� � /$TIT91� �� � �Td�T0�ThP�TU5�V6�V7�V8�V9�W0�W�WOQ�U�W�gQ�U�W1�W1�W1��W1�W2�R!SBoN_CF�!@$<!J� ; ;2�1�_CMNT�$�FLAGS]�C�HEK"$�b_O�PTJB � ELL�SETUP � `@HO8@9 P�R�1%�c#�aREPR�hu0D+�@���b{uHM9 MN�B;1�@UTOB�J U�0 }49DEVIC�STI/@�� �@b3�4pB�d�"VAL��#ISP_UNI�tp_DOcv7�yFR_F�@|%u13���A0s�C_WAx�t,q�zOFF_T@]N�DEL�Lw0pdq�1�Vr?^q��#S?�o`Q"U��t#*�QTB����MO� �E 	� [M�����wREV�BIL��͋� XI� v�R / !D�`���$NOc`M@�|����ɂ/#`ǆ� ԅ�������@Ded p �E RD_E��h��$FSSB6�`K�BD_SE�uAG*� G�2Q"_��2b�� V!�k5p`(��C��00q_ED� �� � t2�$!SL�p-D%$� �#r�B�ʀ_OK1��0] P_C� ʑ0tx��U �`LACI�!��a�Y�� �qCOsMM� # $D
�� ��@���J_\R BIGALLOW�G (Ku2-B�@�VAR���!�AB ��*�BL�@� �C ,K�q���`S�p��@M_O]˥���CCFS_UT��0 "�A�Cp'���+pXG��b�0 4�� IMCM ��#S@�p�9���i �_��"t�C��M�1 �h$�IMPEE_F�s��s��� t�����D_�����DR��F����_����0 T@L���L�DI�s@G�� ��P�$�I�'�� �CFned X@GRU@���Mb�NFLIx�\Ì@UIRE�xi42� SWITn$�`0_N�`S 2CFz�0M� �#u�D��!��v`���J�`J�tV��[ E���.p�`�ʗELBOF� �շ�p@`0���3����� F�2�T��A`�rq1J1,��z _To!��pЩ�g���G� }�r0WARNM�p�#tC�v`�ç` � C�OR-UrFLT�R��TRAT9 T|%p� $ACCVq���� ��r$OR�I�_&�RT��S\<��0CHG�0I�E��TW��A�I'��T��!D��� ��202�a1��HD)R�2��2�2J; ST���3��4��5��U6��7��8��9 1�׀
 �2 @.� TRQ�$vf��4'�1�<�_U<�G�z�Oec  <� �P�b�t�53>B_�LL�EC��!~�MULTI�4�"u�Q;2�CHILD��&s0wDET� "'�STY92	r��=���)2���ױ��ec# |r056$J ���`���uTOt���E^	EXTt�����2��22"(M����$`@D	��`&��X������ %�"��`%�ak�����s�����&'�E�A�u��Mw�9 �% ���TR�� ' L@U#9 ���=At�$JOB���мP�TRIG��( dp������^'�#j�~�x�pOR��) t$�FL��
RNG%Q@�TBAΰ �v&r�*`1t(@��0 �x!�0�+P�pX�%���*��͐�U��q�!�;2J�_)R��>�C<J�8*&<J D`5CF9��`�x"�@J��P_p��7p+ \@RO0"pF�0��IT�s�0NOM��>Ҹ4s�2��� @U<PPgў�P�8,|Pn��0�P�9�͗ RA���l�8?C�� �
$TͰt�MD3�0T��pU(�`�΀+AHlr>�T1�JE�1\�J����PQ��\Q��hQCYN�T�P��PDBGDd̰�0-���PU6$`$Po�|�u�AX�܆��TAI�sBU�F,����C�1. �����F�`PI|�U-@PvWMuXM�Y��@�VFvWSIMQ�STO�q$KEE�SPA��  ?B�B�>C�B?�P��/�`��MARG�u2��FACq�>�SLEW*1!0����
��17_MCW$0'����pJB�Ї�qDE�Cj�eN"s�V%w1 Ħ�CHNR�;MPs�$G_@�g�D�_�@s��1_FP�5�@TC�fFӓC@�Й���qC��+�VK��*��"*�JRx���SoEGFR$`IOh!v�0STN�LIN>��csPVZ��R�A�D2 ����r 2��hr�r�R~��3` +^? ���եq�`Kҥq|`������t��|aSIZ#�!� �T�_@%�I��qRS�*s��@2y{�Ip{�pTpLF�8�@�`��CRC����CCTѲ�Ipڈ�a���bL�MIN��a1�순���D<iC �C /���!uc���4�n j�SEVj���F��_!uF��N����|a��=h�?KNLA�C2��AVSCA�@AP��2�@�4�  �cSF�$�;�Ir ��C�a�05��	 D-Oo%g��,,m�����ޟ�URRC�6� n���sυ��U��R�0HANC���$LG��ɑDQ�$t�NDɖ��AR۰N��aqg��ѫ�X��ME��^�Y�[PS�RAg�X�AZ�П���:rEOB�FCT��A���`�2�!Sh`0ADI��O��y�"y�n!@�������~#C�G3��!��BMPmt@�Y8�3�afAES$���v��W_;�BAS#?XYZWPR��*��m!��	�QU�87/  ƀI@d��2�8\�p_C:T��n�#  ��_L
 .� 9 ���C�/�Y(zJ�LB�$��3�D��5�FOR�C�b�_AV;�M�OM*�q�SaԫBP�`Ր�y�HBP�ɀE�F�����AYLOAD&$ER�t&3�2��Xrp�!u�R_F}D�� : T`�I�Y3��E�&��Clt��MS�PU
a$(kpD��9 �rb�;�B�	EVId��
�!_IDX��$���B@X��X<&�SY5� ��0R_H�0e�<>��ALARM��2W��rMER��0=C hb Pnq�`M\q�J@$PL`A&�M#�$�`��� 8�	�P��V�]�0���U�P�M{�U��>�TI-Tu�
%�![q�Y�Z_;���? ��B pQk��6NO_HEADE^az��} ѯ��`􂳃���dF� ق�t� ���@�@|��uCIRTR�`$��ڈL��D�CB@4�RJ����[Q���cA�2>���OR�r���O����T`UN_OO�Ҁ$����T(�����I�VaC|q= � PXWOY���=B}p$SKADR�Y�DBT�TRL
��C��րfpbDs�L�~�DJj4 _�bDQ}��PL�q�wbWA���WcD��A��A=�2�U�MMY9��10��+����D;[QP�R�� 
��D8�Z���E O�Y1�$�a$8�9K�L)F!/�2����0GG/���PC�1Hf/���PE+NEA@Tf�I�/�#��RECOR`"J�H @ �E$L�#F$#PR��`�+jp��nq�_D$�qPROSS]�
����R�r�` u�$TRIyG96PAUS73>ltETURN72�+MR:�U 0Ł0�EW$��SIGNsALA�QR$LA�м�5�1G$PD�'H$Pİ�AI�0�Ab�C�4�C��DO��D�2�!�6GO_oAWAY2MOZq��Z�W DCS��CwSCBg�K Իa\#���ERI�0Nn�!T�`$�����FCBxPL�@QBGAGE�� �P��ED|BD�wA[CD�OF�q[F0�FoC��MPMAB0XoC�?$FRCIN��2Dxk��@��$NE�@��FDL8�� L� ����=��Rw��_��P� OVR1�0���lҠ�$E�SC_�`uDSB�IO����pTe�E�VIB�� `s��Z�8�V��pSSW��$�&VL��:�Lk��X����ѣ�bQ����US�C�P��A=�	Q��MP1%e&S*`�(bt`:'c5۳ESUd�� -cWg&SWg?cWd�����Wd��Wd.���AUT�O$�Ya҃�ac�SB ����-d��&SwB[���GB�f$VOLTr�g ��  � GAOD!�q���@:ЗORQҀKra�$DH_THE&0��Rgp� qtnwALPAHnt��o��w0 Vp]�$�.�Ra�[��s�5 �`r�CQ#BUD�S� %F1M��sV
���;��Lb�tk����BRTHR��L��T(`�Z��VɖL��DE  �1��2�⋅�������� kѯ�aәTt0V�ꆸ� �����̈Я�-�"��N~��sS2����IwNHB��ILTG0 ɡ�T?��3$�w��E���PqQxQ�TqPe��0Y�AF}�O�ນ�� ڗ��qPڳē��`��bPܙ���PL?�x��3���TMOU�� ēS���� ��s�/�S1H8���O�Aܙ��I�����CDIƑ˩o�S#TI��գ�O:ҋ�,0���AN��Qg`�S��+r�#x$�Ј���w�_����PR	A�P`vC����GMCNeQe�����VERS��r�oPIw�FPåǲШ۷-G.�DN��G>���B��F�2�Ƿ�Mʪ7�F��_�MN�D ̠,����d�{ƭa����OB���U˱z���DI���#���3� ����A���w�Fx���3�ON�5��Q��VAL�CR[�_�SIZ��b�;Qn�REQ�Rb��]2b���CHq�΂�ڃ��`������:�n�S_U���X��wWFLG����wU$CV�iM8GP�QδFLXP�92`3R�u���EAL�P�-�C	��+rT��W���� �R�c���NGDMS7� ��K>S��P_M'0h�STW`v������AL�P ���Q���U���U�IAG,�o��d�U�J-�T"A-`� �� �A�����H`��Q`��6��Pq_D&��1s ��.�P�F�>2�=T�� ?7 @1A>��#�#L��?_=i @@>�LD�c���0�FRI�0 `Ѐ��1}ѲIV\1�*�^1�UP`��a��C�LW��
`�L=S&-c&&S�C .w�� L���!����d�Q$w�҇��$w�����
�P�5R�SM���V0h b� r��d^2AW�a�_TRp}�8@NS_PEA����< ��$�SAVG�8�6G]%8���CAR �`0�!�$���"CRa����$ d�#E�@��"STD���!Fpo��'�QOF��%��"RC���&RC۠�(F��2A�R#7���%, gMEA�Q_�a��
QQ�(�al2��u4Ib�r7�I�R�9wQ�7�8M�/��!CpR�  ��p�2F<�SDNH�a   E
P2QM P $Mi� �s$cA�$C�cm�9����4�AT�0CY_ N LS!IG1x'yB��y@@H2Y�NO�����SDEVI�@ �O@$�RBT�:VSP�3�CuT�DB�Y|�A	W`3CHNwDGDAP H@�GRP�HE iXL��U��VS�Fx2� DL1p Q6ROp��sFB�\]�FEN�@���S��ChAR �d�@DOd�PMCSb�P薇P�R��HOTSWz42�D�MpELE�1/e�8C8`�RS T�@��`�r� hf��`OL�GCHA�Fk�Fs����C�A@T � �$MDLUb 2S@�E���q�6�q	0P�i�c�e�cJ��	u�ݢ�#~5t+w�PTO���� �b��DS�LAVS� U  ��INP �	V��t�yA_;�ENUAwV $R�PC_�q*�2 1bL�waD�p�SHO+� W  ���A�a�q�2�r�v��u�vS_CF� ?X` ,f��r�OG gE��%D�h���pC�Iߣi�M�A��D�x AY?�W�� p�NTV	�D�V�E�0@�SKI��T��`g?Ň2�� JZs�! Cꆻ��f��_SV� �`XCL�U��H���ONLd��'�Y�T��OT:e�HI_V,11 AP7PLY��HI4`;��U�_ML�� $VRFY8�	�U�=M{IOC_I���"J 1"��߃O�@X��LSw"`@$DUMMY4���ڑ�C=d L_TP���8kC��^1CNFf��@�E��@T�y� D_#�UQ_��ݥ�YPCP���=�� �������uJ �� Y �+�
0RT_;P��uNOCCb Z�r�TE���=�פrOdG�@[ D��P_BAe`Lkc�!��_���H��d��E �\�pAb=cAR�GI�!$���`[� B�SGNA]� ��`U��IGN��Տ��� ��V�������ANNUN���&�˳�EU�J'�ATCH��J��8pt�rA^ <@g������:c$Va��`�����QEF] }I�� _ @@�FͲITb�	$TOTi �C�O�c��u�M�@NI�a`(tB��c���A>����DAY@CLOAD��D\�n���� ��EF7�XI�Ra���K���O%��a:?�ADJ_R�!@Eb��>�H2�"[Ӑ
 c�%��`a͠MPI8�J��D �A��?�Ac 0��х�� $��Z�ϡ�Ui ���CTRL� Yp ;d��TRA8 ?3IDLE_PW  ЏѠ��Q��V�GV_���`c O`p�;Q@?e� 1$��6`<cTAC-3��P�LQH�Z�Rz\ A-u6:ɰSW;�A \���"J��`b�K�;OH�(OPP; �#�IRO� �"BRK��#AB �O��� ���� _ ���F���`�d͠, j@S�RQDMW��MS�P6X�'�z��IFECAL,�� 10^tN��V―�豊�V�(0}f�C)P
��N� Yb� !gFLA_#�OVL ��HE���"SUPCPO��ޑ\�L�pH��&2X�$Y-
Z-
W-
��/��0�GR�XZ�q�$Y2&�CO�PJ�SA�X2 R��*r�!��:��"�byI�0)�f `�@/CACHE��c؛�0�s0LAZ SU7FFI, C��q\���6o��1M�SW�g 8�K�EYIMAG#TM�@S��n
2j�r|�2��OCVIE���~�h �aBGL����`�?�@��@��j�i��!`STπ!�������x���EMAI�`�N��`A�@Z�FAUD� �j�"�qa��U�3G�u E}�?k< $I#�U�S�� �IT'�BU!F`��DNB���'SUBu$�DC_���8J"��"SAV�%�"�k������';��P��$�UORD��UP_pu �%��8OTT��1_B`��8@LMl�F4���C7AX@Cv���XXu 	��#_G��
 @'YN_���l6���UD�E��M����T��F� caC�D]I`BEDT)@C���~�m�rI�G�!c�&���l`���a�P��F�ZP n (�pSV� )d\�ρ��E��?o� �����>"$3C_R�IK ��kB��hD{pRfgE�.(ADSP~KBP�`�IIM�#�C�Aa��A��U�G���iCM! IP��KC��� �DCTH� �S�B*�T���CHS�3�CBSC��� ��V�dYVSP�#�[T_DrcCONV��Grc[T� �Fu F��ቐd�C�0j1��SqC5�e]CMER;d>AFBCMP;c@�ETBc p\FMU DUi ��+�~�CD�I%P702#@O���qWӏ�SQb��QǀSU��MSS�1ju�4`�T��Aa��}A�1r� "��<���4$ZO@s�D��l�U6�&��eP���eCNc�l��l�l�i�GROU�W)��S c�MN�kNu�eNu@�eNpR|b|�i�cH�ppi��z
 �0CYC����s�w�c��zDEfL�_D��RO�a@���qVf���v{�O� 2���1��t��:R�ua��.#�:���AL� �1sˢI1¡�J0��PB���AR^�T�Gbt ,!@��5h��aGI1LcR1s�0"�0R����1u����H�����P����Cڠ	���������J0��0vH *	�L U�1#J�Q��V
�[�7A z���z��z��z�Ѩz�Fz�7w�8w�9Pw���y���1��1��U1��1��1Ě1њU1ޚ1�2��2�����2��2��2��2�Ě2њ2ޚ2�3J��3��3����3��U3��3Ě3њ3ޚe3�4��I�XTF��1w6�.(�0�f�0�U�0ŷ�e>`FDR�5�xTU VE���?1���SR��REr�F���OVM~Cz)�A2�TROV2ɳDT� R�MXa�I�N2���Q�2�IND�p�r�
���0�0�0G@u1��[�G`��{�D_֎[�RIV�P��G�EAR~AIOr�K"N�0�y�p�5`�@�a�Z_MCM�� �����UR�Ryxǀ��!? ���p?nЋ�?n�ER�vт��!�P���zE@:�PXqB�R�I0%L�#ETUP?2_ { ���##TDPR�%TBp��p����I��"BAC�2G| T��"�4)�:�%	`^B��p�IFI��� Mc���.��PT���FLUI�} � ��K UR�c!���B�1SP�x E�EMP�p�2$���S^�?x��J8ق0
3VRT���0_x$SHO��Lq�6 ASScP=1��PӴBG_���������FOR�C:dh�d~)"F%UY�1�2\�2�1�Q�h� p� |��N�AV�a��������S!"��$VI�SI��#�SCM4S�E����:0E�V�O���$���M����$��I��@��FMR2��� �5`�r�@ �� �2�I�9 F�"��_���LIMI�T_1�dC_LM�������DGCLFl����DY�LD��B��5�������M��Fc��u	 T��FS0Ed� P�QC�0$EX_QhQ1i0�P�ajQ3�5��GoQ���� ����RSW�%ON�PX�EBU1G��'�GRBp�@mU�SBK)qO1L�7 ��POY 
)P��P��M��OXta`SM��E�"������`_E � ��0� �TERMrZ%�c%�ORI�1r_ �c%�0�SMep	O��_ ��&>`�`�(وc%�QUP>� ��� -���bQ���q#� ���G�*� ELTOQ�p�0�PFIrc�1Y��P|�$�$�$UFR�$��1L0e� OTY7�PT4q�k3wNST�pPAT�q=4PTHJ�a`�EG`*C�p1ART�� !5� y2$2REyL�:)ASHFTR(1�1�8_��R�PcJ�& � $�'@��  ��s�1 @I�0��U�R G�PAYLyO�@�qDYN_k����.b�1|��'PERV��RA��H��g7�p��2�J�E-�J�RC����ASYMFL3TR�1WJ*7�����E�ӱ1�I��aU�T�pbA�5�F�5P��PlC�Q1FOR�pMF�I!���W���/&�0F0�a  �9H��Ed� �m2N�,��5`OC1!?�$OP����c������bRE��PR.3�1a�F��3e��R�5e�X�1(�e$PWR��_����@R_�S�4��et$3�UD�ҸПQ72 ]���$H'�!�`�ADDR�fHL!GP�2�a�a�a:��R���U�� H��SSC ����e-��e���e���SEE��aSCD���� $���P_"�_ B!rP����}I�HTTP_���HU�� (�OB�J��b(�$�fL�Ex3Us�� �� ���ะ_��T�?#�rS�P��z�KRN�LgHIT܇5��P ���P�r������PL���PSS<�ҴJQUERY_FLA 1��qB_WEBSOC���HW�1U����`6PINCP	U���Oh��q�����d���d���� �I�HMI_ED� T� �RH�?$��FAV� d�Ł��wOLN
� 8��yR�@$SLiR�$INPUT_�($
`��P�� �؁SLA� ����5�1��C���BMIO6pF_AuS7��$L%�}w%�A��\b.1��0���T@HYķ��SCHg�UOP4� `y�ґ�f�� ��������`PCC
`�����#���aIP�_ME�񵁗 X�y�IP�`�U�_N#ET�9���Rĳ8s�)��DSP(�Op�=��BG��Я�M��A��� lp:CTiAjB�pAF TI�`-U��Y ޥ�0PSݦBUY IDI�rF ���P��!�� �y0��,����Ҥ�N�Q�Y R��IRCA|�i� � ěym0�CY�`EA������񘼀�CC����R�0�A�7QDAY_<���NTVA�����$��5 ���SCAd@��CL����e���𵁛8�Y��2e�o�N_�PCP�q������,�N����
�xr࿀�:p�N� 2!��Ы�(ᵁ����xr۠LABy1��Y .��UNIR��Ë �ITY듭��e�R�#�5���R_U{RL���$AL0 �EN��ҭ� ;�T��T_U��ABKsY_z��2DISԐ��AH�Jg�����P�$���E��g�R���З A�/���J����FLs��7 Ȁ|���
�UJR� ��pF{0G��E7��J7 O^ R$J8I�7�H�R�d�7��E�8{��H�APHIQ�S��DeJ7J8�B��L_KE*� � �K��LM�[� � <X�X�Rl�u���WATCH_VA��o@D�tvOFIELc��cy� L��4� � o1Vx@��-�CT[�9�m�<���LGH���� $��LG_SIZ�t�z�2y�p�y�FD��Ix���+!�� w�\ ����v��S��� 2��p�������\ ��h�A�0_gCM]3NzU
RFQ\v�v�d(u�"B ��2�p����I��+ �\ ��jv�Rː_�0  ��ZIPDUƣE�L)N=��ސ�p��z6���f�>sD�PL�MCDAUiEA`Fp���TuGH�R���|�BOO�a��� C��I�IT0+���`��RE����SCR� �s��DIr��SF0�`RGIO"$D�����T("�t|�S�s{�W$|�XJGM^'MNC�H;�|�FN��a&K�'uЅ)UF�(1@�(�FWD�(HL�)STP�*V�(%Г(��(RS9HIP�+��C[T�# R��&p:'^9U=q�$9'�H%C�2�"Gw)�0PO�7�*���#W}$���)EX.��TUI�%I���� ����rCO#C� *�'$S��	)���B@�NOFANA|��Q
�AI|�t:��EDCS��c�C�c*�BO�HO�GS���Br�HS�H(IGN������!O���DDEmV<7LL��H��-��Ц(�;�T��$��2�p�����(1R�Q�ѧ(�`뀸{�Y��POS1�U2��U3�Q��2�@�Ш# ��{�PtD�� ��&q)��0�d��V+STӐR�Yl�\@~ ` �$E.fC.k�p<p=fPfX��3�ѩ LRТ� �� x�c�p��<�Fp�did^�_ ������Kq&���c��MC�7� ��pCL�DPӐ��TRQLaI#ѽ�ytFL��,r�5s8�D�5wS��LD5ut5uORG���91HrCRESE�RV���t���t�� ��c�� � 	`u95t5u��PTp���	xq�t�vRCLMC������D�q>�M��k�������$DEBUGMCAS��ް��?U8$�T@��Ee�g���M�FRQՔ� �� j�HRS_R%U7��a��A��k5�FREQ� �$</@x�OVER���n��V#�P�!EFI�%�a��g��t����t� \R�ԁd�s$U�P��?A���PS�P��	߃C ��͢a��U\�l��?( 	oQMI;SC� d@�QkRQ��	��TB �� Ȗ0A՘AX����ؗ�EXCE�Sj��M��\��§������a��SC>�P � H��̔�_��Ƙǰ]���C�MKHԳK�J� �m�B_K�FLIC��dB�QUIREG3MO��O˫3��quL�`MGմ �`���T��R�NDU�]��>��k��G�Df��INAU9T���RSM>�a��@N)b]3-���5��PSTL\�� 4nX�LOC�VRI%�v�UEXɶANGuB�u��?� A��ŷ�������MF O����Y�b@�e4Ŝ2k�SUP�f�pF�X��IGG� � �A��c���c Q6�dD�%�b|�!`�Ȁ!`��|��3w�ZWa�T!I�V�� M��[��� t��MD��I��)֟@���H8ݰM��DIA��ӂ��W,!�wQ�1�D��)?�O���]��[ 0�CU��VP�(�pu���O!_V���� ���S�X�5������P��0N���P��KES2����-$B� ����ND�2����2_TX�dXTRA�C?�/���M�|q�`�P�v��XҰ�Pt SB�q`�USWCS��Tx��	���PULS��A�NSޔ��R��JOIN��H��~`j�=��b��b�����P=��$��b$���TA����S���S�H�S�E��SCF���J��R��PLQ��a�LO��н.���� ��8��������0�RR2���� 1��eA�q Kd$��Iΐ+�G�A�2+/� ΍PRIN�<$R SW0"�a/�wABC�D_J%�¡��_J3�
��1SPܠe��P���3��р`�B�J/���r�qO8QyIF��CSKP"z�{�{�J���Q�L2LBҰ_A1Z�r�~ELQ��OCMPೕ�T����RT�����1�+���P1��>@�Z�SMG0��=�;JG�`SCL�͵OSPH_�@��%�V�� RTER0`  �< A_�@G1�"�A�@c��\$D�I�
"23UDgF  ǀ~ LW�(7VELqIN�b)@� _BL�@u��$G �q�$�'�'�%`<�� �ECHZR/�TSAY_`� ���E}`B<����5�B��1:}`_�� �)5D2d%�PA4I��N9t&i`�DH�A���ÀP�$V `�#>A$���ł�$Q�R}ӆ��H �$BELvᵆ<!_ACCE�!c��7</��0IRC_] ���pNTT��S$PS�rL� d�/E s��F{�@F
��9�gGCgG36B���_��Q�2�@�A���1_MGăDD�A]"łFW�`���3�EC�2��HDE�KPPAByN>G��SPEE�B �Q%_pB�QY�Y��1>1$USE_��,`]Pk�CTReTYP��0�q P�YN��A e�V)хQM����ķ��@O� YA�TINCo�ڱ�B�DՒ�WG֑ENC����u�.Ax�2Ӕ+@INPOQ�aI6Be��$NT�#>�%NT23_�"ł�IcLO� ł_`��I �œif� œk�? �`� ej�C400fMOS�I�A���ОA䃔�P?ERCH  �c��B" �g��c��lb=������oUu@�@	A6B(uLeT	~�1epT�ljgv�fTRK@%�AY��"sY��q6B��u�s۰�]��RU�McOMq�ՒY�MP�Ĕ�C�s�CJR���DUF �BS_BC?KLSH_C6B)� ���f���St�H��RR�|�QDCLALM-dp���pm0��CHK|���GLRTY����d��Y��)Üd_UM]�ԉC��A!��=PLMT� _L �0��9��E�.�  ��#E)�#H� =��Q�3po�xPC�axHpW�頿EׅCMCE�\�@�GCN_,ND�LΖ�SF�1�iVoR���g<!��6B���CATގSH)�,�D fY��f��7A���f܀PAބ�R_P݅�s_ �v���s,����JG�T]����Y�����TORQU`aP��c�yPOU��0�b��P%�_W�u�t���1D��3C��3C�I*K�IY�I�3F�6������@VC�00RQ�t��1���@ӿ��ȳJRK�����Up�DB M��UpMC� DL�1BrGRV�J�Cĭ3Cĳ3$�H_p��"�j@q�COS~��~�LN���µ�� �0�����u����̓�b�Z���f$�MY���؊���>�THE{T0reNK23�3�hҧ3��CBm�CB�3C! AS� ��u�0�ѭ3��m�SB�3��Nx�GTS$=QC������������$DU��Kw�B�%(�
�%Qq_��a��x�{�K���b(��\�A�`Չ��p�{�{�LP!H~�g�Aeg�Sµ�� ������g������֊��V��V��0��V���V��V��V��V*	�V�V%�H��������G�����H��H���H	�H�H%�OJ��O��OV	��O��UO��O��O��O	�O�O�Fg���	������SPBAL�ANCE_-�LmE��H_`�SP!1��A��A��PFULCElTl��.:{1��UTO_�����T1T2��22N���29`�!anPL�=B�3�qTXpOv |
A4�INSEG�2��aREV��`aD3IF�uS91�8't"1�`OB.!t�M���w2�9`��,�LC�HWARRCBAB�� ��#�`-ФQ 5
�X�qPR��&��2�� 
�""��1e7ROB͠CR6B5��� ��C�1_���T � x $WEIGH�PFrp$��?3àI�Q�g`IFYQ�@LAGĒRq�S�R �RBI�Lx5OD�p�`V2S	T�0V2P!t�W0�1(1�&1/0�30
�P�2<�QA  2řd[6/DEBUg3L_@�2=�MMY9&E qNz�Drp$D_A��a$�0��O�  �DO_@A.1� <B0�6�Hm�Q�B�2�0N-cRdH_p`�P��2O�� �� %��T`"a��T/!�4)@�TICKh3| T1"1@%�C ��@N͠�XC͠R?��Q�"�E�"|�E8@PROMP�S�E~� $IR���Q��R;pZRMA�I)��Q�R4U_r0�2S; �q�PR8�C�OD�3FU�Pd6I�D_[�vU R!G�_SUFFu� �l3�Q;Q�BDO`�G �E�0�FGRr3 �"�T�C�T�"�U�"�UPׁ�T8D�0�B0Hb �_FI�19*cO�RD�1 50�23�6V�+b�Q1@$Z�DT}U���1;E��4 *:!L_NA�mA�@�b�EDEF_I�h�b�F�d�E�2�F��4�F�c�E�e�FIS�P��PAKp�Ds�C��d��44בi��2DP�"�It�3D�O#>OBLOCKEz��S��O�O�Gq�R�PUM �U�b�T�c�T�e�T!r �R�s�U�c�T�d�R�6 �q�S� ���U�b�U@�c�S�Z��X�@P`  t�@qe�)@W�x��:�ss0�TE�<D��( l1LO�MB_��ɇ0V2V�IS;�ITYV2A���O�3A_FRI��a SIq�Q!R�@��@�3�3V2�W��W�4����_e��QEAS^3�Rϡ���_�[p:R�4�5��6_3ORMUL�A_Iz���TH]R^2 �Gtg�30�f��<8�5COEFF_O�A	 ��A���GR�^3Sg0BCAnO/C$��]3���0�GRP� � �G $�p�YBX�@TM~w���u�B�s��bCER, Tttsd$`7�  �LL�TSpS~�_SVNt�ߐĸ�$`���$`� ���SETUsMEA*P�P��W0�1+b>/0� � h��  @ڐo�l�o�cqDz��b�@cqq`t�P�G��R�� Q\p�*q[p��>�c NPR�EC>at��ASKy_$|�� PB1?1_USER�����{ ���VEL@���{ 0�$Ō!I]`���MT�ACFG>���  �@@ =O�"NORE-0l@,o�V�SI.1�d��6��"UXK�fP!��D�E�� $KE�Y_�3�$J3OG��0SV���0���!��}�SW�"�ah\aS�ՐT|�GI��5@| ^�� 4 �h��'d2�!XYZ�c���31�_ERR#�� 8Ԡ�A�fPV�d��1�����$BUF��X����_�MOR|�� HB0CUd�lA�!���GQ\aB�,"!a	$� ���a�����?�G~�� � �$SIՐ���VOx��T�0OBJE_���ADJU)B��EGLAY���%�DR�OU.`=ղВQ0b=��T���0���;BDIR���; I�"0DYNW�#���	T��"R���@�0�"�OPWORK����,%@SYSB9Uy�SOP��$ޑ�U�; P�pN�<�PA�t�>�"��+OP�PUd!0�`!z��l�IMAGw�1B0y�2IM�Õ��INe�d��RGO�VRD��-��o�P q��0��J�Os���"�L�pBa���o�PMGC_Ee`���1Ny M A�21�2U����SL_��� � ?$OVSL�ǫň?q�`��2�" -�_ ��k�P��k�Pu���2�C� �`�Ź����_ZER�D��$G�� 1�>���� @*���%MOh`RI��� 
�JP8+�=!/�L���ح�T� �0AT�US��TRC_T���sB��}fs��9s�1Re`��� DFAm����L���"��00a� ޱ��XEw{�����C0vcUP��+p	qPXPȝj�43 � ��PG\���$S�UBe�%�qe9J?MPWAIT z�}%LO��F�A�R�CVFBQ�@x"�!R��� �x"ACC� R�&�B�'IGNR_{PL9DBTB�0Pqy!BWbP�$w��Uy@�%IGT�PI���TNLN�&2R���rL�NP��PE�ED \HADO!W�06�w��E[q4�jO!�`SPDV!� LbAz�`�07��3UNIr��0"!R��LYZ`� o}��PH_PK���e�RETRIE�9{�q����0'PFI"�� �G`�0D� 2�g�DBG�LV�#LOGSIYZ��EqKT�!U��2VDD�#$0_T�G��MՐCݱ��|@eMR�vC}�3�CHECK�0���PO�V!�2k�I��LE(!���PArpT�2K�W���@P2V!� h $ARIBiR� c��a/�O�P8�ӐATT��2�IF|@z�Aq�4S�3UX����2L9I2V!� $g���OITCHx"[�W �;AS9N2N xR�LLBV!�� /$BA�DYs���BAM!���Y9F�PJ5��Q��R6�V>�Q_KNOW�Cb��U��AD�XV��0�D�+iPAYLOAt��Ic_��Rg��RgZOcL�q��PL�CL_�� !@7��b�QB��d���fF�iC֠�js��d��I�hRؠ�g�ҢdBd����J��q_J�a:���AND��Ĳ`.t�b�a�q�PL0?AL_ �P�0P���QրC��DNc�E���J3CpWv�{ TPPDCK�������P�_ALPHgs�sBE��gy|��K�1�� �s ���HoD_1Oj52ydDP�AR�*���;�&���TIA4�U�5U�6��MOM���a���n���{�Y�B� ADa���n���{�PUB��R��҅n��҅{�A2�Wp��W �/  PMsbT�� BxQ���?� e$PI��81���TgJ��niJ�I
V�Id�Ir��[��3!��>!��r�Ӫ�U3HIG�SU3�% �4얎4�%� ���"�����!
��!�%SAMP���^��_��%�P4s ю���[  	ӝ�3 ���0���&��������^��Sp��H&0	�IN�SpB��� �뤕"��6��6�V�/GAMM�SyI�F� ETْ��;�D�tvA�
$ZpIBR!�62IT�$HIِ_������˶E��ظAҾ���LWͽ�
̀��7���rЖ,0�qC��%CHK��" �~I_A����� Rr�Rqܥ�Ǚ��ԥ�|��Ws �$�x� 1���I7R�CH_D�!� R1N{��#�LE��ǒ�!,��x���90MS�WFL�$�SCR�((100��R@��3 ]B��ç��a����َ0ޤ�PI3A9�ME�THO����%��AXH�XX0԰62�ERI��^�3��R$�0$u	��pF{�_����?ⲣ1�L�L8�_�a�OOP����8wᲡ��APP:���F���@{���أR	T�V�OBp�0T���0�;��� 1�I���� ��r���RA�@MeGA1�ЫSSV-�w�P_@CURg��;�GRO[0S_�SA�Q��Y�#NO�pC!"�tY�� Zolox�������!b��,��&�DO�1A���A ����Х��A���A"�0WS�c �qwP}M)�� � �ãYLH�qܧ��S rZ�]B�o��0��Ĕ�q_�C1��M_W���g���c�M� �`Vq�$Ap�x1o�3"�PMJ�,�� �'A� 9�!YWi:�$�LWQ |ai�tg�tg�tg{t� �N`���S��JSpX�0O�sRqZ���P� *�� ���M��������������@X��� ��@!��q_~R� |�q#(Y����& n��&{�Y�Z��'�&t�|�Q�� ���%J0��@}`�$PQ��PMON_QU�c� � 8�@Q�COU��%PQTH��HO�^0HYSf:PES�R^0UEI0tO��@O|T�  �0�PGõz�RUN_+TO��POْ.�'� PE`�5C��A�<�INDE�ROGGRAnP� 2g��NE_NO�4�5I�T��0�0INFO�1� �Q�:A��ȇOIB� (��SLEQݖFAѕ�F@�6 0OSy�T�� 4�@ENAB|��0PTION.S%0ERVE���G���uPzCGCF�A� �@R0J$Rq�2�
��R�H�O�G�"��EDIT�1� ��v�K�ޓʱE��NU0W*XAUT<u�-UCOPY�ِ(N\����MѱNXP\[^q�PRUT9� _R�N�@OUC�$�G�2�T �$�$CL`?0���0��� �  ��P�S�@�X��PXK�QIRT�U��_�PA� _W�RK 2 e��@ 0  �#5�QMoYhJo|m |l	�`�m�o�� `��o�o�f�e �l}�aI[ct�'`BS�*� 1��Y� < 7������� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t�`��������srCC��gLMT?0���s7  dѴINڿ��дPRE_EXE��)�Ƅ0jP��z�a'`DV��S�@�e)�%sel�ect_macr�o����kϤ�qtIOgCNVVB�� ��P��USňw���0�V 14kP $�$p��a�|�`?��Ɛ >�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o (:L^p��� ���� ��$�Ѱ�LARMRECOV ^�����LMDG ��Ь�LM_IF� ��d  �YST-040 �Operatio�n mode A�UTO S��ed� eed lim�it.(L:6) ������)�;�M�_��q��, 
 ����#�>TELE�OP ǘLINE� 0ǑقABOR�TEDǘJOINTǐ8 %�����C$���1��ᕜA��ATAǒؑ3���גؒ��  clear䀪���ί���NGTOL  ~@� 	 A |����ѰPPINFoO �� f��L�^�p����   ������k���ۿſ�� ���5��Y�C�iϏ�%���ٯ�������� ��'�9�K�]�o߁���ߙ�PPLICATION ?t������Handlin�gToolǖ �
V9.40P/�17���
8813ǀ����F0�	�549���������7DF5�О�ǓN�one��FR=A�� 69��_ACTIVE1�s  �� �  ��.ڀMOD���������CHGAPON�L�� �OUP�L[�1	��� �>�B�T�f���CUR�EQ 1
��  UTp�p�p�	�� ������l��������������i3l�;p���^�H��A�t
HTTHKY�FXv |��*<N `������� �//&/8/J/\/�/ �/�/�/�/�/�/�/�/ ?"?4?F?X?�?|?�? �?�?�?�?�?�?OO 0OBOTO�OxO�O�O�O �O�O�O�O__,_>_ P_�_t_�_�_�_�_�_ �_�_oo(o:oLo�o po�o�o�o�o�o�o�o  $6H�l~ ��������  �2�D���h�z����� ��ԏ���
��.� @���d�v���������Ƃ�TO�����DO?_CLEAN���E�NM  �� p�������ɯۯ�v�DSPDRYRLL���HI��o�@�� G�Y�k�}�������ſ�׿����ϻ�MA�X��,�呿��=�X�,�<�9�<���PLU�GG,�-�9���PRUC��Bm�q�6��(ϗ�O����SEGF�K���� �m� �G�Y�k�}ߏ�����LAP$�7ޡ���� ��+�=�O�a�s������ �TOTA�L_ƈ� �USENU$�1� �������RGDISPM+MC�d�C�O��@@�1�O"�D���-�_STRIN�G 1��
��M��S��
~��_ITEM1��  n���������  $6HZl~ ��������I/O SI�GNAL��T�ryout Mo{de��InpN�Simulate�d��Out`�OVERR!� �= 100��I?n cyclT���Prog Ab�orj��JSt�atus��	Heartbeat���MH Faul<��Aler�! /!/3/E/W/i/{/�/�/�/ (���(� ���/??&?8?J?\? n?�?�?�?�?�?�?�?��?O"O4OFO�/WORИ�~A�/XO�O�O �O�O�O __$_6_H_ Z_l_~_�_�_�_�_�_�_�^PO���"` �KoEoWoio{o�o�o �o�o�o�o�o/�ASew��bDEV%n�p9o��� �#�5�G�Y�k�}��� ����ŏ׏�����|1�C�PALT�- j��OD�������ȟڟ ����"�4�F�X�j��|�������į֯X�GRIB�������6� H�Z�l�~�������ƿ ؿ���� �2�D�V�h�z�����R�-��&� ���������"�4�F� X�j�|ߎߠ߲�������������PREGn�W���0�~��� ����������� �2� D�V�h�z���������~$�$ARG_~@�D ?	����� � 	$$	[]�$:	���SBN_CONF�IG�XW�qRCII_SAVE  $zm���TCELLSE�TUP 
%�  OME_IO�$$%MOV_qH� ��REP���#��UTOBAC�K� 	t�FRA:\D� �.D�z '`��D�w� �s � 25/1�1/29 20:_26:16D�;�D���#//h�� C/j/|/�/�/�/�/D��X/�/??(?:?L? �/p?�?�?�?�?�?�? g? OO$O6OHOZO�? ~O�O�O�O�O�O�O��ׁ  c_F_\�ATBCKCTL.TM�)_;_M___\q_8INIm���j~CMESSA�G� �Qz �[ODGE_D� �j�X�O�p�_@PAUS�6` !� , 	�; :oHg,		2oloVo �ozo�o�o�o�o�o�o  
D.Pz}d`?TSK  mw<}_CUPDT�P�W�d�p�VXWZD�_ENB�Tf
�vS�TA�U�u��XI}SX UNT 2�v�wy � 	�p	�C���� ��x��>�?����gD�R�W  C��#��'���4��&m�����R�����k`��;� B�' ����問��y����.�1�ME�T��2@��y P�Q�A�IAIz��A���A҅��A�h=B5�s�u�>��>i�Hy>yK�?
�0]?��?	��95�SCRDC�FG 1�Y ��  ����%�7�I�pD�Q��ݟ������Я ���[���<�N�`��r�������7���FG�R9��p�_ԳPNA�� 	FѶ_�ED�P1��� �
 �%-PEDT-¿ R�v����E�<�GE�D��;9/�>���  ����2�����B�  ����{�����j�����3��#� �G�Y���@G�ߠ�6�����4�W������Zݨ�� Z�l������5K��� ���Y�t���&�8���\���6��d��Yހ@����(��7 �S0wY�w��f���8����{�IZ��C/��2/����9{/��//L Zݤ/?V/h/�/�/��CR���?�?Tn?��? ?2?�?V?԰!�N�O_DEL�ҲGE_UNUSE޿�дIGALLOW� 1�   �(*SYST�EM*
�	$S?ERV_GR[�@n`REG�E$�C
��@NUM�J�C�M�PMU?@
��LAYK�
��PMPAL�PUCOYC10 N3^P<!^YSULSU_�M�5Ra�CLo_�TB�OXORI�ECU�R_�P�MPMC�NVV�P10|I^�PT4DLI�p��_�I	*PROG�RA�DPG_cMI!^Ko]`AL+e�joTe]`B�o�N�$FLUI_RE�SU9W�o�O�o�dMR�N�@�<�?�; M_q����� ����%�7�I�[� m��������Ǐُ돀���!�3�E�W�2BL�AL_OUT ��K���WD_A�BOR:PcO��IT�R_RTN  ��$�빸�NONS�TO�� lHC�CFS_UTIL� �̷CC_�AUXAXIS ;3$� h}�j��|�����ƽCE_R�IA_I`@��נ��FCFGG $�/�#��o_LIM�B2+�w �� � 	��SB\���$� 
Ԡ���)�Z���/�����[�����.R��H�!�����L��(
5������PA�`GP7 1H������A�S�e�w�6�CCV� C7��J��]���p������� CU������������U���é�̩�ձ�Uߩ�������ę;���PCk������������������R��ɱ���������� D� DU!�!�!�!�� ��&?��HE@ONFIpCѷG_P�P1H� +EH��ߟ߱�����������C�KPA�US�Q1H�ף IR�S�H�A��e� ������������� �E�+�i�{�a����A?Iץ�MؐN�FO 1��� �3��$4��A��PA�w��ǼiA�'.��gEB<���* D<Ş�B�Q_DF�C�@���B�I�Pb�O�� � ��LL/ECT_�!�����EN+`�ʒ��n�NDE�#��/�1234?567890�" �A��/ҵHw��#)j��<i{��; ��/��/`/+/ =/O/�/s/�/�/�/�/ �/�/8???'?�?K? ]?o?�?�?�?�?O�?t��$� �>�IO &��"S▒O�O�O�O`G[TR�2'DM(��0^�?�NN�(oM Z���_MOR)q3)H��7ىU3��Y�_ �_�_�_�_�[bR�kQ�*H�,S�?<�<ѠD<cz�KFd���P	,��;ϒo�o�o@˿�o�oœh�UY�@E�oS ��sja�PDB�.���4cpmidbg3��Рs:��>uqpz��v_  ��>x��}.��}�`��|�<�mgP���t���~f������@ud1:�?��Xq?DEF -��zC�)*�cO�buf.txtJ��|K�[`��/DM��>����R�A��MCiR2�0_{RCd���hS2�1����G���Cz�A�d4�EI�jA���	C-]�G�/X"B�e;F�]�H�j�C�1�aF�%J���iE&�mI�؂�LڒY�F��I�!o�N��mH�?aGMSo�������6f23DLD�	>�z�!� 2��}���yc
�@x9� C}�Ĵ  D4G��E���  E�%q�F�� E�p�u�F�P� E��fF�3H ��G�M��Ъ5�>�33���?�xn9�q@��Q5����RpA�?a��=L��<#�QU�@,�Cϒ����RSMOFST� +i�����P_�T1Ɠ4DMA �=ք�MODE 5dm�@��	Q�M�;��%��?����<�M>�{�Ͷ�TESTc�)2i�`�R�6�OߊK�CN�AB���n� �8��\�n�CdB͖��Cpp������p:d�QS ��� ������4ѕI7>���>B8rm5$�RT_c�PROG %j�%��d�1�h@NUS�ER��x�KEY_?TBL  e������	
��� !"#$%&�'()*+,-.�/(:;<=>?�@ABCc�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������>��͓���������������������������������耇�������������������s��4A8�LCK��xF�y��STAT��z2�X�_ALM������_AUTO_�DO�E�FD�R 3:i�2h�&q[~�� �BUOSYST-�322 Auto� status �check time out ����i�$TEL�EO8�i� ���)qA�ʜ@�Ĭ�����?��ڛMsB��õ�?*?���?Mf=��o�TR���-���D.��B���C��ϾB�N�*p��4�N4�J5H�j5H��>�i�B�J�d�BF��pZ��[~�bbt�����5/�M*F�B��GA+$����@R��J�}BQ�H�����������2>��@�@���&��CBxHCKH<B��6> Tbt��/��u�AUS�H?Z?l?i�$7? �?:�� mϸ?�?p�� �?�?OO�?,OfOxO �M6?�O�O�O~?�O	_ �?*_$_BOD_6_p_~_ T_�_�_�_�_�Oo)o ;o�OLoqo_�o�o�_ �o�o�o�o�o�oF Xo��No�� �o����@�N� $�b�x�����n��� ���A��b�\�z� |�n�������ʟ��� (�֏O�a�s������ T�ʯį��֯�� ��2�H�~���>���ɿ ۿ���ϼ�2�,�J� L�>�xφ�\Ϛϰ��� �Ϧ��1�C��T�y� $Ϛߔ߲ϴߦ����� ����N�`�߇�� ��V߼�������� ��H�V�,�j����� ��v�����$I ��jd���v�� ���0��Wi {&��\��� ��/&/�:/P/�/ �/F�/�/�/��/? �:?4?R/T?F?�?�? d?�?�?�? O�/'O9O KO�/\O�O,?�O�O�? �O�O�O�O�O
_ _V_ h_O�_�_�_^O�_�_ �O
oo"_$ooPo^o 4oro�o�o�o~_�o	 �_,Q�_rl�o �~�����&� 8��o_�q���.���� dڏԏ��� �.� �B�X�����N�ǟٟ 럖���!�̏B�<�Z� \�N�����l������� ���/�A�S���d��� 4�����¯Ŀ����� Կ�(�^�p���ϩ� ��f����Ϝ���*� ,��X�f�<�zߐ��� �߆����#���4�Y� �z�t�ߔ������ ������.�@���g�y� ��6����l������� ����(6J`� �V������) ��JDbdV�� t���/�7/I/ [/l/�/<�/�/� �/�/�/?�/?0?f? x?&/�?�?�?n/�?�? �/OO2?4O&O`OnO DO�O�O�O�O�?__ +_�?<_a_O�_|_�O �_�_�_�_�_�_ o6o Ho�Ooo�o�o>_�o�o t_�o�oo�o0> Rh��^o�� ��o�1��oR�L�j l�^�����|���Џ� ��?�Q�c��t��� D�����ҏԟƟ �� �"�8�n���.����� ˯v�ܯ���"��:� <�.�h�v�L�����ֿ 迖��!�3�ޯD�i� ��τϢ��ϖ����� �����>�P���w߉� ��FϬ���|�����
� ���8�F��Z�p�� ��f���������9� ��Z�T�r�t�f����� ������ ��GY k�|�L����� ���*@v �6���~�	/ �*/$/BD/6/p/~/ T/�/�/�/�/�?)? ;?�L?q?/�?�?�/ �?�?�?�?�?�?OFO XO?O�O�ON?�O�O �?�O�OO__@_N_ $_b_x_�_�_nO�_�_ o�OoAo�Obo\oz_ |ono�o�o�o�o�o (�_Oaso�� To���o���� �2�H�~���>��ɏ ۏ����2�,�J� L�>�x���\������ �����1�C��T�y� $������������� į��N�`������ ��V���ῌ����� ��H�V�,�jπ϶� ��v����߾�$�I� ��j�d߂τ�v߰߾� �������0���W�i� {�&ߌ��\������� �����&���:�P��� ��F���������� ��:4R�TF�� d��� ��'9 K��\�,��� �����
/ /V/ h/�/�/�/^�/�/ �
??"/$??P?^? 4?r?�?�?�?~/�?	O O�/,OQO�/rOlO�? �O~O�O�O�O�O�O&_ 8_�?__q_�_.O�_�_ dO�_�_�O�_�_ o.o�oBoXo�otc�$C�R_FDR_CF�G ;re��Q
UD1�:�W�P�aJ�d  ��`�\�bHIST� 3<rf  �`�  ?�R�@tAtB�b�C�P1pDtE�tItg�Ppo�tw�_��bIND�T_EN6p�T��q�bT1_DO  �U̫u�sT2��wVAoR 2=�gp� hq  7��R��|4�|�m[��RZ��`STOP��rT�RL_DELET�Np�t ��_SCREEN re~�rkcsc�r�Uw�MMENU �1>��  <�\%�_��T�� R��S/�U���e�w�ğ ������џ�	�B�� +�x�O�a��������� ��ͯ߯,���b�9� K�q�������࿷�ɿ ����%�^�5�Gϔ� k�}��ϡϳ������ ��H��1�~�U�gߍ� �ߝ߯�������2�	� �A�z�Q�c���� �������.���d� ;�M���q�������������YӃ_MAN�UAL{��rZCDƳa?�y�rG +���R�f"
�^"
?|(��PdT�GRP 2@�y��B� � s���� �$DBCO�pRIG���v��G_ERRLOG' A��Q�I�[m �NUM�LIM�s��u
��PXWORK 1B�8����//�}DBTB_�� C%����S"� �aDB_A�WAY��QGC;P �r=�ןm"G_AL�F�_��Yz����p�vk  �1D� , 
���/"�/%?/(_Mؘpqw,@�=5ON�TIM����t��_6�)
�0�'MOTNENFpF�;�RECORD 2�J� �-?�SG�O��1�?"x"!O 3OEOWO�8_O�O�?�O O�O�O�O�O�O(_�O L_�Op_�_�_�_A_�_ 9_�_]_o$o6oHo�_ lo�_�o�_�o�o�o�o Yo}o2�oVhz ��o��C�
� �.��R��K���� ����Џ?��ߏ�*� ����+�b�t�㏘��� ��Ο=�O�����:� %���p�ߟ񟦯��O� ǯ�]������H�Z� ��������#�5�����ϩ�i"TOLEoRENCv$Bȿ"� L��� CSS�_CCSCB 2%K�\0"?" {ϰϟ���7��
�� ��@�R�d�3߈ߚ�"�x���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg0y��� ���d���R�LL]��La�m1T#2 7C�C��F\�^ A�C�pC�ɴ�#�0� 	� A���B<���?�  �$�0���\0袰�0��B��`#s�K/]/(o/�ϓ/�/�/�s/�/�/�J��a�L~�?�I��:$z�:�5{OȦ��/��/T`?;�@��O? �?�?�?Ȏ0AF��?{F�A OO�7�1 ���9M	AB
AZO dBAE�9$O�O�O�Oi:�P��`�@0�DzJCA� @���
X-.
[#_   M?�>O�ڴ࿀q_�_�_�_:W�A< o:[<ǲ/o�/�_+oPoboto�eASCHC�V�WB$�Dz�cD�`�a=/�o@�oo�oW�a.+!⠲2=t,yD���Yr9��I?�-t �s�js�w�yj��������Q��� �@`��$�����A�� ��Bމ�o��'�9� �_]�o�N���r���ɟ ۟_�B�ʄ��YZ�>`� 9Bk��B�W@���?H�(�RE���Z�l�~���� `_м¯���
��� ̯9�,�]�o��� �H� ����ٿ뿊��ƿ3� E�W�iϬ���$ϱ��� �� Ϟ����/�A�S� ��w�V�h߭ߌ��S���ߐ�_�f	�� H�?�Q�~�u���� ���������D�� -�g�q����������� ��
@7Ic�m��߾�   �����)M@ qdv����� ��//I/P�m/� v/�/�/�/�/�/�/�/ ?3?*?<?i?`?r?�? ^/�?�?�?�?�?O/O &O8OJO\O�O�O�O�O�O�O�O�g	 � Q�P�s� �PC4p*�p�p6U6P\Cu9p/p�� ]VT^PM]�6P�:P�>P��VJ_�^P�bP�0fP�Vr]v��Tp Q�
k���_oo�id1Q&oNo ;o_cox�oˏUUA   �o<�k1Q@�  �o�kt�b����逡Up �� 1��6��1C���C�cPfL��?#�c>�{����`�cP�@@��d��r�`B�cP>�s�qC��p�����b�t<�o?��PH�)S�B���tq�q�p�r�`B���eIC�&�Q�4(� �oz�UU5�@�=�@9�^=��A��ϹRF9Q�-R��q�aA����tV@B��=�by��`ځ`  ?�p����U�[?����}t��$���$DC�SS_CLLB2� 2M���p�P�^?�NSTC�Y 2N��?�  ��� ����ʟ؟���� � 2�D�Z�h�z��������¯ԯ��SA�DEV�ICE 2O��!�$��4&V�h��� ����˿¿Կ���
� 7�.�[�R�ϑϣϵ������4(A�HNDG�D P��*�Cz|�A�LS 2Q��_�Q�c�u߇ߙ߫������?�PARAM RP��1�`�&տRBT 2T��/ 8�P<C�'pG �qi�l��sF@"�R��(qI�X���0�pB CW  ��B\x�N��Z��&���%��)���X�@j��p����zq�����B �(s,�F�p��V��q���b��B ��4&c �S�e�l�4+�����H1~�����D�C�$Z|��b���A,� �4�u@�X@��^@w���]�B���B�cP%���C4�C3�:^C4��n��� ��p8�-B�{B��A����� l��C��C3�JC4jC3��yn�+�3 Dff 2�A PB W4+@:�]o�W�� ���/�/P/'/ 9/K/]/o/�/�/�/�/ ?�/�/�/?#?5?�? Y?k?�?�?�o�?�?O �?6O!OZOlOWO�O�E s�?�?�?�O�O_�O �OL_#_5_G_Y_k_}_ �_�_�_ o�_�_�_o o1o~oUogo�o�o�o �o�owO D/A ze����O�o�o 
��o��R�)�;��� _�q����������ݏ �<��%�r�I�[�m� �������ǟٟ&�8� �\�G���k������� گů�����F�� /�A�S�e�w�Ŀ���� ��ѿ�����+�x� O�aϮυϗϩϻ��� ��,���b�t�ﯘ� �߼ߧ��������� :��C�U߂�Y�k�� ����������6�� �l�C�U�g�y����� ������ ��	- ?Q������ �@+dvQ� ������� *///%/r/I/[/�/ /�/�/�/�/�/&?�/ ?\?3?E?�?i?{?�? �?U�?�?"O4OOXO CO|OgO�O{��?�O �?�O�O0___f_=_ O_a_s_�_�_�_�_�_ o�_oo'o9oKo�o oo�o�o�o�o�o�O :%^I�������H�$DCS�S_SLAVE �U���	����z_4D�  	��AR_MENU V	� �j�|�������ď��BY�� ��~?�S�HOW 2W	� � �b�aG�Q� X�v���������П֏���� @�:�d�a� s����������߯� �*�$�N�K�]�o��� ����̯ɿۿ��� 8�5�G�Y�k�}Ϗ϶� ����������"��1� C�U�g�yߠϝ߯��� �����	��-�?�Q� c��s��������� ����)�;�M�t��� �������������� %7Ip�m�� ��������! 3ZWi���J ����//DA/ S/e/��/��/�/�/ �/�/?./+?=?O?v/ p?�/�?�?�?�?�?�? ?O'O9O`?ZO�?�O �O�O�O�O�OO�O_ #_JOD_nOk_}_�_�_ �_�_�O�_�_o4_.o X_Uogoyo�o�o�o�_ �o�o�ooBo?Q cu���o:��~�CFG X)��3�3q5p��FRA:\!�L�+�%04d.CS�V|	p}� ��qA g�CHo�z@v�	����3q�����́܏� ���4��JP����q�p1� �RC_�OUT Y���C��_C_�FSI ?i� .����� ��͟�����>�9� K�]���������ίɯ ۯ���#�5�^�Y� k�}�������ſ�� ���6�1�C�U�~�y� �ϝ����������	� �-�V�Q�c�uߞߙ� �߽��������.�)� ;�M�v�q����� �������%�N�I� [�m������������� ����&!3Eni {������� FASe�� ������// +/=/f/a/s/�/�/�/ �/�/�/�/??>?9? K?]?�?�?�?�?�?�? �?�?OO#O5O^OYO kO}O�O�O�O�O�O�O �O_6_1_C_U_~_y_ �_�_�_�_�_�_o	o o-oVoQocouo�o�o �o�o�o�o�o.) ;Mvq���� �����%�N�I� [�m���������ޏُ ���&�!�3�E�n�i� {�������ß՟���� ��F�A�S�e����� ����֯ѯ����� +�=�f�a�s������� ��Ϳ�����>�9� K�]φρϓϥ����� ������#�5�^�Y� k�}ߦߡ߳������� ���6�1�C�U�~�y� ������������	� �-�V�Q�c�u����� ����������.) ;Mvq���� ��%NI [m������ ��&/!/3/E/n/i/ {/�/�/�/�/�/�/�/�3�$DCS_C�_FSO ?����71 P ??T? }?x?�?�?�?�?�?�? OOO,OUOPObOtO �O�O�O�O�O�O�O_ -_(_:_L_u_p_�_�_ �_�_�_�_o oo$o MoHoZolo�o�o�o�o �o�o�o�o% 2D mhz����� ��
��E�@�R�d� ��������ՏЏ�� ��*�<�e�`�r��� ������̟����� =�8�J�\�������?_C_RPI4>F? �������3?�&��o����� >SLү@ d������%�7�`� [�m�Ϩϣϵ����� �����8�3�E�W߀� {ߍߟ���������� ��/�X�S�e�w�� �����������0� +�=�O�x�s������� ������'P K]o����� ���(#5Gp k}�����Q�� �/6/1/C/U/~/y/ �/�/�/�/�/�/?	? ?-?V?Q?c?u?�?�? �?�?�?�?�?O.O)O ;OMOvOqO�O�O�O�O �O�O___%_N_I_ [_m_�_�_�_�_�_�_ �_�_&o!o3oEonoio {o�o�o�o�o�o�o�o FASe�������>�NOC�ODE ZU���?�PRE_CHK \U���pA �p�< ��pU�]�o�U� 	 <Q����� ���ۏ�Ǐ�#��� �Y�k�E�����{�ş ן��ß����C�U� /�y�����s���ӯm� ��	���?��+�u� ��a�������ɿ�Ϳ ߿)�;��_�q�K�}� �ϝ������ω���%� ���[�m�Gߑߣ�}� ���߳����!���E� W�1�c��g�y����� ���������A�S�-� w���c����������� ��+=asM _������ '�]o	�� ����/#/� G/Y/3/e/�/i/{/�/ �/�/�/?�/?C?9 Ky?�?%?�?�?�?�? �?	O�?-O?OOKOuO OOaO�O�O�O�O�O�O �O)_____q_K_�_ �_a?�_�_�_�_o%o �_Io[o5oGo�o�o}o �o�o�o�o�o�oE W1{�g���_ ����/�A��M� w�Q�c���������� Ϗ�+���a�s�M� ��������ߟ��� '���3�]�7�I����� �ɯۯ������� G�Y�3�}���i���ſ ��������1�C��� +�yϋ�eϯ��ϛ��� ������-�?��c�u� Oߙ߫߅ߗ������� �)��M�_�U�G�� ��A����������� ��I�[�5����k��� ����������3E Q{q���] ����/Ae wQ������ �/+//7/a/;/M/ �/�/�/�/�/��/? '??K?]?7?�?�?m? ?�?�?�?�?O�?5O GO!O3O}O�OiO�O�O �O�O�O�/�O1_C_�O g_y_S_�_�_�_�_�_ �_�_o-oo9oco=o Oo�o�o�o�o�o�o�o __M_�ok� o������� �I�#�5����k��� Ǐ��ӏ��׏�3�E� �i�{�5c���ß�� ���ӟ�/�	��e� w�Q�������ѯ㯽� ϯ�+��O�a�;��� �����Ϳ߿y��� �!�K�%�7ρϓ�m� ���ϣ���������5� G�!�k�}�W߉߳ߩ� �����ߕ��1��� g�y�S������� �����-��Q�c�=� o���s��������� ����M_9�� o����� 7I#mYk� �����!/3/) /i/{//�/�/�/�/ �/�/�/?/?	?S?e? ??q?�?u?�?�?�?�? OO�?%OOOE/W/�O �O1O�O�O�O�O__ �O9_K_%_W_�_[_m_ �_�_�_�_�_�_o5o o!oko}oWo�o�omO �o�o�o�o1U gAS����� �	����Q�c�=� ����s���Ϗ�o��� ���;�M�'�Y���]� o���˟����۟� 7��#�m��Y����� �������!�3�ͯ ?�i�C�U�������տ �������	�S�e� ?ωϛ�uϧ��ϫϽ�������$DC�S_SGN ]�	�E��-����30-NOV�-25 19:4{4 ��29R՟20:27_�x��x� [}�t��q�т�xҚك�J����EƼÞ�o ��ǖ�  1ԿHOW ^	�? x�/��VERSION �=�V4.�5.2��EFLO�GIC 1_���  	������C��R�%�PROG_ENB  ���:�{�s�ULSE�  X��%�_�ACCLIM������d��WR�STJNT��E��-�EMO|�zя��$���INIT �`2����OPT?_SL ?		�	��
 	R57Y5��]�74b�6c�-7c�50��1����C���@�TO  �L��� �V�DKEX��dE�x�PATH A=ڇA\k}��H�CP_CLNTI�D ?�:� �D�ռ��IAG_GRP 2e	�����z�	� @�  
?ff?aG���B�  2��/�8[I@c����!�7@�z��@^�@
�!���mp2m1�5 890123�4567�����  ?���?�=q?��
�?޸R?�Q�?��?������(�?�z�����x�@�  A�_�Ap !7A�88_�B4��� ��L�x�
�@��@��\@�~�R@xQ�@�q�@j�H@�c�
@\��@U�@Mp���//'$�; �O)H���@Ct >d 9@4�/\)�@)� #t {@��/�/�/�/��/P'?���?����_ ?}p��?u?n{�?s ?\�Q��? ?2?D?V?h8�
�=?����0w5��z�H?p�h?��?^�R�?�?��?�?�?h8��t0����@�?��0�;@&O8OJO\O nOP'�$_�_Y_k_ �O?_�_�_�_�_�_s_ �_�_1oCo!ogoyoo �o��Bj"� �2{1�@^"?���f�t0��d"5!�
u4V��u"�B3t�AT>u��?@[q��@�`,=q�=b���=�E1>��J�>�n�>�{�H"<�o �z��s�q��� �zx�C�@<(�Uzҗ 4�� ����A@x�?*�o� �m*�P�b���tn����2���Ώ�����i>wJ��&�bN2��"��G�N��o@��@v���0����@�ffr!l ��s33���(��"�C�� ƒI��CH�)C.dBت"8"����'���"~�A?�&"�K����pf�B��@��p�������p��>6��N?y�I���!c?I������8?�#?�ߎ�TS��G��D<ŞB�?Q_DFxВ�@�����3��N��T����C��@���B�I� ����ÿ���ҿ俀�Ϥ��<�o��C�T_CONFIG� f��|��egY��ST�BF_TTS��
@����О�}���1��MAU������MS�W_CF��g� � # ��OCVIE�W��h!�-�� �s߅ߗߩ߻��ߟ� a�����,�>�P��� t�������]��� ��(�:�L�^���� ����������k�  $6HZ��~�� ����y 2 DVh�����X��v�RC�i���!���/S/B/w/�f/�/�/�/��SBL�_FAULT �j*6��!GPMS�K���'��TDIAOG k��-�������UD1�: 6789012345I2��=1����P\υ?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�Od696���r�
t?�O|�TREC	P"?4:
B44_[7�� s?p_�_�_�_�_�_�_ �_ oo$o6oHoZolo�~o�o�O�O�O�o7�U�MP_OPTIO2=��.�aTR���:�)uPME���Y_TEMP  �È�3BC�rgp�B�QtUNI�����gq�YN_BR�K lL�7�EDITOR�a�a@�r�_
PENT 1m�)  ,&?TELEOP^P �z���pPSNA��:�&MTPG �p+�=��/��I�z��� ��ۏ����5�� Y�k�R���v���ş�� �П����C�*�g� N�v�������������ޯ��?�Q���E�MGDI_STA�zuV�gq�uNC_I?NFO 1n!��b���X�������솳n�1o!� �P�o����
�d�o U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫��� u�� ��
��*�B�*�P�b� t����������� ��(�:�L�^�p��� ������2������� 9�CUgy�� �����	- ?Qcu���� ����//1;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?��?�?�? O)/OEOWOiO{O�O �O�O�O�O�O�O__ /_A_S_e_w_�_�_�_ �?�?�_�_o�_3O=o Ooaoso�o�o�o�o�o �o�o'9K] o����_�_�� ��+o5�G�Y�k�}� ������ŏ׏���� �1�C�U�g�y����� ���ӟ���	�#�-� ?�Q�c�u��������� ϯ����)�;�M� _�q���������˿ݿ ����7�I�[�m� ϑϣϵ��������� �!�3�E�W�i�{ߍ� �߹����������%� /�A�S�e�w���� ����������+�=� O�a�s����������� �����'9K] o������� �#5GYk} �	������ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?��? �?�?�?/O)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�?�_�_�_�_O �_!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��_�_ ����o�+�=� O�a�s���������͏ ߏ���'�9�K�]� o�������ɟ۟� ��#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߝ��߹����� �����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ����������� /ASew��� ����+= Oas������� ���//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?� ��?�?�?�?��?O O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�?�_�_�_ �_�?�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m �_u����_�� �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e������ ��u������+�=� O�a�s���������ͯ ߯���'�9�K�]� w���������ɿ�� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g߁��ߝ� ����ۿ����	��-� ?�Q�c�u����� ��������)�;�M� _�y߃����������� ��%7I[m ������� !3EWq�c� ��������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?i{�?�?�?�?� �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_�?s?}_ �_�_�_�?�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qk_u����_ �����)�;�M� _�q���������ˏݏ ���%�7�I�cQ� ��������ٟ��� �!�3�E�W�i�{��� ����ïկ������/�A�[� �$EN�ETMODE 1�p��� W k�k�f������j�OATCF�G q��e��Ѵ��C���DATA 1rw�uӰ���*	ρ*��'�9�K�]�l�dlύ�e��ϻ��� ������'ߡϳ�]� o߁ߓߥ߷�1���U� ���#�5�G�Y����� ������������u� ��1�C�U�g�y���� ��)�������	- ����cu������j�RPOST_KLO��t�[
׶�#5Gi�RROoR_PR� %w��%L�XTABL/E  w�ȟ�����RSEV_�NUM ��  ����  �_�AUTO_ENB�  ���X_N�O5! uw����"  *�x �Jx �x �x + +w �/�/�/Q$FLTR=/O&HIS#]��J+_ALM 1v.w� �[x,e�+�/Q?c?u?�?�?�?�/_"W   �w�v!���:j�TC�P_VER !�w�!x�?$EXT�� _REQ�&�H)BCSIZKO=DSkTKhIf%�?B�TOL  ]D�z�"�A =D_BWD�0�@�&�A��v�CDI�A wķ����]�KSTEP��O�Oj�POP_D�O�Oh�FDR_G�RP 1xw��!d� 	�?�_��yPs��Y�Q'�M�"���l��T� ����V�yS�_�]yPA8���B/}A՚��A�@�d��B3���]]An��^�Qab�� oEo�_Bo{ofo�o�o��o�o@5�@"���@ P�>�����n
 M �� a�a�bB�� �o(2�o�oZE~�]y@`�t@S33�u�]@�q�g��yP�F@ ��|yPG��  @�Fg�f�C�8RL��]?��  h��6�X�����875t���5���5`+���~����3�� {� �A$�� M6���5��FEATURE� y���@���HandlingTool ��]Engli�sh Dicti�onary�4Dw St��ard���Analog �I/O>�G�gle� ShiftZ�u�to Softw�are Upda�te�matic Backup����ground �Edit ��Ca�meraU�FY�CnrRndIm����ommon calib UI���nˑ�Moni�tor$�tr�R�eliabn��D�HCP �[�ata Acquis3�~\�iagnos���R�v�isplay~ΑLicensZ��`�ocument? Viewe?�^��ual Chec�k Safety���hancedh���s�Frܐ��xt. DIO� /�fi��@�en]d�Err>�L���\�4�s[�rP�K� ��@
�FCTN M�enu��vZ���T�P In��fac<ĵ�GigE־��Đp Mask �Exc�g=�HT�԰Proxy S�v��igh-S;pe�Ski�� ����O�mmunicn��onsV�ur���q�V�ײconn�ect 2��nc=rְstru!��ʒ��eۡ��J��X�K�AREL Cmd7. L�ua��ÿRun-Ti<�E�nv�Ȟ�el +:��s��S/W�ƥ����r�Book(System)
�MACROs,M�?/Offseu�p�aHO���o�u�MR8��4���MechSt�op+�t����p�im�q���x�R������odo�witch��ӟ�.��4�Op�tmF��,�fil�䬳�g��p�ult�i-T�Γ�PC�M fun�Ǽ�o���������Regi�e�rq���riݠF����S�Num S�el��/�:� Ad�jua�*�W�q�h�t�atu��ߪ�R�DM Robot>�scove'����ea��<�Freq� Anlyq�Re�m��O�n5�����S�ervoO�!��S�NPX b-�v�SN԰Cliܡ?r��Libr&�_�� ���q +oJ�t��sGsag��X�@ �����	�@/Iս�M�ILIB��P OFirm���P���AccŐ͛TPT9Xk��eln��������orqu>o�imula=��|u(�Pa&��ĐtX�B�&+�ev.�成ri��TUSB port ��iPf�aݠ&R �EVNT� nexcept�����X%5��VC�rl�c���V���"�%q��+SR SCN�/S�GE�/�%UI	�Web Pl��>���A43��ۡ��ZD?T Applj�
�{1EOAT����x&0?�7Grid�񸾡�=�?iR�".�5� F���/גRX-�10iA/L�?A�larm Cau�se/��ed(�A�ll Smoot�h5���C�scii<+�V�Load䠌J�Upl�@w�toS� ��rityAv�oidM(�s7�t�@�ycn�����_�CS+���.3 c��XJo��� -T3_H�.RX��U����Xcollabo����RA�:�.9D���in���NR�THI
�On��e Hel����ֿ������1trU�ROS Eth$��A������;,�G �B�,�|HUpV�%�W�t ԰�_iRS�ݐ��64MB DRA9M�o�cFRO���L8F FlD�����22M �A:�opm�ԕ1ex@V�
�sh�q�"�wce�u��p��|�tyn�sA�
�%�r ����J��^�.v� P)Q/sbS�`���O�N��mai��U�h��R�q�T1�^cFC+Ԍ%̋Fs9�pˌk̋��Typ߽�FC%�hױV�N Sp�ForްK��Ԭ��lu!����cp�PG� j�֡�RJ�[L`Sup"}��֐�f��crFP��lu�� ��al�����r ��i�
q�4@а��uest,IMPLE ׀6*|HZ�p��c0�BTea(�8|���$rtu���V��9HMI�¤��U;IFc�pono2D�BC�:�L�y�p��� ������ʿܿ	� �� ?�6�H�u�l�~ϫϢ� ����������;�2� D�q�h�zߧߞ߰��� �����
�7�.�@�m� d�v��������� ���3�*�<�i�`�r� �������������� /&8e\n�� ������+" 4aXj���� ����'//0/]/ T/f/�/�/�/�/�/�/ �/�/#??,?Y?P?b? �?�?�?�?�?�?�?�? OO(OUOLO^O�O�O �O�O�O�O�O�O__ $_Q_H_Z_�_~_�_�_ �_�_�_�_oo oMo DoVo�ozo�o�o�o�o �o�o
I@R v������ ���E�<�N�{�r� ������Տ̏ޏ�� �A�8�J�w�n����� ��џȟڟ����=� 4�F�s�j�|�����ͯ į֯����9�0�B� o�f�x�����ɿ��ҿ �����5�,�>�k�b� tφϘ��ϼ������� �1�(�:�g�^�p߂� ���߸������� �-� $�6�c�Z�l�~��� ����������)� �2� _�V�h�z��������� ������%.[R dv������ �!*WN`r �������/ /&/S/J/\/n/�/�/ �/�/�/�/�/??"? O?F?X?j?|?�?�?�? �?�?�?OOOKOBO TOfOxO�O�O�O�O�O �O___G_>_P_b_ t_�_�_�_�_�_�_o ooCo:oLo^opo�o �o�o�o�o�o	  ?6HZl��� ������;�2� D�V�h�������ˏ ԏ���
�7�.�@�R� d�������ǟ��П�� ���3�*�<�N�`��� ����ï��̯���� /�&�8�J�\������� ����ȿ�����+�"� 4�F�Xυ�|ώϻϲ� ��������'��0�B� T߁�xߊ߷߮����� ����#��,�>�P�}� t����������� ��(�:�L�y�p��� ������������ $6Hul~������  �H552��2�1R7850�J614AT�UP'545'6�VCAMCR�IbUIF'28ncNRE52VwR63SCH�LIC�DOCV��CSU869z'02EIOC��4R69VES�ET?UJ7UR{68MASK�PRXY{7OCO#(3?+ &m3j&J6%53��H�(LCHR&OP�LG?0�&MHCuRS&S�'MCS>�0.'552MDS�W+7u'OPu'MP�Rv&��(0&PCMzR0q7+ 2� ��'51J51�80nJPRS"'69j&�FRDbFREQnMCN93&�SNBA��'SH�LBFM1G�82�&HTC>TMI�L�TPA�T7PTXcFELF� ��8J95n�TUTv'95j&wUEV"&UECR&wUFRbVCC
X�O�&VIPnFCS�C�FCSG��I�WEB>HTT�>R6��H;RVC�GiWIGQWIPGmS�VRCnFDGu'�H7�7R66J5t'R�8R51
(�6�(2�(5V�J8�86�L=I% ږ84g662R6�4NVD"&R6n�'R84�g79�(�4�S5i'J76�j&D0�gF xRT�SFCR�gCRX�v&CLIZ8ICMqS�Sp>STYnG6)7CTO>���7�NNj&ORS��&C &FCB�F�CF�7CH>FC�R"&FCI�VFCR�'J�PO7GBfM�8�OLaxENDS&L]U�&CPR�7LW�S�xC�STxTE�gS60FVR6�IN�7IHaF� я�����+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯۯ��� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q����������� ��%�7�I�[�m�� �������������� !3EWi{�� �����/ ASew���� ���//+/=/O/ a/s/�/�/�/�/�/�/ �/??'?9?K?]?o? �?�?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_ �_�_�_�_	oo-o?o Qocouo�o�o�o�o�o �o�o);M_ q������� ��%�7�I�[�m���������Ǐُ� � H552���21�R78��50�J614��ATUP7�54�57�6�VCAM��CRI��UIFv7�28��NRE��52v�R63�S�CH�LICƚDwOCV�CSU��8697�0F�EI�OCǛ4�R69�v�ESETW�u�J�7u�R68�MA{SK�PRXY��]7�OCO��3W�h���6�3�J65��536�H$�LCH^ƪOPLGW�0��MHCRǪS��MkCSV�0��55F��MDSW���OP���MPR���6�0n6�PCM��R0E˰��F���6�51f�5u1��0f�PRS���69�FRD��FwREQ�MCN�{936�SNBAכ^%�SHLB�ME�t�ּ26�HTCV��TMIL�6�TP�AV�TPTX��ELړ�6�8%�#��wJ95��TUT���95�UEV��U�ECƪUFR��V�CCf�O��VIP��CSC��CSGtƚ$�I�WEBV�7HTTV�R6՜��lS���CG��IG��oIPGS'�RC���DG��H7��R6�6f�5�u�R��R�51f�6�2�5�v�#�J׼��6��L�U�5�s�v�4��66�F�R64�NVDv��R6��R84�k79�4��S5嫷J76�D0uFnRTS&�CR�wCRX��CLI&̎e�CMSV�sV�S�TY��6�CTOhV�#�V�75�NN��ORS����6�FC�BV�FCF��CH�V�FCR��FCI�F�FC��J#��G�
M��OL�EN�DǪLU��CPR���Lu�S�C$�SvtTE�S60��FVRV�IN��IH���m??�?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� ������������ '9K]o��� �����#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s����������͏ߏ��STD�LANG���0�B� T�f�x���������ҟ �����,�>�P�b� t���������ί�� ��(�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢ� ����������� �2� D�V�h�zߌߞ߰����RBT
�OPTN ������'�9�K�]� o�����������DPN	���)�;� M�_�q����������� ����%7I[ m������ ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ� ����������'�9� K�]�o߁ߓߥ߷��� �������#�5�G�Y� k�}���������� ����1�C�U�g�y� ��������������	 -?Qc�f�������99���$FEAT_�ADD ?	����  	�#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙπ�Ͻ��������D�EMO y   �L�B� T߁�xߊ߷߮����� ������G�>�P�}� t����������� ��C�:�L�y�p��� ������������ ?6Hul~�� ����;2 Dqhz���� �� /
/7/./@/m/ d/v/�/�/�/�/�/�/ �/?3?*?<?i?`?r? �?�?�?�?�?�?�?O /O&O8OeO\OnO�O�O �O�O�O�O�O�O+_"_ 4_a_X_j_�_�_�_�_ �_�_�_�_'oo0o]o Tofo�o�o�o�o�o�o �o�o#,YPb �������� ��(�U�L�^����� ������ʏ���� $�Q�H�Z���~����� ��Ɵ����� �M� D�V���z�������¯ ܯ��
��I�@�R� �v���������ؿ� ���E�<�N�{�r� �ϱϨϺ������� �A�8�J�w�n߀߭� �߶���������=� 4�F�s�j�|���� ��������9�0�B� o�f�x����������� ����5,>kb t������� 1(:g^p� ������ /-/ $/6/c/Z/l/�/�/�/ �/�/�/�/�/)? ?2? _?V?h?�?�?�?�?�? �?�?�?%OO.O[ORO dO�O�O�O�O�O�O�O �O!__*_W_N_`_�_ �_�_�_�_�_�_�_o o&oSoJo\o�o�o�o �o�o�o�o�o" OFX�|��� ������K�B� T���x�������ۏҏ ����G�>�P�}� t�������ןΟ��� ��C�:�L�y�p��� ����ӯʯܯ	� �� ?�6�H�u�l�~����� Ͽƿؿ����;�2� D�q�h�zϔϞ����� �����
�7�.�@�m� d�vߐߚ��߾����� ���3�*�<�i�`�r� ������������� /�&�8�e�\�n����� ������������+" 4aXj���� ����'0] Tf������ ��#//,/Y/P/b/ |/�/�/�/�/�/�/�/ ??(?U?L?^?x?�? �?�?�?�?�?�?OO $OQOHOZOtO~O�O�O �O�O�O�O__ _M_ D_V_p_z_�_�_�_�_ �_�_o
ooIo@oRo lovo�o�o�o�o�o�o E<Nhr �������� �A�8�J�d�n����� ��яȏڏ����=� 4�F�`�j�������͟ ğ֟����9�0�B� \�f�������ɯ��ү �����5�,�>�X�b� ������ſ��ο��� �1�(�:�T�^ϋς� ���ϸ������� �-� $�6�P�Z߇�~ߐ߽� ����������)� �2� L�V��z������ ������%��.�H�R� �v������������� ��!*DN{r ������� &@Jwn�� �����//"/ </F/s/j/|/�/�/�/ �/�/�/???8?B? o?f?x?�?�?�?�?�? �?OOO4O>OkObO tO�O�O�O�O�O�O_|_0]  'X F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ����������
��.�  /�)�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o�o "4FXj|�� �������0� B�T�f�x��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@� R�d�v߈ߚ߬߾��� ������*�<�N�`� r����������� ��&�8�J�\�n��� �������������� "4FXj|�� �����0 BTfx���� ���//,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�?�? O O$O6OHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Rodovo�o�o�o�o�o �o�o*<N` r������� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P� b�t���������ο� ���(�:�L�^�p� �ϔϦϸ������� �(�$�4�8�+�N� `�r߄ߖߨߺ����� ����&�8�J�\�n� ������������� �"�4�F�X�j�|��� ������������ 0BTfx��� ����,> Pbt����� ��//(/:/L/^/ p/�/�/�/�/�/�/�/  ??$?6?H?Z?l?~? �?�?�?�?�?�?�?O  O2ODOVOhOzO�O�O �O�O�O�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ� ����������
��.� @�R�d�v����� ��������*�<�N� `�r������������� ��&8J\n �������� "4FXj|� ������// 0/B/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?t?�?�?�?�?�? �?�?OO(O:OLO^O pO�O�O�O�O�O�O�O� __$_6Y�$FE�AT_DEMOIoN  ;T�fP��<PNTINDE�X[[jQ�NPIL�ECOMP z�����Q�iRIU�PSETUPo2 {�U�R?�  N �Q�S�_AP2BCK �1|�Y  �)7Xok%�_8o<P�P&oco9U�_�oo �oBo�o�oxo�o1 C�og�o��,� P�����?�� L�u����(���Ϗ^� 󏂏�)���M�܏q� �����6�˟Z�؟� ��%���I�[���� ����D�ٯh������ 3�¯W��d������ @�տ�v�Ϛ�/�A� пe����ϛ�*Ͽ�N� ��r���ߨ�=���a� s�ߗ�&߻���\��� ���'��K���o��� |��4���X������ #���G�Y���}���� ��B���f�����1t�Y�PP�_ 2�P*.VR8���*��������l PC���F'R6:�2�V�TzPz�w��]PG���*.F�o/��	�:,8�^/�STMi/�/ /�-M/�/�H�/?�'?�/�/g?�GIFq?�?�%�?pD?V?�?�JPG�?�O�%O�?�?oO�
JSyO�O��5C�OMO�%
JavaSc�ript�O�?CS�O&_�&_�O %�Cascadin�g Style ?SheetsR_���
ARGNAME�.DT�_��� \@�_S_�A�T�_�_�P�DISP*�_����To�_�QLaZooCLLB.ZIwo,2o$ :\�a\�o�i��ACollab�o�o�o
TPEI?NS.XML�_�:\![o�QCus�tom Tool�barbiPAS�SWORDQo��FRS:\�dB`�Password Config� ��/��(�e���� ����N��r����� =�̏a������&��� J���񟀟���9�K� ڟo�������4�ɯX� �|���#���G�֯@� }����0�ſ׿f��� ���1���U��y�� ϯ�>���b���	ߘ� -߼�Q�c��χ�߫� ��L���p��ߦ�;� ��_���X��$��H� ����~����7�I��� m���� �2���V��� z���!��E��i{ 
�.��d�� ��S�wp �<�`�/�+/ �O/a/��//�/8/ J/�/n/?�/�/9?�/ ]?�/�?�?"?�?F?�? �?|?O�?5O�?�?kO �?�OO�O�OTO�OxO __�OC_�Og_y__ �_,_�_P_b_�_�_o �_oQo�_uoo�o�o :o�o^o�o�o)�o M�o�o��6� �l��%�7��[� ���� ���D�ُh� z����3�,�i��� �����ßR��v�������$FILE�_DGBCK 1�|������ < ��)
SUMMAR�Y.DG!�͜M�D:U���ِD�iag Summ�ary����
CONSLOG��n����ٯ���Console log����	TPACCN��t�%\�����T�P Accoun�tin;���FR�6:IPKDMPO.ZIPͿј
��ϥ���Excep�tion"�ӻ��MEMCHECK���������-�Mem�ory Data|����>n )��RIPE�~ϐ�%���%�� Pa?cket L:����L�$�c���ST�AT��߭� �%A�Stat�us��^�	FTP�����	��/�m�ment TBD�2�^� >I)E?THERNEw�
��d�u�﨡Eth�ernJ�1�fig�uraAϩ��DCSVRF&���7������ veri?fy all:���� 4��DIF�F/��'���;�Q�d�iff��r�d���CHG01������A�����it�2���2 70���fx�3���I ��p�VTRNDIAG.LSu�&8���� O�pe��L� ��no�stic��GϿ)VDEV�D�AT�������Vis�Devisce�+IMG���,/>/�/:�i$I�magu/+UP� ES/�/FR�S:\?Z=��U�pdates L�istZ?��� FLEXEVEN��в/�/�?���1 UIF EvM�M����-vZ)CR?SENSPK�/˞��\!O���CR�_TAOR_PEA�KbOͩPSRBW�LD.CM�O͜�E2�O\?.�PS_R?OBOWELS���:GIG��@_�?d_>��GigE�(O~��N�@�)UQHADOW__D_V_��_��Shado�w Change�����1dt�RRCMERR�_�_�_oo���4`CFG E�rroro tai}lo MA�k�CMSGLIBgo�No`o�o|R�e��z0iyc�o�a�)�`�ZD0_O�os���ZD�Pad�l= �RNOTI�R�d���Noti�fic����,�AG��P�ӟt����� ����Ώ]�����(� ��L�^�폂������ G�ܟk� ����6�ş Z��~������C�د �y����2�D�ӯh� �������¿Q��u� 
�ϫ�@�Ͽd�v�� ��)Ͼ���_��σ�� ��%�N���r�ߖߨ� 7���[�����&�� J�\��߀���3�� ��i����"�4���X� ��|������A����� w���0��=f�� ���O�s �>�bt� '�K���/� :/L/�p/��/�/5/ �/Y/�/ ?�/$?�/H? �/U?~??�?1?�?�? g?�?�? O2O�?VO�? zO�OO�O?O�OcO�O 
_�O._�OR_d_�O�_ _�_�_M_�_q_oo �_<o�_`o�_mo�o%o �oIo�o�oo�o8 J�on�o��3� W�{�"��F�� j�|����/�ď֏e�������0��$FI�LE_FRSPRT  ������?��MDONLY 1�|S�� 
 ��)MD:_V�DAEXTP.Z�ZZ1�⏹�ț�6%NO Ba�ck file <���S�6P��� ��>��K�t�����'� ��ί]�򯁯�(��� L�ۯp������5�ʿ Y�׿ Ϗ�$ϳ�H�Z� �~�Ϣϴ�C���g� ��ߝ�2���V���c� ��߰�?�����u�
� ��.�@���d��߈��~C�VISBCKq�|[���*.VD��|��S�FR:\���ION\DATA�\��v�S�Vision VD� ��Y�k����y�� B�����x���1C ��g���,�P ����?�P u�(��^� �/��M/�q/�/ >/�/6/�/Z/�/?�/ %?�/I?[?�/??�?�2?D?�?9�LUI_�CONFIG �}S����; '$ �3v�{S�;O�MO_OqO�O�O�I#@|x�?�O�O�O__%\ �OH_Z_l_~_�_'_�_ �_�_�_�_o�_2oDo Vohozo�o#o�o�o�o �o�o
�o.@Rd v������ ��*�<�N�`�r��� �����̏ޏ����� &�8�J�\�n������ ��ȟڟ쟃���"�4� F�X�j��������į ֯����0�B�T� f�����������ҿ� {���,�>�P�b��� �ϘϪϼ�����w�� �(�:�L�^��ςߔ� �߸�����s� ��$� 6�H���Y�~���� ��]������ �2�D� ��h�z���������Y� ����
.@��d v����U�� *<�`r� ���Q��// &/8/�\/n/�/�/�/ ;/�/�/�/�/?"?�/ F?X?j?|?�?�?7?�? �?�?�?OO�?BOTO fOxO�O�O3O�O�O�O �O__�O>_P_b_t_ �_�_/_�_�_�_�_o o�_:oLo^opo�o�o>$h  x�o�c��$FLUI_D�ATA ~�����a�(a�dRESULT� 3�ep ��T�/wi�zard/gui�ded/step�s/Expert �o=Oas��������z�C�ontinue �with Gpance�:�L�^�p� ��������ʏ܏� �� �b-�a�e�0 �0`��c�a6?��ps��� ������ҟ����� ,�>�P��0ow����� ����ѯ�����+��=�O�a�?�1�C�U�e�cllbs�ֿ� ����0�B�T�f�x� �Ϝ�[���������� �,�>�P�b�t߆ߘ�@��i�{��ߟ�]�e�rip(pſ-�?�Q� c�u��������� ����)�;�M�_�q� �������������� ������`�e�#p�TimeUS/DST	��������!3E�Enabl(�y� ������	//(-/?/Q/�b�)0�/M_q24|�/ �/??)?;?M?_?q? �?�?Tf�?�?�?O O%O7OIO[OmOO�O �Ob/t/�/�/Z�"q?Region�O5_ G_Y_k_}_�_�_�_�_��_�_�America!�#o5oGoYo ko}o�o�o�o�o�o�o��Ay�O�O3�O_~qEditor�o ����������+�=� � Tou�ch Panel� rs (reco/mmenp�)K��� ����Ə؏���� �2�D�|�%��I|[qacceso ܟ� ��$�6�H�Z��l�~�����Con�nect to Network�� ֯�����0�B�T��f�x�����x��@���}����,!��s I�ntroduct !_4�F�X�j�|ώϠ� �����������0� B�T�f�xߊߜ߮��������� ɿ� �"�i�{���� ����������/�A�  �e�w����������������+=�H�3��+�O� ���� 2D Vhz�K���� ��
//./@/R/d/ v/�/�/Yk}�/� ??*?<?N?`?r?�? �?�?�?�?�?��?O &O8OJO\OnO�O�O�O �O�O�O�O�/_�/1_ �/X_j_|_�_�_�_�_ �_�_�_oo0oBoS_ foxo�o�o�o�o�o�o �o,>�O_!_ �E_������ �(�:�L�^�p����� So��ʏ܏� ��$� 6�H�Z�l�~���O�� s՟���� �2�D� V�h�z�������¯ԯ 毥�
��.�@�R�d� v���������п⿡� �ş'�9���`�rτ� �ϨϺ��������� &�8���\�n߀ߒߤ� �����������"�4� �=��a��Mϲ��� ��������0�B�T� f�x���I߮������� ��,>Pbt �E��i���� (:L^p�� ������ //$/ 6/H/Z/l/~/�/�/�/ �/�/����/?� V?h?z?�?�?�?�?�? �?�?
OO.O�ROdO vO�O�O�O�O�O�O�O __*_<_�/??�_ C?�_�_�_�_�_oo &o8oJo\ono�o?O�o �o�o�o�o�o"4 FXj|�M___q_ ��_���0�B�T� f�x���������ҏ�o ���,�>�P�b�t� ��������Ο���� �%��L�^�p����� ����ʯܯ� ��$� 6�G�Z�l�~������� ƿؿ���� �2�� S��w�9��ϰ����� ����
��.�@�R�d� v߈�G��߾������� ��*�<�N�`�r�� Cϥ�g���ύ��� &�8�J�\�n������� ����������"4 FXj|���� ������-��T fx������ �//,/��P/b/t/ �/�/�/�/�/�/�/? ?(?�1U??A �?�?�?�?�? OO$O 6OHOZOlO~O=/�O�O �O�O�O�O_ _2_D_ V_h_z_9?�?]?�_�_ �?�_
oo.o@oRodo vo�o�o�o�o�o�O�o *<N`r� �����_�_�_�_ #��_J�\�n������� ��ȏڏ����"��o F�X�j�|�������ğ ֟�����0��� �u�7�������ү� ����,�>�P�b�t� 3�������ο��� �(�:�L�^�pς�A� S�e��ω��� ��$� 6�H�Z�l�~ߐߢߴ� �߅������ �2�D� V�h�z�������� ��������@�R�d� v��������������� *;�N`r� ������ &��G	�k-��� �����/"/4/ F/X/j/|/;�/�/�/ �/�/�/??0?B?T? f?x?7�?[�?�? �?OO,O>OPObOtO �O�O�O�O�O�/�O_ _(_:_L_^_p_�_�_ �_�_�_�?�_�?o!o �OHoZolo~o�o�o�o �o�o�o�o �OD Vhz����� ��
���_%o�_I� s�5o������Џ�� ��*�<�N�`�r�1 ������̟ޟ��� &�8�J�\�n�-�w�Q� ��ů������"�4� F�X�j�|�������Ŀ �������0�B�T� f�xϊϜϮ������ �����ٯ>�P�b�t� �ߘߪ߼�������� �տ:�L�^�p��� ��������� ��$� �����i�+ߐ����� �������� 2D Vh'����� ��
.@Rd v5�G�Y��}��� //*/</N/`/r/�/ �/�/�/y�/�/?? &?8?J?\?n?�?�?�? �?�?��?�O�4O FOXOjO|O�O�O�O�O �O�O�O__/OB_T_ f_x_�_�_�_�_�_�_ �_oo�?;o�?_o!O �o�o�o�o�o�o�o (:L^p/_� ����� ��$� 6�H�Z�l�+o��Oo�� sou����� �2�D� V�h�z�������� ���
��.�@�R�d� v���������}�߯�� ��ٟ<�N�`�r��� ������̿޿��� ӟ8�J�\�nπϒϤ� �����������ϯ� �=�g�)��ߠ߲��� ��������0�B�T� f�%ϊ��������� ����,�>�P�b�!� k�Eߏ���{����� (:L^p�� ��w��� $ 6HZl~��� s�������/��2/D/ V/h/z/�/�/�/�/�/ �/�/
?�.?@?R?d? v?�?�?�?�?�?�?�? OO���]O/�O �O�O�O�O�O�O__ &_8_J_\_?�_�_�_ �_�_�_�_�_o"o4o FoXojo)O;OMO�oqO �o�o�o0BT fx���m_�� ���,�>�P�b�t� ��������{oݏ�o� �o(�:�L�^�p����� ����ʟܟ� ��#� 6�H�Z�l�~������� Ưد����͏/�� S��z�������¿Կ ���
��.�@�R�d� #��ϚϬϾ������� ��*�<�N�`���� C���g�i������� &�8�J�\�n���� ��u��������"�4� F�X�j�|�������q� ������	��0BT fx������ ���,>Pbt �������/ ����1/[/�/�/ �/�/�/�/�/ ??$? 6?H?Z?~?�?�?�? �?�?�?�?O O2ODO VO/_/9/�O�Oo/�O �O�O
__._@_R_d_ v_�_�_�_k?�_�_�_ oo*o<oNo`oro�o �o�ogOyO�O�O�o�O &8J\n��� ������_"�4� F�X�j�|�������ď ֏�����o�o�oQ� x���������ҟ� ����,�>�P��t� ��������ί��� �(�:�L�^��/�A� ��e�ʿܿ� ��$� 6�H�Z�l�~ϐϢ�a� ��������� �2�D� V�h�zߌߞ߰�o��� ���߷��.�@�R�d� v����������� ��*�<�N�`�r��� �������������� #��G	�n��� �����"4 FX�|���� ���//0/B/T/ u/7�/[]/�/�/ �/??,?>?P?b?t? �?�?�?i�?�?�?O O(O:OLO^OpO�O�O �Oe/�O�/�O�O�?$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_�? o2oDo Vohozo�o�o�o�o�o �o�o�O_�O%O_ v������� ��*�<�N�or��� ������̏ޏ���� &�8�J�	S-w��� cȟڟ����"�4� F�X�j�|�����_�į ֯�����0�B�T� f�x�����[�m���� 󿵟�,�>�P�b�t� �ϘϪϼ������ϱ� �(�:�L�^�p߂ߔ� �߸������� ￿ѿ �E��l�~���� ��������� �2�D� �h�z����������� ����
.@R� #�5�Y���� *<N`r� �U�����// &/8/J/\/n/�/�/�/ c�/��/�?"?4? F?X?j?|?�?�?�?�? �?�?�??O0OBOTO fOxO�O�O�O�O�O�O �O�/_�/;_�/b_t_ �_�_�_�_�_�_�_o o(o:oLoOpo�o�o �o�o�o�o�o $ 6H_i+_�O_Q ����� �2�D� V�h�z�����]oԏ ���
��.�@�R�d� v�����Y��}ߟ� ���*�<�N�`�r��� ������̯ޯ𯯏� &�8�J�\�n������� ��ȿڿ쿫���ϟ� C��j�|ώϠϲ��� ��������0�B�� f�xߊߜ߮������� ����,�>���G�!� k��Wϼ�������� �(�:�L�^�p����� S߸������� $ 6HZl~�O�a� s����� 2D Vhz����� ���
//./@/R/d/ v/�/�/�/�/�/�/�/ ���9?�`?r?�? �?�?�?�?�?�?OO &O8O�\OnO�O�O�O �O�O�O�O�O_"_4_ F_??)?�_M?�_�_ �_�_�_oo0oBoTo foxo�oIO�o�o�o�o �o,>Pbt ��W_�{_��_� �(�:�L�^�p����� ����ʏ܏���$� 6�H�Z�l�~������� Ɵ؟꟩��/�� V�h�z�������¯ԯ ���
��.�@���d� v���������п��� ��*�<���]���� C�EϺ��������� &�8�J�\�n߀ߒ�Q� �����������"�4� F�X�j�|��Mϯ�q� �������0�B�T� f�x������������� ��,>Pbt ���������� ��7��^p�� ����� //$/ 6/��Z/l/~/�/�/�/ �/�/�/�/? ?2?� ;_?�?K�?�?�? �?�?
OO.O@OROdO vO�OG/�O�O�O�O�O __*_<_N_`_r_�_ C?U?g?y?�_�?oo &o8oJo\ono�o�o�o �o�o�o�O�o"4 FXj|���� ���_�_�_-��_T� f�x���������ҏ� ����,��oP�b�t� ��������Ο���� �(�:�����A� ����ʯܯ� ��$� 6�H�Z�l�~�=����� ƿؿ���� �2�D� V�h�zό�K���o��� ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�� ������������� #���J�\�n������� ����������"4 ��Xj|���� ���0��Q �u7�9���� �//,/>/P/b/t/ �/E�/�/�/�/�/? ?(?:?L?^?p?�?A �?e�?�?�/ OO$O 6OHOZOlO~O�O�O�O �O�O�/�O_ _2_D_ V_h_z_�_�_�_�_�_ �?�?�?o+o�?Rodo vo�o�o�o�o�o�o�o *�ON`r� �������� &��_/o	oS�}�?o�� ��ȏڏ����"�4� F�X�j�|�;����ğ ֟�����0�B�T� f�x�7�I�[�m�ϯ�� ����,�>�P�b�t� ��������ο���� �(�:�L�^�pςϔ� �ϸ����ϛ�����!� �H�Z�l�~ߐߢߴ� ��������� �߿D� V�h�z�������� ����
��.������ s�5ߚ����������� *<N`r1� ������ &8J\n�?�� c������/"/4/ F/X/j/|/�/�/�/�/ �/��/??0?B?T? f?x?�?�?�?�?�?� �?�O�>OPObOtO �O�O�O�O�O�O�O_ _(_�/L_^_p_�_�_ �_�_�_�_�_ oo$o �?EoOio+O-o�o�o �o�o�o�o 2D Vhz9_���� ��
��.�@�R�d� v�5o��Yo��͏�� ��*�<�N�`�r��� ������̟���� &�8�J�\�n������� ��ȯ��я������ F�X�j�|�������Ŀ ֿ�����ݟB�T� f�xϊϜϮ������� ����ٯ#���G�q� 3��ߪ߼�������� �(�:�L�^�p�/ϔ� ��������� ��$� 6�H�Z�l�+�=�O�a� �������� 2D Vhz������ ��
.@Rd v��������� ��/��</N/`/r/�/ �/�/�/�/�/�/?? �8?J?\?n?�?�?�? �?�?�?�?�?O"O� �/gO)/�O�O�O�O �O�O�O__0_B_T_ f_%?w_�_�_�_�_�_ �_oo,o>oPoboto 3O�oWO�o{O�o�o (:L^p�� ����o� ��$� 6�H�Z�l�~������� Ə�o珩o��o2�D� V�h�z�������ԟ ���
���@�R�d� v���������Я��� ��׏9���]��!� ������̿޿��� &�8�J�\�n�-��Ϥ� �����������"�4� F�X�j�)���M����� ��������0�B�T� f�x��������� ����,�>�P�b�t� ��������{��ߟ��� ��:L^p�� ����� �� 6HZl~��� ����/���� ;/e/'�/�/�/�/�/ �/�/
??.?@?R?d? #�?�?�?�?�?�?�? OO*O<ONO`O/1/ C/U/�Oy/�O�O__ &_8_J_\_n_�_�_�_ �_u?�_�_�_o"o4o FoXojo|o�o�o�o�o �O�O�O	�O0BT fx������ ���_,�>�P�b�t� ��������Ώ���� ��o�o�o[����� ����ʟܟ� ��$� 6�H�Z��k������� Ưد���� �2�D� V�h�'���K���o�Կ ���
��.�@�R�d� vψϚϬϾ�Ͽ���� ��*�<�N�`�r߄� �ߨߺ�y��ߝ����� &�8�J�\�n���� �������������4� F�X�j�|��������� ��������-��Q ������� �,>Pb!� �������/ /(/:/L/^//A �/�/y�/�/ ??$? 6?H?Z?l?~?�?�?�? s�?�?�?O O2ODO VOhOzO�O�O�Oo/�/ �/�O_�/._@_R_d_ v_�_�_�_�_�_�_�_ o�?*o<oNo`oro�o �o�o�o�o�o�o�O _�O/Y_��� ������"�4� F�X�o|�������ď ֏�����0�B�T� %7I��mҟ� ����,�>�P�b�t� ������i�ί��� �(�:�L�^�p����� ����w���������$� 6�H�Z�l�~ϐϢϴ� �������ϻ� �2�D� V�h�zߌߞ߰����� ����
�ɿۿ�O�� v����������� ��*�<�N��_��� ������������ &8J\�}?� c�����"4 FXj|���� ���//0/B/T/ f/x/�/�/�/m�/� �/�?,?>?P?b?t? �?�?�?�?�?�?�?O �(O:OLO^OpO�O�O �O�O�O�O�O _�/!_ �/E_?	_~_�_�_�_ �_�_�_�_o o2oDo VoOzo�o�o�o�o�o �o�o
.@R_ s5_��mo��� ��*�<�N�`�r��� ����gȍޏ���� &�8�J�\�n������� c��џ���"�4� F�X�j�|�������į ֯������0�B�T� f�x���������ҿ� ������ٟ#�M��t� �ϘϪϼ�������� �(�:�L��p߂ߔ� �߸������� ��$� 6�H���+�=ϟ�a� ��������� �2�D� V�h�z�����]����� ����
.@Rd v���k�}������$FMR2_�GRP 1���� ��C4  B��	� ��9K6F�@ a@�6G��  �Fg�f�C�8R�y?��  ��66�X����875t���5���5`+=�yA�  /+�BH�w-%@S3	39%�5[/l-6@6!�/xl/�/�/�/ �/?�/&??J?5?G?��?k?�?��_CF/G �TK�?��? OO�9NO �
F0FA �K@�<RM_CHK?TYP  ��p$&� ROMa@�_MINg@������@�R XSS�B�3�� 7�O���C�O��O�5TP_DEF�_OW  ��|$WIRCOMf@�_�$GENOV_RD_DO�F��fE]TH��D dbU�dKT_ENB7_ �KPRAVC�:�G�@ �Y�O�_�?oyo&oI*� �QOU��NAIRI<�@��oGo�o�o,�o��C�p3�P�O:��B�+spL�i�O�PSMTኹY(�@
t�$HoOSTC�21�ε@�5 M5C��R{���  27.00�=1�  e�]� o�������K�ď֏���������	ano?nymous!�O�a�s����� �4��������D�!�3� E�W�i���������ï 柀�.���/�A�S� ��课�П����Ŀ ����+�r�O�a�s� �ϗϺ�������� �'�n��������ϓ� ڿ����������F�#� 5�G�Y�k���υ�� ��������B�T�f�C� z�g��ߋ�������� ����	-P����� u������(� :�<)p�M_q� �������/$ ZlI/[/m//�/� ���//�/D!?3? E?W?/?�?�?�?�? �/�?./OO/OAOSO �/�/�/�/�?�O?�O �O__+_r?O_a_s_ �_�_�O�?O�_�_o�o'o�t�qENT {1�hk P!�_.no  �p\o�o �o�o�o�o�o�o �o:_"�F�j �����%��I� �m�0���T�f�Ǐ�� 돮��ҏ3���,�i� X���P���t�՟��� ��
�/��S��w�:� ��^�������������ܯ=� �QUIC�C0J�&�!19�2.168.1.10c�X�1��v�8���\�2�ƿؿ9�!ROUTER:���!��a��P�CJOG��e�!�* ��0��U�C�AMPRT�϶�!1�����RTS����x� !Sof�tware Op�erator PanelU߇���7kNAME !Kj?!ROBO�����S_CFG 1��Ki ��Auto-sta�rted�DFTP�Oa�O�_���O ����������E_�.� @�R�u�c�	������� ����cN:�L�^�;r� ��R������� �%H�[m ���jO|O�O�O 4!/hE/W/i/{/�/ T�/�/�/�/�//�/ /?A?S?e?w?�?�� ��??�?</O+O=O OO?sO�O�O�O�O�? `O�O__'_9_K_�? �?�?�?�O�_�?�_�_ �_o#o�OGoYoko}o �o�_4o�o�o�o�o f_x_�_g�o��_ �����o��-� ?�Q�tu�������� Ϗ�(:L^`�2� �q�����������ݟ ���%�H�ʟ[�m� ���������� �ί 4�!�h�E�W�i�{��� T���ÿտ�
�Ϟ��/�A�S�e�w����_?ERR ��ڇ����PDUSIZ � �^6�����>��WRD ?�(����  ?guest����+�=�O�a���SC�D_GROUP [3�(� ,�"�wIFT��$PA��wOMP�� �޷_SH��ED�� �$C��COM��T�TP_AUTH �1��� <!iPendanm��x�#�+!KAR�EL:*x����KC������V�ISION SET��(����?�-�W�R���v������������������G�CTR/L ���a��
��FFF�9E3��FR�S:DEFAUL�T�FANU�C Web Server�
tdG� ���/� 2D�V��WR_CON�FIG ���������ID�L_CPU_PC�� �B���� ;BH�MIN���~�GNR_IO�������ȰHMI_EDIT ���
 ($/C/��2/ k/V/�/z/�/�/�/�/ �/?�/1??U?@?y? d?�?�?./�?�?�?�? OO?OQO<OuO`O�O �O�O�O�O�O�O__�;_�NPT_SI�M_DO�*N�STAL_SCR�N� �\UQTPMODNTOL�Wl[�RTYbX�qV\�K�ENB�W����OLNK 1�����o%o7oIo[o�moo�RMASTE���Y%OSLA�VE ��ϮeRAMCACHE�o��ROM�O_CFG�o�S�cUO'��b?CMT_OP�  "��5sYCL�ou� _ASG 1����
 �o��� ����"�4�F�X��j�|����kwrNUMj����
�bIP�o��gRTRY_CNx@uQ_UPD�Êa��� �bp�bA��n��M��аP}T{?��k ��._ ������ɟ۟퟈S�� �)�;�M�_�q� ��� ����˯ݯ�~��%� 7�I�[�m�������� ǿٿ�����!�3�E� W�i�{�
ϟϱ����� ���ψϚ�/�A�S�e� w߉�߭߿������� ��+�=�O�a�s�� �&���������� ��9�K�]�o�����"� �������������� GYk}��0� ����CU gy��,>�� �	//-/�Q/c/u/ �/�/�/:/�/�/�/? ?)?�/�/_?q?�?�? �?�?H?�?�?OO%O 7O�?[OmOO�O�O�O DOVO�O�O_!_3_E_ �Oi_{_�_�_�_�_R_ �_�_oo/oAo�_�_ wo�o�o�o�o�o`o�o +=O�os� ����\n�� '�9�K�]��������ාɏۏi�c�_ME�MBERS 2��:�  � $:� ����v���1���RCA_ACC 2���  � [~�v eL�Kl�6M@��  �!l�l��6L%Pl������$�����a�BUF001 �2�n�= ���u0  u0�ɪ��������T�$�"�"�("�U5"�D"�Q"�`"�Ul"�y"��"��"�U�"��"��"��"���"��"���������"��/��=���L��Z��i��v���y�  �[����������"�"�"�**"�7"�E"�R"�a��m"�z� $��Ȑ����'��3�B�N�[��j�w����J�����ߙ2� ��������� !��(�-�1�-�9�-� A�-�I�-�Q�-�Y�-� a�-�i�-�q�-�y�-� ��-�-�-�-� ��-©�-±�-¹�� ����ɠ��Ѡ��٠�� ��������������t� x�
�� ���!��(�-�1� -�9�-�A�-�I�-�Q� -�Y�-�j�h�-�q�� y�z������ ��¡�©�±�� ������ɰ�Ѱ� ٰ���ߙ3���� �����!�/�6� 1�?�6�A�O�6�Q�_� 6�a�o�6�q��6⁢ ��6③��6⡢��6� ����l�������Ѣ�� ������������� ��	����'�l�(� 7�6�9�G�6�I�W�6� Y�g�6�i�w��y��� ≲��♲��⩲ ��⹲���ɲ����ٲ����d�CFG ;2�n� 4��*l�l�<l�47]��HIS钜n�� �� 2025-11-3��l�   � # &f � ' "珪� � ��6X�`�hdl��pl�ʐx {��8 �l�;  ��   7 ����9 �9, ����7[}�Rq29 }	7v��������)� % �� �  -�RO  *� l��B��aN/`/r/�/�/ �/�/�/�/�/'/9/&? 8?J?\?n?�?�?�?�? �?�/?�?O"O4OFO XOjO|O�O�O�?�?�O �O�O__0_B_T_f_ x_�O�O�O�_�_�_�_ oo,o>oPo�O���[m
8 c� 8@���o�o�6d� ��b� �b� +  �X�  X� 6dT6c	,: J{�|!r0  Q!1 
 R)!r�� !r9K]���� �����:�a��2�a ,*q 1  \�_�_m���� ����Ǐُ�����_ X�E�W�i�{������� ß՟��0���/�A� S�e�w����������� ����+�=�O�a� s���������߿� ��'�9�K�]�oρ� J�Ѐo�o

eq� ��������� �� � ��� ��� eq� �Geq	$"��eqeq!� "n� Vpn�^p������� �� ��$�6���� �� Z� �־�п ������������ &�8�o��n������� ����������G�Y� FXj|���� ��1�0BT fx�����	 //,/>/P/b/t/��/�/�Ϙ�I_CF�G 2��� H�
Cycle �Time�Bu{sy�Idl�"^�min�+1�Up�&�R�ead�'Do�w8?�` 1�#C�ount�	Num �"����<��zb�qaPROG�"�������)�/softpar�t/genlin�k?curren�t=menupa�ge,1133,1�/OO/OAO3b5�leSDT_ISO_LC  ���p��/J23_DSP_ENBL�vK0~�@INC ��M|�ӄ@A   ?&p�=���<#�
<�A�I:�oJp�N`_���O<_�GOB�0�C�CF�1�FVQG_�GROUP 1�vvK	r<�P�C�٢_D_?���?�_��Q�_o.o@o�_ dovo�o�o��,_NY�G_IN_AUT�ODԫMPOSRE�^_pVKANJI_�MASK v�HqR�ELMON ��˔?��y_ox������.6r�3��7ĲC���u�o�DKCwL_L�`NUML���EYLOGGINGDЫ���Q�E�0�LANGUAGE� ��~���DEFAULT� ����LG�!���:2�?�W��80H  ���'~��  � 
���囊�GOUF ;���
��(UT13:\��  �-� ?�Q�h�u���������ϟ�����(g4�8�i�N_DISP ���O8�_�_��L�OCTOL����D�z`�A�A��GBO_OK ���d�1
�
�۠#���� �#�5�G�Y�i���3{�W�	��쉞QQJ�¿Կ1��_BU�FF 2�vK 	���25
�ڢVB�&�7 Coll�aborativ �=�OΗώϠϲ��� ������'��0�]�T��fߓߊߜ��DCS ��9�B�Ax����Rh�%�-�?�Q���I�O 2��� ���Q���� ����������*�<� N�b�r����������������&:e�E_R_ITMsNd�o ������� #5GYk}����������hS�EV�`�MdTYPsN�c/u/�/
-��aRST5���SC�RN_FL 2�
s��0����/??`1?C?U?g?�/TPK��sOR"��NGNA�M�D��~�N�UPS�_ACR� �4D�IGI�8+)U_�LOAD[PG �%�:%T_NO�VICEt?��MA?XUALRM2��a����E
ZB�1_�P�5�` ��y�Z@CY��˭�O+���ۡ��D|PP 2�˫ �Uf	R/_
_C_ ._g_y_\_�_�_�_�_ �_�_�_oo?oQo4o uo`o�o|o�o�o�o�o �o)M8qT f������� %��I�,�>��j��� ��Ǐُ�����!�� �W�B�{�f������� ՟����ܟ�/��S� >�w���l�����ѯ�� Ư��+��O�a�D����p���RHDBGDEF ��E�ѱO���_LDXDIS�A�0�;c�MEMO�_AP�0E ?�;
 ױ��3� E�W�i�{ύϟϱ�Z@�FRQ_CFG k��G۳A ���@��Ô�<��d%��� ������B��K{��*i�=/k� **:tҔ� g�y�ߔ��߱����� �����J�Es��J d�����,( H���[�����@�'� Q�v�]����������������*NPJI�SC 1��9Z� ������ܿ������	Zl_MST�R �#-,SC/D 1�"͠{ �������� //A/,/e/P/�/t/ �/�/�/�/�/?�/+? ?O?:?L?�?p?�?�? �?�?�?�?O'OOKO 6OoOZO�O~O�O�O�O �O�O_�O5_ _Y_D_ i_�_z_�_�_�_�_�_ �_o
ooUo@oyodo �o�o�o�o�o�o�o�?*cN�M�K���;љ$�MLTARM��u�N��r ���հ��İMETP�U��zr��CN�DSP_ADCO�L%�ٰ0�CMNT6F� 9�FNb�f�>7�FSTLI��x�4 �;ڎ�s�����9�POSCFz��q�PRPMe���STD�1�;; 4�#�
v��q v�����r�������� ̟ޟ ���V�8�J� ��n���¯��������9�SING_CH�K  ��$MODA���t�{�~~2�DEV 	��	MC:f�HS�IZE��zp�2�T�ASK %�%�$1234567�89 ӿ�0�TR�IG 1�; lĵ�2ϻ�!�bϻ�F��YP����H�1��EM_INF 1��N�`)AT&FV0E0g����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ��2��H6�^���R����A�߶�q�������� ��5������ ߏ�B߳�������� ���1�C�*�g��,� ��P�b�t������ R�?���u0�� ������������� M q���Z� ��/�%/��[/  2�/�/h�// �/�/�3?�/W?>?{? �?@/�?d/v/�/�/O �//OAOx?eO?�ODO��O�O�O�O_�NIT�ORÀG ?z� �  	EXESC1~s&R2,X3,XE4,X5,X��.V7,X8,X9~s'R�2�T +R�T7R�TCR�TOR�T [R�TgR�TsR�TR�TT�R�S2�X2�X2�XU2�X2�X2�X2�XU2�X2�X2h3�X�3�X37R2�R_G�RP_SV 1��� (�>���R>15����s?	zQ��*�V?R�a���_�D�B���cION_�DB<��@�zq W �2p�2p�Y��1t �zp�>w�/  �^p�Y��@�N   `rpa�>{ep�Y�-ud1�����8��PG_JOG ��ʏ�{
�2��:�o�=���?����0�B��~\�n��������0H�?��C�@�ŏ׏����rp�����qL�_NAME !�ĵ8��!De�fault Pe�rsonalit�y (from �FD)qp0�RMK_ENONLY��_�R2�a 1�L�XL�8�gpl d����ş ן�����1�C�U� g�y���������ӯ� ��	����
�<�N�`� r���������̿޿� :��)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+��<�Sew����������A;�yq  B�Bw��Pf��� ���/!/3/E/W/ i/{/�/�/�/���/ �/??/?A?S?e?w? �?�?�?�?�?�?�?�/ �/+O=OOOaOsO�O�O �O�O�O�O�O__'_`9_&O�S���x_�]�rdtS���_�]�_ �_�W�����S"oe_oXoa ��qogo yo�o�o�o�o�ouP�p("|����	upE Wi{~9pK�A\��8��s� A ��y�@h�Q�Q��"����Tk\$�� W ��P�PE�x?C�  �I�@o a�<o��p�������ߏ 
f�Q*�����0��P�Cr� � �3r �.� @D��  A�?�G�-�?x.I�.@I�A�����  ;�	l�Y�	 �X?  ������� �, ǀ �����uPK��o�����]K���K]�K	�.��w�r_	����@
�)�b�1������I�Y������T;fY�{{S���3�����I�>J���;Î?v߮>��=@�����E��RѯעZ����wp��u�� D�!�3��7pg  �  �9��͏W���	'� �� u�I� ��  ��u��:��È��È=�s�ͱ���@��@ǰ�3��\�3�E��&���N�pC�  'AY�&�Z�i�b�@f��i�n�C����I�Ch����b��r0����ڟ.�B�p����q���}ر�.Dz Ə<ߛ�`�K�pߖ���w������А 4P�����.z��d  ��Pؠ?�ff0�_��	�� 2p>��P���8.f�t�>L����U���(.��P ���٨�����É���{ x��;e�m����KZ;�=g;�4�<<����%�G��3����p�?fff?ذ?&�S���@=0e�?��q�+�rN�Z� ��I���G���7���(� ����!E0iT�����+��F �p���#��D�� w����� ��//=/(/a/L/ �/p/��/�p�6�/ Z#?�/ ?Y?k?}?� �?�?>?�?�?�?�?�?�1O�����KD�y^KC�O�OO�O����`�O�O�O�Oai���1J��}�DD1���.B�D��@�AmQa��9N�,ȴA;�^@���T@|j@�$�?�V�>��z�ý��=�#�
>\)?��
=�G�-]��{=���,���C+��B�p���P��6���C98R����?N@��(��5�-]G�p�G�sb�F�}�G��>.E�VD��Kn���I��� F�W�E���'E���D���;n���I���`E�G���cE�vmD���-_�oQ_�o�o �o �o$H3X ~i������ ���D�/�h�S��� w��������я
��� .��R�=�v�a�s��� ��П����ߟ��(� N�9�r�]��������� ޯɯۯ���8�#�\� G���k�������ڿſ ���"��F�1�C�|� gϠϋ��ϯ����������P(�Q34�] �����Q�	�9�O��53~�mm��a�ǀ5Q�߫�aғ�����ߵ1��� ����1��U�C�y�g�J�%P�P���!�/���'���
���.������4�;�t�_��� ������������ :%��/�/d�������� 7%[Im���027�  B��S@J@�CH#PzS@�0@ZO/1/C/U/g/y/�-�#��/�/0�/�/�/�3?�3�� @�3��0ĵ0�13��5
 ?f?x?�?�?�?�? �?�?�?OO,O>OPO��Z@1 ���ۯ��c/�$MR_CABLE 2ƕ� ��TT �����ڰO���O�)�@ ���C_���_O_u_ 7_I__�_�_�_�_�_ o�_�_oKoqo3oEo {o�o�o�o�o�o�o�o �oGm/�K!�"���O����ذp�$�6���*Y��** �COM }ȖI���0�* e.�%% �2345678901���� ��Ï��R� � !� �!�
���Mnot sent b���W��TE�STFECSAL?GR  eg�*!�d[�41�
k�������$pB����������� 9UD1�:\mainte�nances.xsmlğ�  C:��DEFAU�LT�,�BGRP {2�z�  ��"���%  �%!1�st clean�ing of c�ont. v�i�lation 56��ڧ�!0�����+B��*������+��"%��mec�h��cal ch�eck1�  �Bk�0u�|��ԯ�����Ϳ߿�@���rollerS�e�w�ū��m�ϑϣϵ��@�Basic �quarterl!y�*�<�ƪ,\�)�`;�M�_�q�8�MJ�,�ߓ "8��� ���ߕ �����+�=��C�g�ߋ�ʦ�߹��������@��Overhaul�ߔ��?� x� I�P����}���������� $n������ �)l�ASew��� ��� �+ =O�s���� ���/R�9/� (/��/�/�/�/�// �/�/N/#?r/G?Y?k? }?�?�/�???�?8? OO1OCOUO�?yO�? �?�O�?�O�O�O	__ jO?_�O�Ou_�O�_�_ �_�_�_0_oT_f_;o �__oqo�o�o�o�_�o o,oPo%7I[ m�o��o�o�� ��!�3��W��� �����ÏՏ�6��� �l����e�w����� ����џ�2��V�+� =�O�a�s������ ͯ����'�9��� ]�������⯷�ɿۿ ���N�#�r���YϨ� }Ϗϡϳ������8� J��n�C�U�g�yߋ� �ϯ������4�	�� -�?�Q��u������� ����������f�;� ������������� ���P���t�I[ m������ :!3EW�{ ��� ���/ /lA/��w/��/��/�/�/�/X*�"	 �X�/?.?@?�)B  a/o?m/o%w?�?�?}? �?�?OO�?�?OOaO sO1OCO�O�O�O�O�O __'_�O�O]_o_�_ ?_Q_�_�_�_�_�_�\� Џ!?�  @�! M?HoZo�lo�&4o�o�o�o�(�*�o** F�@ �Q�V�`o'�9�o]o�����/^&�o���� �/�A�S�e���#� ����я�����+� q�����7�������k� ͟ߟ��I�[���K� ]�o���C�����ɯ���o$�!�$MR�_HIST 2���U#�� 
 \�7"$ 23456789013�;��
�b2�90/����[� ��./����ǿٿF� X�j�!�3ρϲ���{� �ϟ�����B���f� x�/ߜ�S����߉��� ���,���P��t���=��$�SKCF�MAP  �UK&��b
�� �����ONREL  �$#������EXCFENB�q
����&�FNC-���JOGOVLI�M�d#�v���KE�Y�y���_P�AN������RU�Ni�y���SF?SPDTYPM�����SIGN��TO1MOTk�����_CE_GRP 1��U��+�0 �ow�#d��� ���&�6\ �7y�m�� �/�4/F/-/j/!/ t/�/�/�/{/�/�/�/�?�+��QZ_ED�IT
����TCO�M_CFG 1����0�}?�?�? 
>^1SI �N�!���?�?���?$O�����?XO78T_/ARC_*�X��T_MN_MOD�E
�U:_SP�L{O;�UAP_C�PL�O<�NOCH�ECK ?�� �� _#_5_ G_Y_k_}_�_�_�_�_��_�_�_oo��NO_WAIT_L	lS7> NTf1�����%��qa_ERR&H2�������?o�o�o�o��OGj�@O�cӦm| e#LOGOo��<���?���t��a~�b_PARAM�b����v_��w
�.�@� = n�]�o� w�Q�����������`Ϗ�)���w�[��m� �����ODRD�SP�C8�OFFSET_CARI0��OǖDISԟœS;_A�@ARK
T9�OPEN_FIL�E��1T6�0OPTION_IO�����K�M_PRG ;%��%$*�����'�WO��N�s�ǥ�� ���u����	� ����Ӧ������RG_DSBL'  ����jN����RIENTTO����C�����A� ��U�@IM_D�S���r��V��LCT �{mP2ڢȪ3̹��dҩ��_P�EX�@���RAT��G d8��̐UOP װ�:�����S�e�Kωϗ��$��r2G�L�X�LȚ�l 㰂�������'�9� K�]�o߁ߓߥ߷��� �������#�5�G���2��v������� ������e�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?�q1�~?�?�?�? �?�?�?�?O O2ODO^�yA�a�m? ~N��~O�O�P�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�O �Oo$o6oHoZolo~o �o�o�o�o�o�o�o  �_oVhz�� �����
��.��@�R�d�QOES��(����B�d�ӏ� ʏ��������Y�D�}�0��r������� ��ԟڟ���p���=�4M��q�	`����x����c�:�o��¯ԯ����A�C  �k�C�C�ڰe"ڰ���O���  ����-���)�C�  �t�k���g�����Կ ��ѿ
�5���_:�ĳ��OU���2��2�H��n��� � ^��\� @D�  &p�?�v�\�?:px��:qC4r�p�(�� � ;�	l��	 ��X � ������ ��, � �x������Hʪ�������H���Hw�zH����ϝ�8�B���B��  Xѐ�`�o�*��'3����t�>u����fC{ߍ��:pB\��
�Ѵ9:qK�t�� �����$���*��� D�P�^��b�g  �  �h������)�	'� �� ��I� ��  ��'�=��������t�@����!�b��^;bt�U�(�N��r� ' '��E�C�И�t�C�И��ߗ���jA��@�����%�B �� ��,���H:qDz�k�ߏz����������А 4P���:uz:���	�f��?�faf'�&8� ]��m�8:p��>!L�����$�(:p�P��	������:�� x�;e�m�"�KZ;�=g�;�4�<<�0��E/Tv��b����?fff?�?y&� )�@=0�%?��%_9��}! ��$�x��/v��/f'�� W,??P?;?t?_?�? �?�?�?�?�?O�?(O OLO�/�/�/EO�OAO �O�O�O�O_�O_H_ 3_l_W_�_{_�_�_1� �_A���eO+o�ORoo Oo�o�o�oK/�o�omo �o*'`+�,�zt���CL�H<��}?����X�
������u�����D1�/n�t�x�p�q��@I�h~�,ȴA;�^@���T@|j@�$�?�V�n��z�ý��=�#�
>\)?��
=�G�����{=��,���C+��B�p����6���C98R����?}p��(��5���G�p�G�sb�F�}�G��>.E�VD��KL����I��� F�W�E���'E���D���;L����I���`E�G���cE�vmD���\�՟��ҟ� ��/��S�>�w�b��� ����ѯ������� =�(�:�s�^������� ��߿ʿ�� �9�$� ]�Hρ�lϥϐϢ��� ������#��G�2�W� }�hߡߌ��߰����� ���
�C�.�g�R�� v��������	��� -��Q�<�u�`�r��� ����������'�M�(�34�]O!���8h~�%3~�m���ǀ5Q��������!���   `N�r��J	eP@"P��Q�_�/V/9/$/]/H)����c/j/�/�/�/ �/�/�/�/!??E?0? i?T?"&�_�_�?�?�8��?�?O�?OBO 0OfOTO�OxO�O�O�O��O2f?_  B���pyp$QCHR�z�p@�N_`_r_�_�_�_�]c�O�_�_0oo+o?�Bc�� @d4��QJc�D
 2o�o�o�o�o�o�o %7I[m���oa ������c/�$PARA�M_MENU ?� � � DEF�PULSE��	�WAITTMOU�T�{RCV� �SHELL_�WRK.$CUR�_STYL�p�"�OPT8Q8�PT�BM�G�C�R_DECSN�p����� ���������-�(� :�L�u�p��������q�SSREL_ID�  ��̕U�SE_PROG �%�z%���͓C�CR�pޒ��s1�_HOST !�z#!6�s�+�T�=����V�h���˯*�_�TIME�rޖF�~�pGDEBUGܐ��{͓GINP_F�LMSK��#�TR\2�#�PGAP� ���_b�CH1�"�TWYPE�|�P�� ������0�Y�T� f�xϡϜϮ������� ���1�,�>�P�y�t� �ߘ��߼�����	�� �(�Q�L�^�p��%�WORD ?	�{
 	PR��p#MAI��q"3SUd���TE��p#��	1���COL�n%��!���L�� �!��F�d�T�RACECTL �1� �q }�~ #�����_�DT Q�� ��z�D �� �^a����c`�������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I?�[?m??�  �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_ J_\_n_�_�_�_�_�_ �]��5oo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�.�oP�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/Dϒ/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D��V�h�z�����������$PGTRACE�LEN  �� � ������Ά_UP _�����������΁_CFoG ����*��
���*�:�D��O���O�  ��O��DEFSPD� ��������΀H_CONF�IG ����� ����dĔ�&݂ ��ǑP^�a�l㑹��΀IN�?TRL ��=��8^���PE��������*�ÑO��΀LID���	~T�LLB 1ⳙ_ ��BӐsB4��O� �𼧶��Q� <<7 ��?��� ����M�3�U���i� ��������ӿ��	�7�T�Ϣk�b�tϡπ诚��������S�G�RP 1爬����@A!���4�I���A �C�u�C�OCWjVF�/��Ȕ`a�zي�ÑÐ�t�0�ޯs���´�ӿ���B������������A�S�&�B3�4�_������j���������	� B�-���Q���M�������  Dz����.� ����&L7p[ ��������6!Zh)w�
V7.10be�ta1*�Ɛ@��*�@�) @ߺ+A Ē?���
?fff>�����B33�A�Q�0�B(���A���AK��h����//('/9/P�p*�W�ӑ��n/�/�%���R��fh���� *���P2�LR��/�/@�/�/�/H?�Ĕ�I�u�&:���?��x?��?A���P!\3 Bfu�B��?�5BH�3�[4��o��4�I�[45��/B\3x3Dx�?YO�?aOkO}O�<<�R@��O�C�O�O��O�O�DA�X�KNO?W_M  Z�%��X�SV 賚ڒ���_�_�_?��_�_�_o����W�M�+�鳛 ��	~@�3#���_��o�\A��
]bV4�@u��u��e��o�l,�X�MR+��JmT3?��W�1C{��OADBANFW�DL_V�ST+�1 k1����P4C� ��[��i/��� ��?�1�C���g�y� �������ӏ�*�	�@�`�?�Q�c��w2�|8Va�up�<ʟ����p3��Ɵ؟Ꟃw4 ��+�=��w5Z�l�~����w6����ѯ㯂�w7 ��$�6��w8`S�e�w����wMAmp�������OVL/D  ��yo���rPARNUM � �{+þ�?υqS[CH�� �
��pX���{s��UPDX��)ź��Ϧ�_CMPa_@`���p|P'yu~�ER_CHK���yqbb3��.��RSpp?Q_MO�m��_}ߥ�_REWS_G�p쩻
� e�����0�#�T�G�x� k�}��������������׳�������� �:�Y�^���Y�y��� ���Ӭ����������� ����R�6UZ��ӥ�u����V �1�FvpVa@k��p��THR_ICNRp��(byudoMASS Z)�MNGMON_�QUEUE �P�uyvup\!��N��UZ�NW��ENqD��߶EXE�����BE���O�PTIO��ۚP�ROGRAM %z%��~Ϙ?TASK_I��.OCFG �zx+�n/� DATACcm�+�0��up 2 �?�?/?A?S?]51  s?�?�?�?�?�6p1�?��?�?O"O,F�!IN+FOCc��-��bd lO~O�O�O�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_�_�_�/A@FD���, 	��!��K�_�!�)fN!fECNB��0m��Pf2Yo�khG�!2�0k �X,		d�=���·o���e�a$��pd��i�i�g_E?DIT ��/%�7����*SYS�TEM*upV9.�40107 cr7�/23/2021� A��Pw���PRGADJ_�p  h $X|[�p $Y�xZ�xW�xқtZқt?SPEED_�p�p�$NEXT_C�YCLE�p���q�FG�p ���pALGO_V� �pNYQ_F�REQ�WIN_�TYP�q)�SIuZ1�O�LAP�r�!�[��M+����qC?REATED�r��IFY�r@!NAM��p%h�_GJ�S�TATU��J�DE�BUG�rMAIL�TI����EVE<U��LAST������tELEM� �� $ENAB<�rN�EASI򁼁�AXIS�p$P�߄�����qROT�_RA" �rMAX� ��qE��LC�A�B
���C D_L9VՁ`�BAS��`��1�{���_� ��Y$x���RM� RB��;�DIS����X_cSPo�΁�� �u|�P� | 	�� 2 \�AN�� �;����8�Ӓ�� �0�PAYLO��3�V�_DOU�qS���p��tPREF� �( $GRID*�E
���R���9Y��rOTOƀ�q�  �p��!��p��k�OXY�� � $L��_�PO|�נVa�S�RV��)���DI?RECT_1� �U2(�3(�4(�5(��6(�7(�8��qFꔑA�� $V�ALu�GROU�P�������� !��@!��8�����RAN泲�⚁R��/���TOTaA��F��PW��I=!%�REGEN #�8�������/��фڶnTzЉ���#�_!S����8�(�V[�'�8��4���GRE��w����H��D�����V_]H��DAY3�V���S_Y�Œ;�SU�MMAR��2 �$CONFIG�_SEȃ���ʅ_�RUN�m�C�С�$�CMPR��P�D�EV���_�I��ZP�*��q��ENH�ANCE�	�
����1���INT���qM)b�q�2Kܖ���OVRo�PG�u�IX��;���OV�CT�����v�
 4� ����a˟��P�SLG"�� \ �;��?�1���qSƁϕc�U� ����Ò�4�U�q]�|Tp� (`�T-��rJ<�O� CK�OIL_MJ���VN�L+��TQn{�N5����C�ULȀD�V(�C6�P_�຀@�mMW�V1V�V1d�U2s�2d�3s�3d�4s�4d��'�	��������p	�IN	VGIB1qp1� 2!�pq/,3 3,4 4,�p?��;���A���N�������PL��TORr3�	���[�SAV���d�MC_F�OLD 	$CSL�����M,�1I��L� �pL��b��KEEP_H/NADD	!Ke��UCCOMc�`k��
�lOP����pl��lREM�k��΢����U��ekHPWv� KSBM��~ŠCOLLAB|��Ӱn��n�+�ITz�O��$NOL��FCALX� �DO�N�r���� �,��FL���$�SYNy,M�C�=����UP_DL�Y�qs"DELAh� ����Y(�AD���$TABTP_�R�#��QSKI�Pj% ����OaR� �E�� P_�� � �)���p7��%9 ��%9A�$:N�$:[�$:@h�$:u�$:��$:9�q��RA�� X������MB�NFGLIC]��0"�U!�<o���NO_H� ��\�< _SWITC�Hk�RA_PAR�AMG� �4�p��U��WJ��:C|ӣ�NGRLT� OO�U�����X�<A���T_Ja1F�rAP�S�WEIGH]�Jg4CH�aDOR��aD��OO��)�2�_FJװ���sA�AV��C��HOB.�.���J2��0�q$�EX��T$�'QIT��'Q�pG�'Q-�G  �RD�C�m" � ��<��
R]��
H���RGEA��4��U�FLG`g��H��sER	�SPC6R��rUM_'P��2T�H2No��@Q ?1 ���0�����  D ��وIi�2_P�2�5cS�ᰁ+�L10�_CI�Ad� �pk����UՖ�D��zaxT�p�Q (�;a��c��޲+�i�p��e��` P`�DESIGRb$�V�L1:i1Gf�c�g10�_DS��D�wp~
`FPOS11�q l�pr��x1C�/#AT�B��U
WusIND��}�mq�Cp�mq`B	�HOMQE�r��?t2GrM�_q���|�?t3Gr��� ��$�`!@s4GrG�Y�k��}����� `a�q5Grď֏�����
��6GrA�S�e�w�L���� �0Ar7Gr��П�����0�8Gr;�M�_�q���䕯0�S �q    �@sM��P���<K@��! T`M�L�M�IO��m�I��:2�OK _OPy���x »Q�cPOWE�" 7�x EQ��b � #s%Ȳ$wDSBo�GNA�b�� C�P2�<rS2;32S�$ �iP��9xc�ICE<@%�cPE`2� @IT���P�OPB7 1�FLOW�TRa@2���U$�CUN��`�AU�XT��2Ѷ�ERF�AC3İUU��   �CH��% t<_9�EЎA�$FREEFROMЦ�A�PX qЎUPD"YbA�PT.�pEEX0���Í!�FA%bҬ���RV�aG� & W ��E�" 1�AL�  �+�jc'���D�  2& ��S\PcP(
  �$7P�%�R�2� ���T�`AXU���DSP���@�W���:`$��RNP�%�@����=K��_MIR����f�MT��AP�`��P"�qD�QSYz�������QPG7�BR�KH���ƅ AXI�  ^��i����1 ����BSOC����N��DUMM�Y16�1$SV�DE��I�FSP_D_OVR79�2 D����OR��֠�N"`��F_����@O�V��SF�RUN���"F0�����UF�"@G�TOd�LCH|�"�%RECOV��9@�@W�`&�ӂH���:`_0�  @>�RTINVE��8A�OFS��CK�KbFWD������1B喻�TR�a�B �FAD� ��1= B1pBL� �6� A1L�V��Kb����#��@+<�AM:��0��j��_M@ ~�@h����T$X`x ��T$HBK���F��A������PPA �
��	������?DVC_DB�3@@pA�A"��X1`�X3`��Se@�`��0��Uꣳ�h�CABPP
R�S #��c�B�@���GUBCP	U�"��S�P�`R���11)ARŲ�!$HW_CGpl�11�� F&A1Ԡ@8p�_$UNITr�l >e ATTRIr@y"���CYC5B�CA���FLTR_2_FI������2b�P��CHK_��S�CT��F_e'F_o,�"�*FS�Jj"CHA�Q�'91Is�82RSD����1���_Tg�`� �i�EM�NPMf�T�&2 8p&2- �6D�IAGpERAIL�ACNTBMw�LOh@�Q��7��PS��b� � ��PRB)SZ`�`BC4&�]	��FUN5s��RIN�PZaߠ�07DFh�RAH@���`� �`C�@�`C�Q�CBOLCURuH�DA�K�!�H�HDAp�aA�H�C�ELD������Cd��jA�1�CTIB�Uu�8p$CE_gRIA�QJ�AF �P��>S�`DUT2b�0C��};OI0DF_LC�H����k�LMLF�aHRgDYO���RG�@�HZ0��ߠ�@�UMUGLSE�P�'3iB$J��J����FAN_ALM�d�bWRNeHAR�D��ƽ�P��k@2�aN�r�J�_}�A�UJ R+4�TO_SBR��~b�Іje �6?A�cMPINF´�{!�d�A�cRE�G�NV��ɣZ�D���NFLW%6r$M�@� ��f� �0� h'uCM4NF�!�ON	 e!e#�p(b*r3F�3	�	 ����q)5�$�3$Y�r��u�_Ѿ�p*$ �/�EaGE�����qAR�Єi���2�3�u�@<�A�XE��ROB��R�ED��WR��c�_���SY`��q� ?�SI�WRI���vE �STհ�ӭ d���Eg!���t8��^a�БB����9�3� O�TO�a����AR�Y��ǂ�1�����F�IE���$LIN]K�QGTH���T_������30���XYZ���!N*�OFF����J�ˀB��,Bl�0��e���m�FI� ���C@Iû�,B��_J $�F�����S`����3-!$1�w0���R2��C��,�DU���3�P�3TUR`XS.�Ձ�bXX�� ݗFL�d���pL�0�按34���� 1�)�K��M�5��5%B'��ORQ��6��fC㘴��0B�O ;�D�,������a�'OVE��rM���� �s2��s2��r1���0�0��0�g /�AN=!� 2�DQ�q���q�}R� *��6����s��V���SER��jA	�2E��H.�C��A���0���XE�2Ӈ�A��AAX ��F��A�N!�SŴ1 _��Q_Ɇ�^ʬ�^ʴ��^��0^ʙ�^ʷ�^�1 &�^ƒP[ɒPkɒP{� �P�ɒP�ɒP�ɒP�� �P�ɒP�����ɪ �R�>�DEBU=#$�8ADc�2����
�AB��7����V� <" 
��i�q��-!�� %��׆��׬��״��� �1�י��׷�JT��DR\�m�LAB��ݥ9 FGRO� ݒ=l� B_�1�u��� }��`����ޥ��qa��AND�����qa� �Eq��1�0�A@�� �NT$`��c�VEL�1��m��1`u���QP��m�NA[w�(�CN1� ��3����  �SERV9Ec�p+ $@@d@n��!��PO
�� _�0T !���򗱬p,  �$TRQ�b
�(� -DR2,�+"P�0_ . ql"@!�&ERR���"I� q���~TO	Q����L�p]�e��ʄ0G��%������RE�@ / �,��/I -��RA~� 2. d�r&�"  0�p�$&��2tPM��?�OC�A8 1 � pCOUNT��� �qFZN_wCFG2 4B �f�"T�:#��Ӝ�� )� `�s/3 ���M:0�R��qC@��/�:0�FA1P��?V�X������r���� �P�:b HELpe�4 5��B_wBAS�cRSR�f� @�S�!QY 1T�Y 2|*3|*4|*U5|*6|*7|*8��L!RO�����NL�q �AB���0Z �ACK��INT�_uUS`�Pta9_cPU�>b%ROU��PH@�h9#�u`w�9��TPFWD_KA1R��ar RE���PqP��A]@QUE�i@&��	�f�>`QaI`���9#�j3r��f�SCEME��6��PA�7STY4SO�0�DI'1�`���18�rQ�_TM�cMANR�QXF�END��$KEYSWIT�CHj31:A�4HE�	�BEATM�3PE�pLE��1��H�U~3F�42S?DD_O_HOMBPO:a60EF��PRr��(*�v�uC�@O�Qo ��OV_Mϒ��E�q�OCM���7��   8%HK�q5# D��g�Uj�2�M�p�4R��FOR]C�cWAR����8%OM�p 6 Q@�Ԣ�v`U|�P�pQ1�V'p�T3�V4��_& �S#O�0�L�R7��hUNLiOE0hdEDVa�  �p�@d8 <�pAQ9�l1MSU�PG�UaCALC__PLANcc1���AYS1�1���@�9O � X`��P  �q;a�թ�w��2��j�M$P�㣒�fyt$��rSC�M�pm�q @���aq��0�tYzZzEU�Q�b�� �T!�Hr�pPv�N�PX_ASf: �0g ADD���$SIZ%a$V�A��MULTI�P�"ns�PA�Q?; � $T9opH�B���rS��j!C~ ��vFRIF�2S��0�YT�pNF[DODBUX�B��u&�!�F��CMtA�Е����������� �S|Z ��< � �pƛTEg�����$SKGL��T��X�&{𷃥㰀��STMT<e�ЃPSEG�2���BW���SHOW�؅�1BAN�`TP�O���gᣥ������� V�_G�= ��$PC���O�kFB�QP\�SP�01A&0^�, VDG���>� �cA00�����P���P��P�P���P��5��6��U7��8��9��A�� b`���P��w᧖��!F����h���1��v�Th�י1�1�1��U1�1�1%�12�U1?�1L�1Y�1f�U2��2��2��2ʙU2י2�2�2��U2�2�2%�22�U2?�2L�2Y�2f�U3��3��3��3ʙ3י3�3���Ȫ�3�3%�32�3�߹3L�3Y�3f�4���4��4��4ʙ4�י4�4�4��4��4�4%�42�4�߹4L�4Y�4f�5���5��5��5ʙ5�י5�5�5��5��5�5%�52�5�߹5L�5Y�5f�6���6��6��6ʙ6�י6��6�6��6��6(�6%�62�6�߹6L�6Y�6f�7���7��7��7ʙ7�י7��7�7��7��7(�7%�72�7*߹7L�7Y�7f���V�`_UPD��?s �c 
]�V���@ x �$TOR�1T�  ��cOP �, ZQ_7RE^��� J���SsC�A��_�U�p��YSLO>A"A � �u$� v��w�@���@��bVALUv10�6�zF�ID_L[C�:HI5I�R$F�ILE_X3eu4u$�CA�SAV���B hM �E_B�LCK�3�ȁ�D_CPU��p��p�5hz�`Y��R3R� C � PaW��� 	�!LAށ�SR�#.!'$RUN�`G@%$D!'$@�@G%e!$e!'%HR0�3$� '$�QT2Pa_�LI�RD  �� G_O�2�0Po_EDI�R  � 7SPD�#E�"i�0ȁ�p	���DC�S9@G)F �? 
$JPC71q��� S:C;C9o$MDL7$5Pf>9TC�`@7UF�@r?8S� ?8COBu ��@
�"|�L�G�P�;;� 9:;�, 
�TABU�I_�!L�HGb�% �FB3G$��3A�sR�LLB_AVAI�B�3�!I $� SEL� NẼ�@RG_rD N��Ta �4{SC�PJ �1�/AB�PT�R=C_9M]`L�K \M f&/QL_��FMj��P�Gi�U9R�6��P+S_�P\� �p�E}E7B�TBC2�e�L ���``�`b$�!FT�P'T�`TDCg�� BPLp��sNU;WTH��qhhTgtWR�2$�pERVE.S�T;S�T�w�R_ACkP ?MX -$�Q�`@.S�T;S�PU@�`ICn�`LOW�GF1�QR2g�`��p�S�ERTIA�d^0i�P�PEkDEUe�LoACEMzCC#c�V�BrpTf�edg�a�TCV�l�adgTRQ�l�e�j|�Scu��e�dcu�J7_ 4JH!��Se@qde�Q�2�0���1�PRcuPJKlvVK<�~qcQ~q�w�spJ0��q�sJJv�sJJ�sAAL�s@�p�s�p�v���r5sS�`N1�l�p�k�`5d�XA_́�0QCF�BN `M GRO�U ��bh�NPC�0sD�REQUIR�R� EBU�C�Q�6=g0 2Mz��P�d�QSGUO�@^�)APPR0C7@֍ 
$� N��CL	O� ǉS^U܉Se�0�BC�@A�"P 䂽 M]P�`�`sR�_MGa!�C���+���0�@,�BRK*�N�OLD*�SHOR�TMO�!m�Z��JWA�SP�tp`�sp`�s�p`�sp`�sp`�A��7§�8sQ�!�QTQG� m��R.Q�<cQ�PATH�*�@ �*��X&���P�NT|@A�"p��� �IN�RUC4`a��-C�`UM��Y
`�)p��>�Q��cP����p��PAYLOA�h�J2L& R_Am@�L ������+�R_F2LSHR�T/�LO���0�8��>���ACRL0z��p�y�ޤsRH5b�$H+���FLEX꺃 �JVR P ��_._�_�_9A���US :�_�Vd` 0�G��_tQd`�_�_lF1G��ũ�o0oBoTofoxo��E�o�o�o �o�o�o�o ���� wz3lt����3EW$F�^zT!��X�'q ju��uu~�W؁� ��p�u�u�u�u������!BJ(�T ��P5�G�Y�' A1T��l�pEL0�_Bԕ�s�J�Sz�JENW�CTR7B`NA���d�HAND_VEB����TUO@�`+�`TSW��T�A�V� $$M��e G��AV�Qs�De�oA@A��@�	$�A5�G�AU�Ad�� 6�T�G�DU�Dd�PD�G/ -STI�5V�5Ng�DYF ��+� x����P&�G�&�A�@�lw�o�Q�k�P�� ����ʕӕܕ��"�JUW 7 ��� ��3%�?!AS�YMT��m�T�Vp�o�A�t�_SH� ~������$����Ưد�J񬢐�#39\"���_VI��`8|�q0V_UNIrS�4��.�Jmu�2��2 A��4X��4�6a�pt� ������&E_������RE��CH( X� ̱���T-Oc�PP�VsSvD�US�RU�P�����z@�D�A}@_5�U��P�EyAa��RPROG�_NA��$�$�LAST���CA�Ns�ISz@XYZ_SPu�DW]R@Ͱb,VSV@�E1QENc���DCUR�H ���H7R_T��YtQ"9S�d��O�TuP?�Z ��I�!A�D���Q���#�S�������3�vP [o � MEѡO��R#B�!T�PP�T0F@1�a�� ̰� h1a%iT0�� $DUMM�Y1��$PS_6��RF��  1�lf�i@FLA*�YP��bc$GLB_TI �U�e`ձ:�wLIF(!\�����g`OW�P��eV�OL#qb �a_2��[d2�[`����b؛P�cZ`TC��$�BAUDv��cST���B�2g`ARIT�Y0sD_WAItAeIyCJ2�OU6��ZqyyTLANS��`�{S�SZc��BUF_�r�fиx�P�yyCHK_�@CE�S��� JO`E�aA�x�bUBYT�����r�.�.�@ ��aA��M�������Q] Xʰ�����ST����SBR�@M21_@��T?$SV_ER�b�����CL�`��A1�Ol�BpPGLh0EW(!�^ 4 $a�$Uq$�q$W �9�A�@R��І�Uم_ "��Dw$GI��}$ف ^	Ӄ�(!�` L�.��"}$�F�"E6�NEAR���B$F}��T|QL�& �J�@�R� a7�$JOINTa�)�х�MSET(!b  "+�Ec�2�^�Se�:��J�_�(!c�  ھ�U�?���LOCK_FO@� �PoBGLV��GL'��TE�@XM���EMP����K��b��$U�؂a�2_���q�`<� �q��^��CE/�?��� �$KARb�M�ST�PDRA܀����VcECX�����IUq��av�HE�TOOiL���V��REǠ'IS3��6��A�CH̐m b^QON$e[d3���IdB�`�@$RAIL_B�OXEa���RO�B�@D�?���HOWWAR0Aa�i`-�ROLMtb��$�*����T��`����O_F�U�!��HTML�58QS�� �$ӂ�(!d���P�@��(!e�������� �oQր}p(!f t��m�^a��t��B�+PO��AIPE�N���O����q��>�AORDED�m ��z�XT`��A),� oQP�O�P go D �`OB� ����ǯ�Uc�`��� ��SYS��ADR���pP`U@^  hs ,"��f$A���E��E�QPVW�VA�Qi � 1�@ق�UPR�B��$EDI�Ad�V/SHWRU�z���cIS�Uq�pND�Px7���G�HEAD�!h @���!i�KEUq�O`CP)P��JMP���L�U:�RACEV�Tj���IL�5S��C��NE���TICK!M�KQ9���HNr�Gk @���HWC��qPHVF�i@STYeB+�LO�a���[�C�el3�
�@�F%$A���D=��S�!$@�1�p a�e�q�ePv �HVSQU��#LO<�b_1TERC`!zO@S?�m 5����R�m@3���ܡ�O`	c IZ�d�A�e�ha�qtb}�hA}pP�~r��_DO�B�Xr�pSSQ�SAXI�qB��v�bS�U�@TL�<��REQ_ܠ��CET���`�CY%���FY'��Af\!�\d9x�P ЂS=R$$nl-�w ������c
�uV
Qh(�A���dC`�A��	�Y��D��p�E"�		CC�C��/�/�/�	4F�SSC�` 7o h5�DSmడf[`SP�@�AT� �
R��L��XbAD�DR�s$Hp� IyF�Ch�_2CH����pO����- �TU�k�Ir p��CQUCp�QV��I�RAq�4���c��
K��
��V*���Pr 	\z�D����|,K� P�"CN��*CƮ���!�TXSCRE�E��s�Pp@�IN!A˃<�4�D�a����`t Tᫀ�b ����O Y6���º�U4h�RR�������R1��TC�UE��u ��j �qz`Ś��RS	ML��U����V�1tPS_��6\��1�9�G\���C��2@4 c2��0Ov�R���&F�AMTN_F�L*�`Q��W���_�BBL_/�WB`N�Pw ����BO ��BLE"�Cg�R"ޙDRIGHtRD<��!CKGRB`�E�T���G�AWIDT�Hs���RB��a�r7�UI��EYհRx d�ʰ�����`=y�BACK��tb4>U���PFO��QW�LAB�?(�PI<��$URm�~P�F�P�PHy1 y� 8 $�PT_��,"�R�PRUp�s�5�da���QO%!t�z�V�ȇ�pU�@�SR ���LUM�S�� GERVJ�рPP���T{ � " G�E�Rh� �¯�LP$AeE��)^g��lh�lh�ki5ik6ik7ikpP`�Z�x�����$u1��p�Q wzQUSRلO| <z��PU2��a#2�FOO 2�PR�I*m9�[�@pTR�IPK�m�UN[DO��})���0Yp��y�����h�����p ~�Rp�qG ��T���-!�rOS2��vR��2�s�CA�����r`�$;Ai�UIaCA���p�3Ib_�sOFFA�*D@���Ob�r�a5�L�t��GU���Ps������+QS�UB`� ��E_�EXE��VeуsW]O� �#��wF��WAl�p΁fP=
 V_DB��N�2SRT�pO�V☖����3OR/�5�RAU@6�TK���y__���� |j ��OWNj�34$GSRC�0`���DA�<��_MPFI����ESP��T�$0��c��g�n�z�E!G� `%�ۂ34J�n��COP��$`��p_���/�+�6����CT�Cہ�ہ��_��DCS��P�w�4�COMp�@�;��O`�=���K�^�/�VUT�q'���Y٤Z��2���@p�w#�SB����2�\0˰_���M��%!]�DIC�#��AY�3G�PEeE�@T�QS�VR1�D��eQL�� a��P �D ��f�z��f�> ����6�QA�t�b# ��L2SHADO�W��#ʱ_UNS3CAd�׳OWD�˰�DGDE#LEG�AC)�q'	�VC�\ C���  v����だm�RF07����7d`C2`7�DRKIVo���ϠC�A�]�(�` ���MY_UBY�d?Ĳ��s�個1��$0�����_hఆ���L��BM�A�$�DEY	�E�Xp@C�/�MU��X��,��0US����;p_R"1�0p#�2�}GPACIN*���RG��c�y�:�y�0�sy�C/�RE�R"!��q�y�D@� )L !�G�P�"��$Tp�R�pD@�&P�P�x1Q��	.���RE6��SWq�_Ar�u@I+�{�Oq�AA/��3�hEZ�U����� �p�HK���PJ��_/�Q0{�EAN��ۀ2�2�X���MRCVCA� �:`ORG��Q�dR�	��L�����REF oG�����!�+`	� p��������<���q�_����r��� S��`C��Ú�1�@D� ���!��#q��ơ�OU����?� 3��Վ2�n 0� 1�*p���l�0 UL�@��3CO�0)��� NT�[��Z�Qf�af% L飏���Q��a�VIAnچ� ��@HD7 �6P$JO�`oB�$Z_UPo�>�2Z_LOW���$�QiBn��1$EP�s�y�� 1!�f � 1¦4�� 5�PA�A� �CACH&�LO�w�ВaB�*��Cn�I#F^��qTm����$HO2�B32{��Uÿ2O�@ ���Ro��=a��Ɛ�VP��ՠA"_SI	Z&�K$Z$�F(�G'����CMPk*FAIjo�G��AD�)�/�MRE���"P'G�P�0е�9�ASY�NBUFǧRTD��%�$P!�COLE_'2D_4�5W�sw��~�UӍQO��%EwCCU��VEM��xv]2�VIRC�!5�#�2�!_>�*&�p�Wp��AG	9R�X#YZ@�3�W���8���4+Qz0T"��I�M�16�2`�GR�ABB�q��;�LE�RD�C ;�F_D��F�f50MH�PER�R [����JR�LAS�@��[_GEb� �H൑~23�ET����"���b¨�I�D�ҙ6m�BG�_LEVnQ{�PK�|Л6\q��GI�@N\P4�[�P��!gI�dr�S� �NRTZLʁc�Ų��#ah��c"!D�qDE�@���Xа�X���(�2��d��pzZ����d�c���D4q��W�2pT��U&�� -$�ITPr9p[Q8��ՓV�VSF$�d��  fp/�f�UmR��SMZu�dr���ADJ`C�� Z�DVf� D�XA�L� � 4 PER�IKB$MSG_Q3$Q!o%Y��p'��dr:g�qQ�^ �XVR\t��B�pT_\��R��ZABC"����Sr����
 Qp�`AC�TVS' � �� $|u�0�cCgTIV�Q!IOu�s&D�IT�x�D�Vϐ
x�P��4�!���pPS����� �#��!���q!L�STD�!�  �_ST�n��aq�;CHx�� L-�@���u�Ɛ*���P G�NA#�C�!q�_�FUN��   o�ZIPu��HR��$L���{p�_ZMPCF"��`b�ƀ�rX�ف��LNK���
	Ł�0#��� $ !��ބCWMCMk�C8�C"�����P{q $J8�2�D6!>�O� H���T���2�����M�怗UX�1݅UXE 1Ѡ��1C���Y�����p����˗7�FTFG�>������Z��A�s@�j�����Y}D'@ � 8n��R� Uӱ$HEgIGHd�:h?(! �'v� ����� � Gd��qp$�B% � E��SHIYF��hRVn�F�`�HpC� 3�(�8�H`O�ѡ�C��+%D,	�"�CE�pV�1�����PHERs� �� ,! M�c�u����$POWERFOL  �p|�����|�p�RG�`��������_�A�  ��?�p����pd��NSb �����?�  Bz|� �l�  <@�|��%���˃���8�ŵ�� 2ӷ��� 	H��l&����>���A� |��t$���*��/�� **:@���p�ϥ��͘���F������ɘ�� |�����5������� %ߟ�I�[߉�ߑ�� ����������w�!�3� a�W�i��������� ��O����9�/�A��� e�w�������'���� �=O}s �������k 'UK]��� ���C/��-/#/ 5/�/Y/k/�/�/�/? �/�/?�/?�?1?C? q?g?y?�?�?�?�?�? �?_O	OOIO?OQO�� 	 �O�O�O_ �E��3_���O`_�O�_��_÷PREF �Ӻ�p�p
��I?ORITY ��|�d���p����pSPL`z����WUT�VqÈ�gODU~����Y�_?�OG��Gx���R��,fHIBqO�y�|kTOENT �1��yP(!A�F_b�`�o�g!�tcp�o}!�ud�o)~!�icm�0bXY�̳�k �|�)�� �����p� ���u����� �N�5�r�Y��������̏�����*/c̳�ӹ���E�W�|�>�+k��F��/��4����|��,�7�A��_,  ��P�����%�|�'���Z@��h�z�����|���ENHANCE S	#�7�A9�d��<���  �,f�T�
�_�S����POSRTe�rb�@�U���_CARTR�EP�Pr|brSKS�TAg�kSLGS6�`�k����@�Unothing������Ϳ>��P�b�To��TEMPG ?isϨE/��_a_seibanm_��i_�����0� �T�?�x�cߜ߇ߙ� �߽�������>�)� N�t�_������� ������:�%�^�I� ��m�����������  ��$H3lWi ������� D/hS�w���uϪ�VERS�I�P=g  disable���SAVE �?j	2670H�705��k/!`�m//*�/ 	�(H%b�O�+�/�Se? 6?H?Z?l?z:%<�/�?4�*'_j` 1
�kX �0ubuE�?xOqG�PURGE��1Bp`�ncqWF<@�a�TӒ*fW�`]Daa��WRUP_DELAY z�f�B_HOT %?e�'b��OnER_NORMAL�HGb�O%_�GSEMI_*_i_��QQSKIP�3.��3x��_��_�_ �_�]?eo+goKo]o oo5o�o�o�o�o�o�o �o�o5GYi �}������ �1�C�U��y�g��� ������я����-��?�7%�$RACF�G �[ќ�3��]�_PARAMr�Q3y��S @И�@`�G�42Cj۠��2��CbFzB�B]�BTIF����J]�CVTMOUړ����]�DC�R�3�Y ���Q@�|1B��Q�B��@���(?ϩ�=L�����Z��i���i��1�h�@����G��x�_����;e�m����KZ;�=g;�4�<<���pf@����� � 5�G�Y�k�}��������ſ׿���xURDI�O_TYPE  ��V�5��EDPR�OT_a�&Y>��4BHbCEސ�SǆQ2c� ��B�ꐪϸ���� �����&�ݹ�W�V_ ~�o����߱����� ����A�O�m�r��� 9����������� ���=�_�d����� ������������' I�Nm���� �����#EJ i+k���� ��//4/F//g/ /�/y/�/�/�/�/�/ 	?+/0?O/?c?Q?�? u?�?�?�?�?�??;?�,O��S�INT 2��I���l�G;�� jO|K��鯤O�f�0 �O�K�?�O�? ___N_<_r_X_�_ �_�_�_�_�_�_�_&o oJo8ono�ofo�o�o �o�o�o�o�o"F 4j|b����������B�O�E�FPOS1 1~"�  xO ��o×O����ݏ鈃� ��Ϗ0��T��x�� ��7���ҟm������ ��>�P����7����� ��W��{�����:� կ^����������S� e��� ��$Ͽ�H�� l��iϢ�=���a��� ��� ߻����h�S� ��'߰�K���o���
� ��.���R���v��#� 5�o���������� <���9�r����1��� U�����������8# \����?�� u��"�FX� ?���_�� /�	/B/�f//�/ %/�/�/[/m/�/?�/ ,?�/P?�/t??q?�? E?�?i?�?�?O(O�? �?OpO[O�O/O�OSO �OwO�O_�O6_�OZ_ �O~_�_+_=_w_�_�_ �_�_ o�_Do�_Aozo<cf�2 1r�o .oho�o�o
o.�o R�oO�#�G� k�����N�9� r����1���U����� �����8�ӏ\���	� �U�����ڟu����� "����X��|���� ;�į_�q������	� B�ݯf����%����� [���ϣ�,�ǿٿ �%φ�qϪ�E���i� �ύ���(���L���p� ߔ�/�A�Sߍ����� ��6���Z���W�� +��O���s����� ����V�A�z����9� ��]���������@ ��d��#]�� �}�*�'` ���C�gy ��&//J/�n/	/ �/-/�/�/c/�/�/? �/4?�/�/�/-?�?y? �?M?�?q?�?�?�?0O �?TO�?xOO�O�o�d3 1�oIO[O�O _�O7_=O[_�O__ |_�_P_�_t_�_�_!o �_�_�_o{ofo�o:o �o^o�o�o�o�oA �oe �$6H� ����+��O�� L��� ���D�͏h�� �������K�6�o�
� ��.���R���퟈�� ��5�ПY�����R� ����ׯr�������� �U��y����8��� \�n�������?�ڿ c�����"τϽ�X��� |�ߠ�)�������"� ��nߧ�B���f��ߊ� ��%���I���m��� ,�>�P��������� 3���W���T���(��� L���p����������� S>w�6�Z ����=�a � Z���z /�'/�$/]/��/�/�/@/�/�O�D4 1�Ov/�/�/@?+? d?j/�?#?�?G?�?�? }?O�?*O�?NO�?�? OGO�O�O�OgO�O�O _�O_J_�On_	_�_ -_�_Q_c_u_�_o�_ 4o�_Xo�_|ooyo�o Mo�oqo�o�o�o�o �oxc�7�[ ����>��b� ���!�3�E����ˏ ���(�ÏL��I��� ���A�ʟe���� ���H�3�l����+� ��O���ꯅ����2� ͯV����O����� Կo�����Ϸ��R� �v�Ϛ�5Ͼ�Y�k� }Ϸ���<���`��� ��߁ߺ�U���y�� ��&���������k� ��?���c������"� ��F���j����)�;� M���������0�� T��Q�%�I��m��/�$5 1 �/���mX�� �P�t�/�3/ �W/�{//(/:/t/ �/�/�/�/?�/A?�/ >?w??�?6?�?Z?�? ~?�?�?�?=O(OaO�? �O O�ODO�O�OzO_ �O'_�OK_�O�O
_D_ �_�_�_d_�_�_o�_ oGo�_koo�o*o�o No`oro�o�o1�o U�oyv�J� n������� u�`���4���X��|� ޏ���;�֏_����� �0�B�|�ݟȟ��� %���I��F����� >�ǯb�믆������ E�0�i����(���L� ��翂�Ϧ�/�ʿS� � ��LϭϘ���l� �ϐ�ߴ��O���s� ߗ�2߻�V�h�zߴ� � �9���]��߁�� ~��R���v����#�<	6 1&�� �������������}� ��<��`��� �CUg�� &�J�n	k� ?�c��/�� �	/j/U/�/)/�/M/ �/q/�/?�/0?�/T? �/x??%?7?q?�?�? �?�?O�?>O�?;OtO O�O3O�OWO�O{O�O �O�O:_%_^_�O�__ �_A_�_�_w_ o�_$o �_Ho�_�_oAo�o�o �oao�o�o�oD �oh�'�K] o�
��.��R�� v��s���G�Џk�� �����ŏ׏�r�]� ��1���U�ޟy�۟� ��8�ӟ\������-� ?�y�گů����"��� F��C�|����;�Ŀ _�迃������B�-� f�ϊ�%Ϯ�Iϫ��� �ߣ�,���P�6�H�7 1S����I� �߲�������3��� 0�i���(��L��� p�����/��S��� w����6�����l��� ����=������6 ���V�z�  9�]��� @Rd���#/� G/�k//h/�/</�/ `/�/�/?�/�/�/? g?R?�?&?�?J?�?n? �?	O�?-O�?QO�?uO O"O4OnO�O�O�O�O _�O;_�O8_q__�_ 0_�_T_�_x_�_�_�_ 7o"o[o�_oo�o>o �o�oto�o�o!�oE �o�o>���^ �����A��e�  ���$���H�Z�l��� ��+�ƏO��s�� p���D�͟h�񟌟� ��ԟ�o�Z���.� ��R�ۯv�د���5��ЯY���}�c�u�8 1��*�<�v���߿ ��<�׿`���]ϖ� 1Ϻ�U���y�ߝϯ� ����\�G߀�ߤ�?� ��c����ߙ�"��F� ��j���)�c���� ������0���-�f� ���%���I���m�� ����,P��t �3��i�� �:���3� �S�w /��6/ �Z/�~//�/=/O/ a/�/�/�/ ?�/D?�/ h??e?�?9?�?]?�? �?
O�?�?�?OdOOO �O#O�OGO�OkO�O_ �O*_�ON_�Or___ 1_k_�_�_�_�_o�_ 8o�_5ono	o�o-o�o Qo�ouo�o�o�o4 X�o|�;�� q����B��� �;�������[��� ����>�ُb������!�������MASKW 1 ��������ΗXNO  �ݟ���MOTE � ���S�_CFG' !Z���N������PL_RANG�V�N������OWE/R "��Ϡ���SM_DRYPRoG %���%W���եTART �#Ǯ�UME_P�RO���q���_E�XEC_ENB � ����GSPD�J�������TD�B����RMп��I�A_OPTION��������N�GVERS���`�řI_AIoRPUR�� R��+���ÛMT_֐T� X���ΐOBOT_ISOLC�����������NA�ME8��H�ĚOB?_CATEG�ϣ�,��S�[�.�OR�D_NUM ?�Ǩ��H705  N��ߨ����ΐPC_TIMoEOUT�� xΐoS232s�1$���� LTE�ACH PEND�AN��o���)���V�T�Mai�ntenance_ ConsN�&��M�"B�P�No Use6�r�8���������̒��NPO�$��Ҏ�"���C�H_LM�Q���	�a�,�!UD1�:��.�RՐVAI�Lw��粥*�S�R  t� ����5�R_INTVAL���� ����V_DATA_?GRP 2'���_� D��P�� �����	���� ��B0RT f������/ �/>/,/b/P/�/t/ �/�/�/�/�/?�/(? ?L?:?p?^?�?�?�? �?�?�?�?O O"O$O 6OlOZO�O~O�O�O�O �O�O_�O2_ _V_D_ z_h_�_�_�_�_�_�_ �_o
o@o.oPovodo��o��$SAF_DO_PULSW��[�S���i�SCANd�������SCà�(2�3}���S�S�
������q�q�
qN� �L^p ���5��� �X�$��+��r2M�qqdY�P�`�rJ�	t/� @��@������ʋ|��� r �ք��_ @N�T ��'�9�K�X�?T D��X��� ������ɟ۟���� #�5�G�Y�k�}�����x��䅎������Ǧ  "�;G�oR� ���p�"�
�u��D�i���q$q�  � ���uq%�\� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z����珈������ ������g�;�D�V� h�z���������������(�Ӣ0�r�i�y� ��$�7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/?r�+?=?O?a? s?�?�?�?�?�?8��? OO'O9OKO]OoO�O ��$�r�O�O�O�O 	__-_?_Q_c_u_�_ �Y�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4@FXj|�c�路 g�������0� B�T�f�x���������ҏ������:�.Ҧ��y�3�	��	123456�78��h!B!�� \��p0����Ο�� ���(�:�@��c� u���������ϯ�� ��)�;�M�_�q��� ��R���ɿۿ���� #�5�G�Y�k�}Ϗϡ� �����ϖ�����1� C�U�g�yߋߝ߯��� ������	��-���Q� c�u��������� ����)�;�M�_�q� ��B���������� %7I[m� �������! 3EWi{��� ����////� S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?D/�?�?�?�?�? OO'O9OKO]OoO�O@�O�O�O�O�O*��� �O	_�E�?5_G_Y_�yCz  A��z_   ��x2�r� }��)�
�W�  	�*�2�O�_�_ o$o"l�#\��_ho zo�o�o�o�o�o�o�o 
.@Rdv� ���Mo���� *�<�N�`�r������� ��̏ޏ����&�8��J��X #P$P�Q�R<�u� k��Q  ������S�P����Q�Qt  ЌPÙ۟�P(� `�,b����]�PFl��$SCR_GRP� 1*3+�34� � ��,a �U	 v��~������d���%����ɯ���h]���P�D1� D�7n��3��Fl
C�RX-10iA/�L 234567W890�Pd� r���Pd�L ��,aC
1o��������[ ¶~�+fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@�R�d�t�?��H�~����m��ϴ����������,a��1���U�T[�G�imXhuP,��?B�  BƠߞ��Ԛ�A�P��  @�1`�՚�@����� ?���H��������F@ F�` A�I�@�m�X��|�� �������������`:�%�7�I�[�B�i� ��������������� -Q<u`��@En�ٯ���W�P�"+f@_�5��1`4b���x����ͣ�O�,dA����$���Fa�,a �#!"/4/E-!�Z(f/x/G/ (�P�!(� �/�/�/��/�/?#9b�����S7س�M�ECLV�L  ,a���ݲ�Q@f1L_D?EFAULTn4b1_�1`�3?HOTSTR�=���2MIPOWER�Fm0pU�5�4W7FDO�6 �5L��ERVENT 1�+u1u1�3 L!�DUM_EIP�#?5H�j!AF�_INE�0SO,d!'FT)O�NIO�O9!���O ��O�O�!RPC_MAIN�O�H��O>_S'VIS_�I�-_�_?!OPCUf�_�Wy_�_!TMP�PPU�_<Id�_�"o!
PMON_�PROXY#o?Fe ono�R<o8Mf]o�o�!RDM_SR�V�o<Ig�o!�R��"=Hh�oR!%
PM�o9LiA��!RLSYNC̟�y8��!gROS(O��4��6�!
CE�PMT'COM7�?Fk%���{!	K�CONS���>Glq�Ώ!K�WOASRC�o?Fm��v�!K�USB��=Hn	�f�!STM�0��;JoU����O�֟�c����CICE�_KL ?%K� (%SVCPGRG1��G�1�2G�DL�6�3o�t�6�4��D��6�5��į6�6��6�7��6���W�R�9_�d�3��� 6�9���6�a�ܿ6��� �6���,�6�ٯT�6� �|�6�)���6�Q��� 6�y���^����^�ʿ D�^��l�^�ϔ�^� Bϼ�^�j���^���� ^���4�^���\�^�
� �2���6��/� ���V��<�'�`�K� ��o����������� ��&J5nY� ������� 4F1jU�y� ����/�0// T/?/x/c/�/�/�/�/ �/�/�/??>?)?P?�t?_?�?
�_DEV� I�M{C:�84���4?GRP 2/E�0�+�bx 	�� 
 ,@�0 �?OD8OJO1OnOUO �O�O�O�O�O�O�O�O "_	_F_-_j_|_c_�_ �[O�_�_�_o�_,o oPo7oIo�omo�o�o �o�o�o�o(:!\^�_  �0i @�������  �=�$�a�s�Z���~� �������؏�l
�@K���qp�W��Q�� ����ϟ��ڟ�)� �M�4�]���j����� ˯ݯ�_����7�� [�B����x�����ٿ �ҿ���3��,�i� Pύ�䯾���^����� ���޹�'��v�]� �߁߾��߷������ *��N��r��;�� �����������&�8� �\�C���g�y����� ������g�4- jQ�u���� �B)fx _����)�� /,//P/7/t/[/m/ �/�/�/�/�/?�/(?�?L?^?E?�?�7d ��[~
�6 �s 	 A;�*=� 6?�=����D�>ޟ���g�:�0���ī��|@��-�@�5_�eA5�-�=�BG+h�&����6)AB�m�����`x���=�?7O%TEL�EOP8OcN[~�y��5�o�ʾ�TF�����������|��ҝ����E��1�E@�*��A`�~�n��!��$�A����M�Y<T�������C=��J����Gc��McO��IJO/_��[~��6r� _�1<�׻���y;��	A�`�ʛ1bP��N	�V�A�&@���@���@)�E�]�1������0ד� x����Q��U?�Q��O�__ _�oDU�NU9���6>���E��bQ�2]�j_ ���rAS��AT�@���@G$�_ ���yC� �Pr�}��Q� 2i?�R�_�o�_�_�o�DU�K�5��l�������S����`
�� 3�>v�ĚM@��@�V�@��%@��Ŀ�qߝ��]V�N���N�!C(u�µ�� �®�ɒow�o �o�DS�I�I���`�"��2�X�%�� ��hoZ�����؏Ə�� � �b�G����z�� ������ԟ��:�� ^��R�@�v�d����� ��Я���6���*�� N�<�r�`������Ͽ �����&��J�8� nϰ��ϧ�^π�Z��� ����"��F߈�m߬� 6ߠߎ߲߰������� �`�E���x�f�� ��������8��\� ��P�>�t�b������� ��$���4���(L :p^������� ���$H6l ���\���� � //D/�k/�4/ �/�/�/�/�/�/�/? ^/C?�/?v?d?�?�? �?�?�?$?	OO�?�? �?<OrO`O�O�O�O�? �O O�O__$_&_8_ n_\_�_�O�_�O�_�_ �_o�_ o"o4ojo�_ �o�_Zo�o�o�o�o �oro�oi�oB� ������J/� n�b��r������� ����"��F�Џ:�(� ^�L�n���������ߟ ���� �6�$�Z�H� j���ҟ�������د ���2� �V���}��� F�h�B����Կ
��� .�p�Uϔ�ψ�vϘ� �Ϭ������H�-�l� ��`�N߄�rߔߖߨ� �� ��D���8�&�\� J��n�������� �����4�"�X�F�|� �����l���h��� ��0T��{��D ������, nS��t�� ���/F+/j� ^/L/�/p/�/�/�// �/?�/�/�/$?Z?H? ~?l?�?�/�??�?�? �?OO OVODOzO�? �O�?jO�O�O�O�O_ 
__R_�Oy_�OB_�_ �_�_�_�_�_oZ_�_ Qo�_*o�oro�o�o�o �o�o2oVo�oJ�o Z�n���
� .�"��F�4�V�|� j����Ǐ������ ��B�0�R�x����� ޏh�ҟ������� >���e�w�.�P�*��� ί�����X�=�|� �p�^�������ʿ�� �0��T�޿H�6�l� Z�|�~ϐ������,� �� ��D�2�h�V�x� ������ߞ������ 
�@�.�d�ߋ���T� ��P���������<� ~�c���,��������� ������V�;z� n\������ .R�F4jX �|������ �/B/0/f/T/�/� �/�z/�/�/�/�/? >?,?b?�/�?�/R?�? �?�?�?�?�?O:O|? aO�?*O�O�O�O�O�O �O�OBOhO9_xO_l_ Z_�_~_�_�_�__�_ >_�_2o�_BohoVo�o zo�o�_�oo�o
�o .>dR��o� �ox����*�� :�`�����P����� ޏ̏���&�h�M�_� �8��������ڟȟ ��@�%�d��X�F�h� j�|�����֯���<� Ư0��T�B�d�f�x� ���տ������,� �P�>�`϶�ܿ��� ���������(��L� ��s߲�<ߦ�8߶��� �� ���$�f�K��� ~�l���������� >�#�b���V�D�z�h� �����������:��� .R@vd��� ������* N<r���b� ����&//J/� q/�:/�/�/�/�/�/ �/�/"?d/I?�/?|? j?�?�?�?�?�?*?P? !O`?�?TOBOxOfO�O �O�OO�O&O�O_�O *_P_>_t_b_�_�O�_ �O�_�_�_oo&oLo :opo�_�o�_`o�o�o �o�o "H�oo �o8������ �P5�G�� ��h� �������(��L� ֏@�.�P�R�d����� �� ��$�����<� *�L�N�`���؟���� ���ޯ��8�&�H� ��į��ԯn�ȿ��� ڿ���4�v�[Ϛ�$� �� Ϟ��ϲ������ N�3�r���f�Tߊ�x� ���߮���&��J��� >�,�b�P��t��� ����"����:�(� ^�L��������r��� n��� 6$Z�� ���J����� �2tY�"� z�����
/L 1/p�d/R/�/v/�/ �/�//8/	?H/�/<? *?`?N?�?r?�?�/�? ?�?O�?O8O&O\O JO�O�?�O�?pO�O�O �O�O_4_"_X_�O_ �OH_�_�_�_�_�_�_�
o0or_Wo�U�P��$SERV_MA_IL  �U�`���QvdOUTPU}T�h�P}@vdRV 20f;  �` (a\o<�ovdSAVE�l�i�TOP10 21��i d 6� s�P6r _�P2oXj|�� �������0� B�T�f�x��������� ҏ�����,�>�P� b�t���������Ο������(�:�guY�P�cFZN_C�FG 2e��c�T�a�e|�GR�P 23��q ?,B   AƠ�Q�D;� BǠ��  B4�SR�B21�fHELL��4ev�`�o���/�>�%RSR >�?�Q���u�����ҿ ������,��P�;��t�_Ϙϩ����?p�¼����Ϸͻ���P�&�'���W��2�Pd��gҾ�HK 15�� ,ߡ߫ߥ����� ����@�;�M�_�� �������������?OMM 6��?���FTOV_EN�B�d�au�OW_?REG_UI_��b�IMIOFWDL�*�7.�ɥ��WAIT\�`ٞ����`����d��TIM������VA�`����_UNIT[�*y�LCy�TRY��Zuv`ME�8����aw֑d ��9�[ �����<��X�Pڠ6p`?�  ��o+`=IpVL�l��fMON_ALI_AS ?e.��`heGo����� �/)/;/M/�q/�/ �/�/�/d/�/�/?? %?�/I?[?m??�?<? �?�?�?�?�?�?!O3O EOWOO{O�O�O�O�O nO�O�O__/_�OS_ e_w_�_�_F_�_�_�_ �_�_o+o=oOoaoo �o�o�o�o�oxo�o '9�o]o�� >������#� 5�G�Y�k�������� ŏ׏������1�C� �g�y�����H���ӟ ���	���-�?�Q�c� u� �������ϯᯌ� ��)�;��L�q��� ����R�˿ݿ��� ��7�I�[�m��*ϣ� �������ϖ��!�3� E���i�{ߍߟ߱�\� ����������A�S� e�w��4������� �����+�=�O���s� ��������f����� '��K]o�� >�����# 5GY}�����l�$SMON�_DEFPROG &����� &*SYSTEM*����RECALL� ?}� ( ��}3xcopy� fra:\*.�* virt:\tmpbackU!�=>192.16�8.56.1:4772 {!�/�/�/��-}7L$s:or�derfil.datY,k/�/?$?6?{}.L"mdb:V/�/2 �/�?�?�?�%2K%T/f/x$~?O!O 3O�!J/�?n/ O�O�O �O�/�/c?�?_!_3_ F?�Oj?�O�_�_�_�? WOiO�?oo/oBO�_��_xO�o�o�o�G
x�yzrate 11 Vohozo/��E�g�l15344 �o�o����C�tpdisc 0Ugphz��/���Etpconn 0 ����������G8�O�O�gp��'��M/K_�^y�� ������CmTo�obu��"�4��@4KoܟY~  ��������oZ�l�~� �!�3�F������ �����n�h�z���/�¯1 ������ȝϯ��EK�s�2796 i�{���0��D˿�����ϊߜ� ��A�S�b�t���)� <�N����߃���:� ����d�v���+��O ЏY��̓�����:_L� g���{�0�_�� ��������FoW i��"4G�Y� ���������`�� {//0/C��y �/�/�/��d/�? ?,??Q�u�?�? �?��j?�OO(O ;/M/�/q/�O�O�O�/ �/\O�/�O_$_6_I? [?�?�O�_�_�_�?b_��?}_o o2oā�$�SNPX_ASG 2:���Va��  �0ā%�7o~o  �?�GfPARAM� ;Ve`a W�	lkP��Ā����d� ���I`OFT_KB_CFG  Ã�\eFcOPIN_S_IM  Vk�b�+=OYsI`RV�NORDY_DO�  �eukrQSTP_DSB~��b�>kSR �<Vi � & ?TELEO�e��{v��W`I`TOP_?ON_ERRxGb~�PTN Ve�P��D:�RING_PRM'���rVCNT_GP� 2=Ve�ac`x 	���DP��я�����BgVD�RP 1>�i�`�Vq؏ 0�B�T�f�x������� ��ҟ�����,�>� e�b�t���������ί ���+�(�:�L�^� p���������ʿ��  ��$�6�H�Z�l�~� �Ϸϴ����������  �2�D�V�}�zߌߞ� ����������
��C� @�R�d�v����� ����	���*�<�N� `�r������������� ��&8J\n �������� "4[Xj|� ������!// 0/B/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?t?�?�?�?�?�?��?�?O�PRG_�COUNT�f�P�)IENBe�+EM�UC�dbO_UPD �1?�{T  
 ODR�O�O�O�O�O_ _A_<_N_`_�_�_�_ �_�_�_�_�_oo&o 8oao\ono�o�o�o�o �o�o�o�o94F X�|����� ����0�Y�T�f� x������������� �1�,�>�P�y�t��� ������Ο��	��� (�Q�L�^�p������� ���ܯ� �)�$�6� H�q�l�~�������ƿ ؿ���� �I�D�V��"L_INFO 1=@�E�@��	 yϽϨ������?���?���>MNe=����� A��PA��w�ǼiA��'.�gEB�<������@ ?j` =@���o� D<Ş�B�Q_DF�C�@���B�I�p߂�-@Y?SDEBUG:@�@��o�d�I��SP_�PASS:EB?~��LOG A��]�A  o�i��v�  �Ao�UD1:\��}���_MPC�ݚEk�}A&�� �AK�SAV B��IA����*�i�1�SV�B�TEM_TIM�E 1C���@k 0o�n��i��{��*���MEMBOK  �EA��������X|f�@� Z�i���� ������h�9
�� ��@�`r� ������� �@Rdv@�����
Le� //(/:/L/^/p/�/ �/�/�/�/�/�/ ??`$?6?H?Z?��SKV��[�EAj��?�?�?��	%�@0]2���?i�  0�o�^
 :O.@R�O�O�O}N��2F ��OBD��O_'_9_-L2�Y_�_�_�_�_�_o�U�_�_�o'o 9oKo]ooo�o�o�o�o �o�o�o�o#5G�Yk_?T1SVG�UNSPD�� '�����p2MOD�E_LIM D���Ҋt2�p�qE��݉uABUI_D�CS H}5���0�G�n��D��|�-�X�>���*���� 
��e��C����r�i�����uE?DIT I��xSCRN J��y�rS�G K��.�(�0߅SK_OPTION��^�����_DI��ENB�  -����BC�2_GRP 2L����MPC��ʓ�|BCCF/�N����� ����`�>�W�B�g���x� ����կ������� �S�>�w�b������� ��Ͽ�����=�(� a�Lυϗ�Ň�϶��� ����v��
�/�U�@� yߧ��`�iМ��߰� ����
���.��>�@� R��v�������� ���*��N�<�r�`� ��������������̀ 4FX��|j ������� B0fTvx� ����/�,// </b/P/�/t/�/�/�/ �/�/�/�/(??L? d?v?�?�?�?6?�?�? �?O O6OHOZO(O~O lO�O�O�O�O�O�O�O  __D_2_h_V_�_z_ �_�_�_�_�_
o�_.o o>o@oRo�ovo�ob? �o�o�o�o<* Lr`����� ���&��6�8�J� ��n�����ȏ���ڏ ��"��F�4�j�X��� |��������֟��o $�6�T�f�x������� ��ү�������>� ,�b�P���t������� �ο��(��L�:� \ς�pϦϔ��ϸ��� ���� ��H�6�l�"� �ߖߴ�����V����� �2� �V�h�z�H�� �������������
� @�.�d�R���v����� ��������*N <^`r����� ��&8�\J l������� �"//F/4/V/X/j/ �/�/�/�/�/�/?�/ ?B?0?f?T?�?x?�? �?�?�?�?O�?,O� DOVOtO�O�OO�O�O��O�O�O_ V4P�$�TBCSG_GR�P 2O U��  �4Q 
 ?�  __ q_[_�__�_�_�_�_��_o%k8R?SQF\_d�HTa?4Q	 HA���#e�>���>$a��\#eAT��A �WR�o�hdjma�G��?Lfg�bp�o�n�;ffhf��ͼb4P�|j��o*}@��R�hf�ff>�33pa#e<qB�o+=xr�Rp�qUy�rt~҃�H�y rIpTv�pBȺt~	xf	x(�;� ��f���N�`���ˏ�ڋ����	V3�.00WR	cr;xlڃ	*���3R~t��HH��� q\�.�]�  c�C.�����8QJ2�?SRF]����CFoG T UPQY SPܚ��r�9ܟ1��1�W� e�	Pe���v�����ӯ ��������Q�<� u�`���������Ϳ� ޿��;�&�_�Jσ� nπϹϤ������� WRq@�0�B���u�`� �߫ߖ��ߺ������ )�;�M��q�\��� ����4Q _���O �� �J�8�n�\������� ����������4" XFhj|��� ���.TB xf��nO��� �//>/,/b/P/�/ t/�/�/�/�/�/�/�/ ?:?(?^?p?�?�?N? �?�?�?�?�?�? O6O $OZOHO~OlO�O�O�O �O�O�O�O __D_2_ T_V_h_�_�_�_�_�_ �_
o�_o@o�Xojo |o&o�o�o�o�o�o �o*N`r�B �������&� �6�\�J���n����� ȏ��؏ڏ�"��F� 4�j�X���|���ğ�� �֟���0��@�B� T���x�����ү䯎o ���̯ʯP�>�t�b� ������������� Կ&�L�:�p�^ϔϦ� ���τ������ �"� H�6�l�Zߐ�~ߴߢ� ���������2� �V� D�z�h�������� �����
�,�.�@�v� ������\������� <*`N�� ��x��� 8J\(��� �����/4/"/ X/F/|/j/�/�/�/�/ �/�/�/??B?0?f? T?v?�?�?�?�?�?�? OO��2ODO�� O�O tO�O�O�O�O�O_�O (_:_L_
__�_p_�_ �_�_�_�_ o�_$oo 4o6oHo~olo�o�o�o �o�o�o�o D2 hV�z���� �
��.��R�@�b� ��v���&OXO֏菒� ����N�<�r�`��� ����̟ޟ🮟�� $�&�8�n�������^� ȯ���گ��� �"� 4�j�X���|�����ֿ Ŀ����0��T�B� x�fψϊϜ������� ����>�P���h�z� ��6߼ߪ��������� �:�(�^�p���R��������� ���  9&�*� *�>��*��$TBJOP_GRP 2U����  ?���C*�i	V�]�Wd������X � *��� ��, � ����*� @&�?���	 �A���~��C�  DD������>v�>\�? ��aG�:��o��;ߴ�AT������A�@<��MX����>���\)?����8Q�����L���>�0 &�;iG.��Ap< � F�A�ff�v��� ):VMՂ.�� S>o*�@w��R�Cр	���������f�f�:�6/�?��33�B    ��/�������>):�S����� �/�/@��H@�%&/�/��=� �<#�
*��v�;7/�ڪ!?���4B�3?'?2	��2? hZ?D?R?�?�?�?F? �?�?�?�?OAOO�?�`OzOdOrO�O�O*�C�*���A��	V�3.00{�crxl��*P��%��%c5Z F�� JZH F6�� F^ F��� F�f F�� G� G�5 G<
 G^�] G� G����G�*�G��S G�; G���ERDu�\E[�� E� F�( F-� FU�` F}  F��N F� F��� Fͺ F��� F�V G�� Gz G?a 9ѷ�Q�L�HefJ4�o,b�*�0c1���OH�E�D_TCH XXd�+X2S�&�&�d$'X�o�o*�1�F�TESTPARS  ��cV��HRpABLE ;1Yd� N`*�H�����g$j�g�h��h)�1��g	�h
��h�hHu*��h��h�h%vRDI0n�GYk}��u	�O�#�-�?�Q�Hc�u�)rS�l� �z 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z���I���m� Fwͩ��ȏڏ쏘������x)r��NUoM  ��n���2� Ep�)r_CFG Z���I���@V�IMEB�F_TTqD��e�޶VER������޳R 1[8{ �8�o*�%�Q� ��د  9�K�]�o� �ϓϥϷ��������� �#�5�G�Y�k�}��� �߳����������� 1���E�W�i�{��� ������������/� A�S�e�w��������� ������+=OR�_���@��`�LIF \��	D`����DR�](FP
�!p�!p�� d� ��MI_�CHAN� � ~DBGLVL���fETHER�AD ?u���0`1�_}�R�OUT�!�j!���SNMA�SKY�j255.%S///A/S��`OOLOFS_�DIp�COR�QCTRL ]8{��1o�-T�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OL�/6O%OZOcPE_�DETAI7�*P�GL_CONFI�G c�������/cell/$�CID$/grp1^O�O�O�O
__|���G_Y_k_}_�_�_ 0_�_�_�_�_oo�_ CoUogoyo�o�o,o>o �o�o�o	-�oQ cu���:�� ���)���_�q� ��������׮}N�� ��%�7�I�a�KOq�P��M�����ʟܟ�  �G�$�6�H�Z�l�~� �����Ưد���� ��2�D�V�h�z���� ��¿Կ���
ϙ�.� @�R�d�vψϚ�)Ͼ� �������ߧ�<�N� `�r߄ߖ�%ߺ����� ����&��J�\�n� ����3��������� �"���F�X�j�|���������@�Us�er View ��I}}1234567890�����+=Ex �e����2��B����@��`r��3� Oas����x4>//'/9/K/]/�~/x5��/�/��/�/�/?p/2?x6 �/k?}?�?�?�?�?$?�?x7Z?O1OCOUO gOyO�?�Ox8O�O �O�O	__-_�ON_TR� lCamera���O�_�_ �_�_�_�_˂E�_o )o;n��Uogoyo�o�o�o�)  mV�	�_�o #5GY o}� ��o������F_�mV=�k�}��� ����ŏl����X� 1�C�U�g�y���2�D� �"�ן�����1� ؏U�g�y�ğ������ ӯ�����D��k��E� W�i�{�����F�ÿտ �2���/�A�S�e� �nUY9���������� ��	߰�-�?�Qߜ�u� �ߙ߽߫���v�D�I f��-�?�Q�c�u�� ����������� )�;���D��I����� ����������) t�M_q���N�`�93��0 B��Sx�1��@���//�J	oU0�U/g/y/�/�/�/ V�/�/�/�?-??? Q?c?u?/./tPv[? �?�?�?OO(O�/LO ^OpO�?�O�O�O�O�O �O�?oU�k�O:_L_^_ p_�_�_;O�_�_�_'_  oo$o6oHoZo_;% N��_�o�o�o�o�o  �_$6H�ol~� ���moe��]� $�6�H�Z�l����� ���؏���� �2� �e&�ɏ~������� Ɵ؟���� �k�D� V�h�z�����E�e�� 5����� �2�D�� h�z���ׯ��¿Կ�x��
ϱ�  �� 9�K�]�oρϓϥϷ����������    ��5�G�Y�k�}ߏ� �߳����������� 1�C�U�g�y���� ��������	��-�?� Q�c�u����������� ����);M_�q�  
��( � �-�( 	 ������� #35G}k����
� � Y�
//./��R/d/v/ �/�/�/����/�/�/ A/?0?B?T?f?x?�/ �?�?�??�?�?OO ,O>O�?bOtO�O�?�O �O�O�O�O_KO]O:_ L_^_�O�_�_�_�_�_ �_#_ oo$ok_HoZo lo~o�o�o�_�o�o�o 1o 2DVh�o �o���	��
� �.�@��d�v���� ����Џ���M�*� <�N���r��������� ̟�%���&�m�J� \�n��������ȯگ �3��"�4�F�X�j� ����������ֿ��� ��0�w���f�xϊ� ѿ�����������O� ,�>�Pߗ�t߆ߘߪ� ���������]�:�L�^�p����߻@� ������������ ��"frh�:\tpgl\r�obots\cr�x!�10ia_l.xml��D�V�h� z�������������������0BTf x�������� �,>Pbt� �������/ (/:/L/^/p/�/�/�/ �/�/�/��/?$?6? H?Z?l?~?�?�?�?�? �?�/�?O O2ODOVO hOzO�O�O�O�O�O�? �O
__._@_R_d_v_ �_�_�_�_�_�O�_o o*o<oNo`oro�o�o��o�o�o�n �6�� ���<< 	� ?��k!�o ;iOq��� ������%�S� 9�k���o�����я�����(�$TPG�L_OUTPUT� f������ �&�8�J� \�n���������ȟڟ ����"�4�F�X�j��|�������į�p��ր2345678901�����1� C�K����r������� ��̿d�п��&�8�J��}T�|ώϠϲ� ��\�n�����0�B� T���bߊߜ߮����� j�����,�>�P��� �߆��������x� ���(�:�L�^���l� ����������t��� $6HZlz� ������ 2 DVh ��� ����/./@/R/ d/v//�/�/�/�/�/��/�/ۂ $$��ί<7*?\?N?�? r?�?�?�?�?�?�?O O4O&OXOJO|OnO�O �O�O�O�O�O_�O0_"_T_}�an_�_�_�_�_�_�]@�_o	z ( 	 V_ Do2ohoVo�ozo�o�o �o�o�o
�o.R @vd����� ����(�*�<�r��`���ܦ�  <<I_ˏݏ��� ����:�L�֪��}� ��)���ş������� k��C�ݟ/�y���e� ������������-� ?��c�u�ӯ]����� W���Ϳ��)χ��� _�q��yϧρϓ��� ��M��%߿��[�5� Gߑߣ�߫���s��� �!���E�W��?�� ��9���������i� ��A�S���w���c�u� ���/�����= )s�����U ���'9�! o	[����� K�#/5/�Y/k/E/ w/�/�/�/�/�/�/ ?�/?U?g?�/�?�? 7?�?�?�?�?	OO���)WGL1.X�ML�_PM�$TP�OFF_LIM ����P����^FN_SVf@  ��TxJP_MOoN g��zD��P�P2ZISTRTCHK h���xFk_aBVTCO�MPAT�HQ|FVWVAR i�M�:X�D �O �R_�P�BbA_D�EFPROG �%�I%TEL�EOPi_�O_DISPLAYm@�N�R�INST_MSK�  �\ �ZI�NUSER_�TL�CKl�[QUIC�KMEN:o�TSC�REY`��Rtpsc�Tat`hyixB�`_�iSTZ�xIRACE_CF�G j�I:T��@	[T
?��hHNL 2k�Z���aA[ gR-?Qcu�����z�eITE�M 2l{ ��%$123456�7890 ��  �=<
�0�B�J�  #!P�X�dP��� [S���"���X�
� |���W���r�֏���� .��0�B�\�f����� 6�\�n�ҟ������ ��>���"���.��� ��ίR����Ŀֿ:� �^�p�9ϔ�Tϸ�x� ����d���H�� l��>�Pߴ�\����� ��v� ������h�(� �ߞ߰�4�L��ߦ�� ���@�R��v�6��� Z�l���������*� ��N��� �������� ����X���J 
n���b� ���"4F�/ |</N/�Z/���/ /�/0/�/?f/?�/ �/e?�/�?�/�?�?�? ,?�?P?b?t?�?�?DO jO|O�?�OOO(O�O �O^O_0_�O<_�O�O �_�O�__�_�_H_�_Pl_~_Go�dS�bm�o>Lj�  �rLj� �a�o�Y
 �o�o�o�o{jUD�1:\|��^aR_GRP 1n�{�� 	 @ �PRd{N�r����~��p���q�+��O�:�?�   j�|�f���������� ҏ����>�,�b�P����t���������	�e���\cSCB ;2ohk U�R� d�v���������Я��RlUTORIAL� phk�o-�WgV�_CONFIG qhm�a�o�o��<��OUTPUT yrhi}����� ܿ� ��$�6�H�Z� l�~ϐϢϴ�z�ɿ�� �� ��$�6�H�Z�l� ~ߐߢߴ��������� � �2�D�V�h�z�� �����������
�� .�@�R�d�v������� ��������*< N`r������ ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/��/�/? ?0?B?T?f?x?�?�? �?�?�/�?�?OO,O >OPObOtO�O�O�O�O �?�O�O__(_:_L_ ^_p_�_�_�_�_�_f� x�ǿoo,o>oPobo to�o�o�o�o�o�o�O (:L^p� ������o �� $�6�H�Z�l�~����� ��Ə؏��� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ���*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b� t���������������>�X���# ��N�_r��� ����&8 J��n����� ���/"/4/F/X/ i|/�/�/�/�/�/�/ �/??0?B?T?e/x? �?�?�?�?�?�?�?O O,O>OPOa?tO�O�O �O�O�O�O�O__(_ :_L_^_oO�_�_�_�_ �_�_�_ oo$o6oHo Zok_~o�o�o�o�o�o �o�o 2DVgo z������� 
��.�@�R�d�u�� ������Џ���� *�<�N�`�q������� ��̟ޟ���&�8��J�\�k��$TX_�SCREEN 1}s% �}�k�����ӯ���	���Z��I�[� m�������,�ٿ� ���!�3Ϫ�W�ο{� �ϟϱ�����L���p� �/�A�S�e�w��� � �߿��������~�+� ��O�a�s���� � ��D�����'�9�K� ��������������� R���v�#5GYk�}����$UAL�RM_MSG ?5����� �n� ��	:-^Q c������ /~�SEV  ��2&�ECFG� u���� � n�@�  A�b!   B�n�
 /u����/�/�/ �/�/�/??%?7?I?�W7>!GRP 2v�H+ 0n�	 �/�?� I_BBL�_NOTE w�H*T���lu���w�T �2D_EFPRO� %� (%�Ow�	O�BO-BTELEOPGO#O�O�O�O�O�O��O�O_�O&_�?�0F�KEYDATA �1x���0p W'n��?�_�_z_�_��_�Z,(�_on�(�POINT E�Ron  IREcCT@oko�PNDUo��oOcCHOICE�]�onTOUCHU`O�o�_�o7 [mT�x�� ����!��E��Z���/frh/�gui/whit�ehome.pn�gQ�������ŏ׏�}h�pointz����/�A�S��  >i�direc����࡟��şןf�/in y��"�4�F�X��m�choicy�����л�ͯ߯�h�touchup���/��A�S�e��h�arwrg�����ÿտ �n���(�:�L�^� p����Ϧϸ������� }��$�6�H�Z�l��� �ߢߴ��������ߋ�  �2�D�V�h�z�	�� ������������.� @�R�d�v���_����� ���������2D Vhz���� ��
�@Rd v��)���� //�</N/`/r/�/ �/%/�/�/�/�/?? &?�/J?\?n?�?�?�? 3?�?�?�?�?O"O�? 4OXOjO|O�O�O�OAO �O�O�O__0_�OT_ f_x_�_�_�_=_�_�_ �_oo,o>o�_boto��o�o�o�oW��k}�b�����o@}�o8J$v,6� {.������� ��/��S�:�w��� p�����я�ʏ�� +��O�a�H���l��� ����ߟ���'�9� Ho]�o���������ɯ X�����#�5�G�֯ k�}�������ſT�� ����1�C�U��y� �ϝϯ�����b���	� �-�?�Q���u߇ߙ� �߽�����p���)� ;�M�_��߃���� ����l���%�7�I� [�m������������ ��z�!3EWi ��������� П/ASew~ ������/� +/=/O/a/s/�//�/ �/�/�/�/?�/'?9? K?]?o?�?�?"?�?�? �?�?�?O�?5OGOYO kO}O�OO�O�O�O�O �O__�OC_U_g_y_ �_�_,_�_�_�_�_	o o�_?oQocouo�o�o �o:o�o�o�o) �oM_q���6 �����%�7��9�����b�t���^�������,��돞����3� E�,�i�P�������ß ���������A�S� :�w�^�������ѯ�� ��ܯ�+�
O�a�s� �������Ϳ߿�� �'�9�ȿ]�oρϓ� �Ϸ�F��������#� 5���Y�k�}ߏߡ߳� ��T�������1�C� ��g�y������P� ����	��-�?�Q��� u�����������^��� );M��q� �����l %7I[��� ���h�/!/3/ E/W/i/@��/�/�/�/ �/�/�??/?A?S? e?w??�?�?�?�?�? �?�?O+O=OOOaOsO O�O�O�O�O�O�O_ �O'_9_K_]_o_�__ �_�_�_�_�_�_�_#o 5oGoYoko}o�oo�o �o�o�o�o�o1C Ugy���� ��	���?�Q�c� u�����(���Ϗ�� ����;�M�_�q���h����~ ���~ ���ҟ���Ο�*��,�[�� �f�������ٯ���� ���3��W�i�P��� t���ÿ���ο�� /�A�(�e�Lωϛ�z/ ����������(�=� O�a�s߅ߗߩ�8��� ������'��K�]� o����4������� ���#�5���Y�k�}� ������B������� 1��Ugy�� ��P��	- ?�cu���� L��//)/;/M/ �q/�/�/�/�/�/Z/ �/??%?7?I?�/m? ?�?�?�?�?�?���? O!O3OEOWO^?{O�O �O�O�O�O�OvO__ /_A_S_e_�O�_�_�_ �_�_�_r_oo+o=o Ooaosoo�o�o�o�o �o�o�o'9K] o�o������ ��#�5�G�Y�k�}� �����ŏ׏����� �1�C�U�g�y���� ����ӟ���	���-� ?�Q�c�u��������@ϯ�����0����0����B�T�f�>�����t�, ��˿~��ֿ�%�� I�0�m��fϣϊ��� ��������!�3��W� >�{�bߟ߱ߘ��߼� ����?/�A�S�e�w� ����������� ���=�O�a�s����� &����������� 9K]o���4 ����#�G Yk}��0�� ��//1/�U/g/ y/�/�/�/>/�/�/�/ 	??-?�/Q?c?u?�? �?�?�?L?�?�?OO )O;O�?_OqO�O�O�O �OHO�O�O__%_7_ I_ �m__�_�_�_�_ �O�_�_o!o3oEoWo �_{o�o�o�o�o�odo �o/AS�ow ������r� �+�=�O�a������ ����͏ߏn���'� 9�K�]�o��������� ɟ۟�|��#�5�G� Y�k���������ůׯ ������1�C�U�g� y��������ӿ��� ���-�?�Q�c�uχ��^P���^P��������ͮ���
���,��;���_�F� �ߕ�|߹ߠ������� ���7�I�0�m�T�� �����������!� �E�,�i�{�Z_���� ���������/A Sew���� ���+=Oa s������ //�9/K/]/o/�/ �/"/�/�/�/�/�/? �/5?G?Y?k?}?�?�? 0?�?�?�?�?OO�? COUOgOyO�O�O,O�O �O�O�O	__-_�OQ_ c_u_�_�_�_:_�_�_ �_oo)o�_Mo_oqo �o�o�o�o���o�o %7>o[m� ���V���!� 3�E��i�{������� ÏR������/�A� S��w���������џ `�����+�=�O�ޟ s���������ͯ߯n� ��'�9�K�]�쯁� ������ɿۿj���� #�5�G�Y�k����ϡ� ��������x���1� C�U�g��ϋߝ߯�����������`���>�`���"�4� F��h�z�T�,f��� ^���������)�� M�_�F���j������� ������7[ B�x���� �o!3EWix� �������� ///A/S/e/w//�/ �/�/�/�/�/�/?+? =?O?a?s?�??�?�? �?�?�?O�?'O9OKO ]OoO�OO�O�O�O�O �O�O_�O5_G_Y_k_ }_�__�_�_�_�_�_ o�_1oCoUogoyo�o �o,o�o�o�o�o	 �o?Qcu��( ������)�  M�_�q��������ˏ ݏ���%�7�Ə[� m��������D�ٟ� ���!�3�W�i�{� ������ïR����� �/�A�Яe�w����� ����N������+� =�O�޿sυϗϩϻ� ��\�����'�9�K� ��o߁ߓߥ߷����� j����#�5�G�Y��� }��������f�����1�C�U�g�>��i��>������������������,��?&cu \������� )M4q�j �����/�%/ /I/[/:�/�/�/�/ �/�/���/?!?3?E? W?i?�/�?�?�?�?�? �?v?OO/OAOSOeO �?�O�O�O�O�O�O�O �O_+_=_O_a_s__ �_�_�_�_�_�_�_o 'o9oKo]ooo�oo�o �o�o�o�o�o�o#5 GYk}��� �����1�C�U� g�y��������ӏ� ��	���-�?�Q�c�u� ����p/��ϟ��� ��;�M�_�q����� ��6�˯ݯ���%� ��I�[�m������2� ǿٿ����!�3�¿ W�i�{ύϟϱ�@��� ������/߾�S�e� w߉ߛ߭߿�N����� ��+�=���a�s�� ����J������� '�9�K���o������� ����X�����#5 G��k}���������������&�HZ4,F/�>/� ����	/�-/?/ &/c/J/�/�/�/�/�/ �/�/�/?�/;?"?_? q?X?�?|?�?�?���? OO%O7OIOXmOO �O�O�O�O�OhO�O_ !_3_E_W_�O{_�_�_ �_�_�_d_�_oo/o AoSoeo�_�o�o�o�o �o�oro+=O a�o������ ���'�9�K�]�o� �������ɏۏ�|� �#�5�G�Y�k�}�� ����şן������ 1�C�U�g�y������ ��ӯ���	��?-�?� Q�c�u���������Ͽ ���Ϧ�;�M�_� qσϕ�$Ϲ������� �ߢ�7�I�[�m�� �ߣ�2���������� !��E�W�i�{��� .�����������/� ��S�e�w�������<� ������+��O as����J� �'9�]o ����F����/#/5/G/�$UI�_INUSER � ���h!��  �H/L/_MENHI�ST 1yh%�  ( �u ��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1�/�/?�?0?�)�/�/13@�/|?�?�?�?�'E?W>71l?�?O#O5O��+�?W5edit~�"TELEOP�?��O�O�O:O�?�?32,2�O	__-_?_�O�Oe,2k?�_�_�_p�_��/f_148�O o"o4oFo��Iono@�o�o�o�o�o��\a �!\o�o/AS Vow�����` ���+�=�O��� ��������͏ߏn�� �'�9�K�]�쏁��� ����ɟ۟j�|��#� 5�G�Y�k��������� ůׯ��o�o�1�C� U�g�y�|�������ӿ ������-�?�Q�c� uχ�ϫϽ������� ߔ�)�;�M�_�q߃� ߧ߹��������� ��7�I�[�m��� � �������������� E�W�i�{��������� ��������AS ew���<�� �+�Oas ���8���/ /'/9/�]/o/�/�/ �/�/F/�/�/�/?#? 5? �2�k?}?�?�?�? �?�/�?�?OO1OCO �?�?yO�O�O�O�O�O bO�O	__-_?_Q_�O u_�_�_�_�_�_^_p_ oo)o;oMo_o�_�o �o�o�o�o�olo�%7I[F?��$�UI_PANED�ATA 1{�����q � 	�}  f�rh/cgtp/�flexdev.�stm?_wid�th=0&_height=10�p��pice=TP&�_lines=1�5&_colum�ns=4�pfon�t=24&_pa�ge=whole��pmI6)  rim�9�  �pP�b� t������������Ǐ ��(�:�!�^�E��� ��{�����ܟ�՟��I6� �  7 Y1�VJ�O� a�s���������ͯ@� ���'�9�K���o� ��h�����ɿۿ¿�� �#�5��Y�@�}Ϗ�vϳ�&��Ɠs��� ��)�;�Mߠ�q�� �ߧ߹�������V�� %��I�0�m��f�� �����������!�� E�W����ύ������� ����:�~�/AS ew����� � =$as Z�~����d� v�'/9/K/]/o/�/� �/�/*�/�/�/?#? 5?�/Y?@?}?�?v?�? �?�?�?�?O�?1OCO *OgONO�O�/�/�O �O�O	__-_�OQ_�/ u_�_�_�_�_�_6_�_ o�_)ooMo_oFo�o jo�o�o�o�o�o�o %7�O�Om�� ���^_�!�3� E�W�i�{������Ï ���������A�S� :�w�^�������џD V��+�=�O�a��� ����
���ͯ߯�� �|�9� �]�o�V��� z���ɿ���Կ�#��
�G�.�k�ޟ�}��|ϵ����������) ��4ߧ�#�`�r߄ߖ� �ߺ�!���������� 8��\�C���y�� �����������������$UI_POSTYPE  ���� 	 ��s�B�QUICKMEN  Q��`�v�D�REST�ORE 1|���  �	�����������mASew�, ������+ =Oan�� ���//�9/K/ ]/o/�/�/6/�/�/�/ �/�/�??0?�/k? }?�?�?�?V?�?�?�? OO�?COUOgOyO�O 6?@O�O�O.O�O	__ -_?_Q_�Ou_�_�_�_ �_`_�_�_oo)o�O 6oHoZo�_�o�o�o�o �o�o%7I[��o������S�CRE��?���u1sc���u2�3�4�5*�6�7�8��swTATM�� ��<��:�USER�p�2�rT�p�ks���U4��5��6��7���8��B�NDO_CFG }Q������B�PDE���?None��v��_INFO 2~j��)���0%� D���2�s�V������� ͟ߟ��'�9���]�o�R���z��OFFSET �Q�-���hs��p��� ��G�>�P�}�t��� Я��׿ο���� C�:�L�^Ϩ����͘ς��
����av��W�ORK �!������.�@ߢ�u�UFRAME  ����RTOL_A�BRT�����EN�B�ߣ�GRP 1������Cz  A������*�<�N�`�r��֐�U������MSK  ��)���N��%�!��%z����_EVN�����+�ׂ�3�«
 h��UEV��!t�d:\event?_user\�u�#C7z���jpF��n��SPs�x�spo�tweld��!�C6��������! ���G|'��5k Y�����> ���1�Ug ���/��	/^/ M/�/-/?/�/c/�/�/ �/�/$?�/H?�/:J��W�3�����8C?�?�? �?�?�?�? O+OOOOaO<O�O�O rO�O�O�O�O_�O'_ 9__]_o_J_�_�_�_��$VALD_C�PC 2�« ��_�_�  w��qd�R�*o_oqo��
hsNbd�j�`��i �da{�oav�_�ooo 3BoWi{�o�o�o �o��o�PA� 0�e�w������ ����(�=�L�a� s�
�������ʏ��� ��$�ޟH�:�o��� ������ڟ؟�����  �2�G�V�k�}����� ��¯ԯ�����.� �R�S�yϋϚ����� �����	��*�<�Q� `�u߇ߖϨϺ����� ����&�8�M�\�q� ���߶���n����� �"�4�F�[�j���� ������������! 0�B�Wf�{���� �������,> teT����� ��/+/:La/ p�/�/./���� �//'?6/H/?l/^? �?�?�/�/�/�/�/? #O�?D?V?kOz?�O�O �?�?�?�?�?_O1_ @ORO9_vOw_�_�_�O �O�O_�__-o<_N_ `_uo�_�o�o�_�_�_ �_o&o;Jo\oq �o����o�o�o�  �"7�FXj�� ���������!� 0�E�T�f�{������� ßҏ����
�,�A� P�b�����x�����Ο �����(�*�O�^� p���������R�ܯ�  ��Ϳ6�K�Z�l�&� ���Ϸ���ؿ���"�  �2�G���h�zϏߞ� ����������
��1� @�U�d�v�]�ߛ��� �������,��<�Q� `�r���������� ����&�;J�_n� ������������ �$F[j|� ������ 0E/Ti/x��/� �/�/�/�//,/.? P/e?t/�/�/�?�?�? �?�/??(?:?L?NO sO�?�?�O�?�O�OvO  OO$O6O�OZOo_~O �OJ_�O�_�_�_�O_� _F_D_V[�$VA�RS_CONFI�G ��Pxa�  FP�]S�\lCMR_�GRP 2�xk� ha	`�` � %1: SC�130EF2 *H�o�`]T�VU�P�h�`�5_Pa?��  A@%pp*`�NVn No9xC VXdv��a��<u�A�%p�q�_R���_R B���#�_Q'��H�� l�;���{�����؏Ï Տ�e��D�/�A�z��-�����ddIA_W�ORK �xe�ܐ�Pf,		�Qxe���G�P ����YǑRTSY�NCSET  �xi�xa-�WINU�RL ?=�`�����������ȯگ�SIONTMO�U9�]Sd� ���_CFG ��S۳�S۵P��` FR:�\��\DATA\�� �� M�C3�LOG@�  � UD13�EX�d�_Q' B@ ����x�e_ſ�x�ɿ�VW �� n6  ����VV��l�q  =���?�]T<��y�Y�TRAIN؎��N� 
gp?�CȞ��TK���b�xk (g����� _���������U�C� y�g߁ߋߝ߯����߮�_GE��xk�`_P�
�P�R���RE��xe*�`h�LEX�xl`1�-e�VMPHA�SE  xec��ecRTD_FILTER 2�xk �u�0��� �0�B�T�f�x����� VW�������� $�6HZl_iSHI�FTMENU 1��xk
 <�\%�������� ��=&sJ\ �������'/��	LIVE/�SNA�c%vs�fliv��9/���� 7�U�`\"menur/w//�/�/������]��MO���y��5`h`ZD�4�V�_Q<��0���$WAITDIN�END��a2p6OK  �i�<���?�S�?�9TIM�����<Gw?M�?*K��?
J�?
J�?�8RELE��:G6p3���r1_ACTO 9Hܑ��8_<� �ԙ��%�/:_af�BRDI�S�`�N�$XV�R��y��$Z�ABC�b1�S;S ,��j�I�2B_�ZmI1�@VSPT ��y��eG�
�*�/o�*!o7o�W�DCSCHG �ԛ(��P\g@��PIPL2�S?�i��o�o�o�ZMPC?F_G 1��ii��0'¯S;Ms�S�4�i��p'��g���e2��  >6��N?y�I���!c?I������8?�#?�ߎ�TS��G��D<ŞB��Q_DFI�1��q>��R>15����s?	z�Q��*V?R�������?�Z�~���Ï��>�C�@���B�I�ڏ�ӈ�����*�@�N�x��$�6�H�6N�`��T�p���o�_CY�LIND�� {� Х� ,(  *=�N�G�:�w�^����� ��ѯ��� 7����<�#�5�r��� ��������޿y�_�� ��8�ύ�nπ�㜻�9� wQ �5�� ���S�����(�ٻϴX�זr�A��S�PHERE 2���ҿ��"ϧ����� �P�c�>�P�̿t�� �ߪ�����'��� ]�o�L���p�W�i���`���������PZZ�F �6