��   �A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG����DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !�� FT� @�� LOG_8	,C�MO>$DNL�D_FILTER��SUBDIRC�APC��8 .� 4� H{AD_DRTYP�H �NGTH�����z +LSq �D $ROBO�TIG �PEER��� MASK�M�RU~OMGDE�V��PINFO�.   $�$$TI ���RCM+T A$( /�QSIZ�!S� �TATUS_%$�MAILSERV~ $PLAN� �<$LIN<�$CLU��<${TO�P$CC�&sFR�&YJEC|!}Z%ENB � �ALAR:!B�TQP,�#,V8 S��_$VAR�)M��ON�&���&APPL�&PA� �%��''POR�Y#_�!�"�ALERT�&i2U�RL }Z3A�TTAC��0ER�R_THROU3UaS�9H!�8� CH- �c%�4MAX?WS�_|1��1MO	D��1I�  �1o �(�1PWD  Ɵ LA��0�ND��1TRYFDEL�A-C�0G'AERS�I��1Q'ROBIC�LK_HM 0Q'� X�ML+ 3SGFReMU3T� !OUU3f G_�-COP1�F33�AQ'C[2�%�B_AU�� 9 R�!�UPDb&PCO�U{!�CFO 3 
$V*W�@�c%ACC_HYQSN}A�UMMY1oW�2"$DM* �$DIS��SN,,	3 �	o!��"%"_WI�CT?Z_INDE�3�PgOFF� ~UR�Y�D��S�  
o t Z!RT�0�N�(cD�)bHOUU#E%A/fVa>fVa�MfLOCA� #{$NS0H_HE����@I�/  �d�PARPH&�_7IPF�W_* O2�F�PQFAsD90�VHO_� 5R42�PS�a?�TEL�� P��\�90WORAXQE� LVO#�FS1�ICE�[p� ��$�c  �S��zq��
��
op��PS�Axw_  XK�qIz0�ALw�q'0 �x
���F�����p�r��u�$� 2�{���r#����� �}��!�qi�����$� _FLTR � �y�p ��
������}�$�}y2}��bSHAR� +1�y Pe���t
�G�6�k�.��� R���v�������П 1���U��y�<���`� r�ӯ�������ޯ?� ��u�8���\����� ῤ�ڿ��;���_� "σ�FϏ�jϸ��Ϡ� ���%���I��m�0� Bߣ�f��ߊ��߮�� ����E��i�,��P� ��t���������/�l��z _LUA1��_x!1.j�08����i�1z���25c5.��q�����uh�2o��������������3����^ 1C��4_��� ������5���N �!3��6O��@�u������Q�J�MA��M?A�P�(�� Q� '��<a/�/�/{/�/�/ �/�/?&?��P?V? h?z?9?�?�?�?�?�?�?
OO��?���u�fOQL
ZDT ?Status�?uO�O�O�O��}iR�Connect:� irc�D//alert�N&_8_J_ \_�G�O�_�_�_�_�_��_���sP 2�q���_o1oCoUogoyo �o�o�o�o�o�o�o�s�$$c962b3�7a-1ac0-�eb2a-f1c�7-8c6eb5�6401a8  (y_J�On���R���ـP(�X"��rZJ�p [D�rcE\!)�,$e"�ـ[� �M�4�q�X�~����� ˏ�����%��I��0�B��f���������w�W�8 DM_�=!W�G�SNT-P�	�%��-��������x�����4#��USTOOM 
�F���W  �3$TCP+IP��XHO%,S"��ELO�W�T!=�E�H!Tb����rj3_t�pdQO \��!KCL������>�v!CRTY�G����O"(�!CO�NS�� ��ib�_smon����