��   F�A��*SYST�EM*��V9.4�0107 7/�23/2021 A 
  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTT��&F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STSTOP�_TPCHG �V LOG_P NT��N�  6 C�OUNT_DOW�N�$ENB_�PCMPWD� �$DV_� IN�� $C� CR5E��A RM9� =T9DIAG9(|�LVCHK >FULLM/��YXT�CNTD��MENU�A�UTO+�FG_wDSP�RLS��U�BURYBA�N��GI�eE�NC/  ~CRYPTE� T  �$$�CL(   �S��[!��	��	P �V� IONX(�M XKl!IR�TUA� Z/�$D�CS_COD?����_%�  W�'_� �/�(S  J�*�� � 6�A�91�"�!	 $b!��0=<? R?`?v?�?�?�?�?�? �?�?OO*O8ONO\O�rO��3SUP� �:�tO�O3F�O�O�O��  !%\"Q��6_ ��� V�[t&W��j��T�O �_��LWJ_��M �V�_��KLUGH 1��) M  9o)o;oMo_oqo�o �o�o�o�o�o�o7o /ASew�� ������+� =�O�a�s��������� ͏ߏ� ��'�9�K� ]�o���������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� 
�
�1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�q߃ߕߧ߹��� ������"�7�I�[� m����������� ����3�E�W�i�{� �������������� ,�ASew�� �����5