��  	vy�A��*SYST�EM*��V9.4�0107 7/�23/2021 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�>#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO"  � A�LM�"ENB���&ON�!� MDG�/ 0 $DEBUG1A�"d
�$3AO� ."��!�_IF� � $ENABL@QC#� P dC#U5K�!MA�B �"��
� OG�f 0COURR_D1P $Q3GLIN@S1I4$C$�AUSO4i OD��"$SEV_AN�D_NOA�#PP�INFOEQ/ �L �0?1�5/_ H �79�EQUIP 2��0NAM� ���2_OVR�$VERSI� �!PCOUPLE, �  $�!PPV1CES0�24G � "PR0�2	� � $SOF�T�T_ID�2TOTAL_EQ� �Q1}@NO�BU SPI_IN�0^�E�X�3CREEN_��43BSIG@�3OEKw@PK_F�I0	$TH{KY�GPANE�D� � DUMMYE1dT�!#U4 Q�!RG1R�
 � $TIT1 d ��� WTdWT� WTT7PWT5UV6UV7UV8UV9UW0UW^WQ�WUrW6QWU�W1�W1*�W1�W1�W2�R!�SBN_CF�!-�0$!J� ; |
2�1_CMNT�$FLAGS]n�CHE"$nb�_OPTB � E�LLSETUP o `�0HO@� PRZ1%�cMA�CRO�bREPR�hD0D+�@��b{��eHM MN�B�
1 UTOB U~�0 9�DEVICTSTI�0�� p@13�p�Bqdf"VAL�#I?SP_UNI�Cp�_DO2v7iyFR_F�@K%D13�[A<�c�C_WA_t�a^�zOFF_#@N�DEL�xLF03q�1�q%r?-q�p�C#?�>`�A�E�C#�s&�ATB�t�cW{4c{� $DB<0�"� S�("{&?��o \� VERq�$F�!��d�_�����dTMP1_5F��2��1_Rs���Rr�MO� �sE � [A��q�����REV�BIL~���AXI� ~�R  � �OD�`(�O
2`M�" �6�/�"3�� A�l�K���@D4d p �E RD_E �7��$FSSB�&w`K�BD_S��VqAG*� G�2 "_��2ϑ� V�t:5?`��qC� �a_EDu �O � C2��`�S�p�4%$l �t'$OP�@qB�q7��_OK���0, P_�C� 7��d&�U �`LACI�!�a{�ƐȤ fqX�M�  @$Dw����@�p�_+R�� BIGALLOW� (KD2�2�@VAR�d!�A�B �BL{@S �C ,M�kp�h`S�p�z@M_O]8��w�CF4d X�0�GR$@��M1�N�FLI�n�[@UIcRE�84U�IT=$�/0_N�`S�"CF�d0Mt� �#PEED��!ʹE`j��pS`JStVҒ`�\��3Np�`
ʗELBOF� �+ŷ+�pH/0̲�3Pϲ� F�2�f���1r�r@1J1[E_y_T>!� �`��g���G�� �A0WARNM��p�d��E`ѳv`NS]T� COR-$r�FLTR��TRA�T T�`� $A�CC%q�� �rb��I�.&��RT���S���`CHGV0I��.�Ti�pA�I�9�T���a�K�� �0�"`a����HDR�2��2B�2J; �C�ѿ�3��U4��5��6��7��%8��9OB`�M���3� @� TRQBt�$Efl���C�N�_U��Y�_�OC� <� b�t���3B^q�LLEC��MULTIV4�"���A
2/�CHILDd��
1 q��@T_Qb�  4� STAY2�b�=��)2�������C�  |@A06$\����i`��d�C1TO���Ep�EXT���U��2��22�0��t�!/@V�Qb.'��B s����	� "�" 	�/%�a}����_s}���#�W�[A��U�qM�� ��" ��:NP�$ L�0�� ��pA��$J�OB ���b�ETR;IG�% d��� ���-'0|������?�_M�r& tf��FL���BNG�A��BAi ���ߑ� /1����0m��R0�aPOp����'���:�$�bq��
2J��_Rҳ�C,J��(8,J��D/5C�X)�͑���@����P*��(�`˻M?P~��ʂ�FACހ��SLEWL! % Y��t!�`�R4d)�ː����qG���@N�HANC��$LG ���aRq��x���ī�!A�p����aR�­��n46���o3P�m5RA�co3AZ�@�8찔�����`FCT��S�_1F���`�SM0�1IK�AE�0��0� ҰD�����U��!���MP�B�a@Ж��HKwAES�@N�G�1BWK�N�S XYZW�`�2l���F	_�g�C�*/  ^0I\��B���+.�STD_C��t�A#n�USTJ��U��,��PU��%�IO�"�P�_hup�q��-|�$��SQOR�shR2p�����`Of0ʢSYېG P�q�Uupx�h`�f�f�9�ڠDBPXW�ORK��.�$�SKP_�p���D�B0�TR�p / ���`��e��0+�b D�q� _C�0[bc,@gPLZc�a��t���"D��DgաcR "E�С9ʨ�ؠ�NQ�1��0�RPQPR�z�
 c�����1 ��3�A�O���L2�i2�o������ y3�o����PCF��4�o3<�E�� c5[҅aRE����b6H $C�E�1$Lhs2$p�c���0y{INEҖ�Q_D;A��ROS ��rֿ���q�s� �P��vPAU�'�RET�URN�rsBMMR��U���CR�pE�WMIP��SIGN�� ��LAL�(�@�3$P��43$P�0+ 5<���#PCW�+[�D#`ސ���t~qY�ҖGO_AW� ��܀HP��rA��PCS"���CY�7�!�15Á3�*̄2Ɗ2ԆNݐ;�x�&KS��DEVI�p� 8 P� @�R)BѓճIԇP)�;��I_BYe�C�R�T�ga�HNDG�b9� H��A.�۰��$DSBLDӟ�ՆЗP?��P��L��:0�P���FB✤�FE�q���Մ��v�
±;� '��A�ö�MCS<�А�TP����BH�0W��%�E����@� ��SLA�0� <  p�IN�P�R������I�=/` ,��S0 P�6�J��x�FI0R�x��\%WQ�rWQW*�NTV�3r�V<��SKI�3TEL�v��j��ӄA�J�CjC_p��SA�F�¤�_SV�EOXCLU��}�� %D�PL��ϳY&������HI_V:@�BPPLY<`����}�����_ML+ }�$�VRFY_c��M�d�IOC��C_�&@��\���O7� �LQS�@}Bvd4\a��Ճk��PP�U�·�6S�AU��NF{F���Յ����+dQCHD`Q��D᮳`�AFSCP���T_�V�B_VALi2n�͢�'@ߑ ><p�PT8P��@|P �RG�9N���� ?��j �Tp��1 ���ɒ_�SGNԡ@�
$ ��"��q�@������ �R�دR��ANNUNp����Յ�$~P/�����&@
�&�bEF�PIqA @��F��.T�OT%�9�vd_�vd��h��b M��NI�b!B���y'��A桲��DAYmSLOAD�-�kd��wc5sa��EFF_AXIђ%C<paaCO���c�`_RTRQԡD� D��Yp� Q�BB(�E��1��� C�@p;?@�.���A� �ԡEp����p�Lt�jDU%�j��R�CABԡFP�2pNYS��IDBW�#hl��1� V-�V_l� � �DI��DG� 1$1��+T"�(!� w�"
_���!E_���VE6 @SWY�!  ��{�N�D��3OH-���PPY ��IRIQ�B�P��� �q'��A ��C�0 �0�-���N�F�@𼳀 RQDW�MS�@AX�G��LIFE`(�F}aRNY�b�W�h� ��Cr@���NT�Y0P�qFLA�Y4�OV;@nHE|��2SUPPO�P|AR`_��ՑC_XhC����Z�W�rA� C�"�BcXZ�0�a3Y2U(EC�pT�P�p!NG�T�JA �_�0��A��10�DH `�CACH��)ѽ#SIZ��ٲ-��@�SUFFI�@�`đkd��wc6b� �PM�@�$I 8��KEYIMAG�sTM|q�3;1�66����qLROCVIE$c �aJ�B�0LK��Ж�?��BD'@�$K�$�j�STw�! �2_��4\`�4��4��>�0EMAIL���p�(����FAULb�bL�B�s�SAX���UP�TTWpԡMO< $C=�Sl�v��IT��BUF�'���'�<P2P�BBD=�C���BIS$@SAV�EOB8 t"B�m �G�P�P�D=�Zp�d��_B@sE-��HOT�r{���P:�d`Z�W�WAXmSC�E�XXB@���C_GY
�P�YN_���N <���D8�)`���M����T��F�p�$�p��DI(��E�`WpX��aO���GcA^�&�Ӕq�Q1��G�F�� P (>pSV��r�kdw�p�p������aQ�dp��Q
C�CC_�p�pK �t:`��5d��R314e��8�QDSPK6bPC{kIM�Crc�a	��Q UOg��u*��0�IPL�c�� qdT!Hs  �eb��T�qrcsHS�STcBSCY�� ��Vޠ"z p9S(t,n��NVԱGQs(tHs ofB@FY1�dTc�P7Q�qSC.�*c�MER���aFBC�MP��`ET�� �R)2FU�DU`6@��J"�CDhi��`P�3�PO��3S$�� qgQ� u-уMS���z��-��u6_���AK�T�� "��O2�T�$ZO�P����U��Ė�P=���CN����������GRO�U������S� �MN����������X/�����HR�b�8{��0�PCYC���`}���s�±��DE��3_D�"��RO���� ��#���|�i����d� ����E�r��.��3M!7 �8�ALV K�U��Qj��P��B,�_3ER�TL �"�V ,�P�.gQL�0r1U 
�0l0NiO����W�0$ǤH��Ǥ��Pf�ɢC��֥j�1�`�ģP���XH *֡L ��3y���v$���w� I�'�G���G���G���G�1G�7D�8D�9PD�YF�P�1]�1j�U1w�1��1��1��U1��1��2ƺ2P��]�2j�2w�2��2���2��2��2��3Jƺ3P�3]�j�3w�U3��3��3��3���3��4Ʋ\QEXT��YlR�8qP��qP��u|P��U�AFDR�ZT"@VE���QR�� rRREr��F\�2OVMKcz��A��TROV�ٳDT�@�MX.�I�N�ٚ���IND�=�?�
i�PZPoPG@BQ�(���bHD,��(�RIV�p�2G�EARKaIO?K�҄�N�P��F�=��W0��2Z_MCM�M R �F�UR��r[��ՠeA?� ���?;�X�?;�E��C� #��OA�p��\05P*Q RI�5���OCETUP2_ g] w�NCTD�`� LET�S����������BACfR^� T�0OB�T)�Z%��p+bl�=�IFI�{�l M0��p��PyTe�!FLUI�4�_ �͑y7@UR�xA��B�Q pE@N�EMP��XR$w]S+ ?x� J����@�CVRTs��0x/$SHOxL>D0ASSp
Q��`��BG_P�����j���w����FORC� B_4f�`�2F%U&�1�R)2�RP��5s Aa |y�N�AVt��w �����S�2�$VI�SI���RSCTS�Ea�� P�BVӐO�|�$w����w��$��I���@��FMR2��b ��������P� ��������������_����LIMI�T_���tC_LM������DGCLFlt��DY�(LDS�b��5����MA��5c@B) T��FS�@�d P���2�SZP$EX_158116Pnp�qj13W;5W6�G<q���e �y��rSW�vEON9P%�EBU1G��1��GR�|`mU�sBK��O1�7 1 PO& �9P�0�p�5�0M��O%�։�SM��E�BX[�2�[���_E �f �p���TE�RM'Eg0E�OR�I�Q,@hIF�PSM2�O��,@iIF�h�zoHj{G_�UP� k� -Z�F��fw >C�@g�yG�J� ELTOL���PWpFI?��Q&��1�pUD�Dh$UFR��$ʠ�APL�u] OT&WWpT����8SNST��PA�T�aLTPTHJ��q�pE���Sv��AART~ �E� ~ FR�B�REL�Z��SHF�T�b�ATQ�X_� R(�p�smF x@$�G�P�j}!�� �����PI�Pz$U�rZ�$PA�YLO�`��DYN_8 d�TQIޥ�`ERVO�am�Xs� 4W���RP� ze�� �RCc�ޥASYM�FLTRޥ�AWJ�Gs�o�Es�~Q�im�qU�d��/a�U� nfUP[p9c[q�VOR2��M�P�GRA��l$�2�6SPP���9H���m �:R,��OC�A�1��$OP��1�����Ѱ �RE��pR�C��.�7�TSe] RRU�u�x�Q��e$PWR��,��R`R_�swTy2��C�UDs�� lqR ]n��$H��!a��ADDR��HAG`VRz�o�h�q�RR�o H��SSC �P����ç�j���w��SE1�"@HSC�D_MN<p���p�ҽ��pAaHO�LL����p�Մ֣�C�ROH�A\ND_�C�ɢNa-�#pGR'OUP[3`r_H�Y�0aq1C���}�Q��� P����ш�j���w������A���k2SAGVED������탞��q $n��p_!Dx��0��PZ�Y}�HTTP_ɠ�H��r (ԠOB�J�h���$s�L�EESG�#�s �� ��f ��_j�T�C��S`pcGKR�L�HITCOU���1�L��p���`s��p�pSSn����JQUERY_�FLA=��`_WE�BSOC��HW����A�1t��4�IONCPUk2yOZ� ��.�3s���r�˄r�~��IOLN��u 8��R��t�$SL6r$INoPUT_�$�pb��P�>��SL��
�1v���������c�˵�b��IO(�F�_AS2w��$!L� o����Q�)���AP ���0��!`HY���x�Q� +�U;OP5x `=����s�M�h�M�o����pP c�p����o�����hA�IP_ME�=y X=�IPo�k2�C_NW�l2+�y1�r0��7֞��SP��A��
� BGk1�|M�|a=z l=0cTiA7bv�AnpTI��`�e� & �՞PPS��BU& ID0Ѣnp����p��M�p���FP�{���Ԗ�ɰN��& ��IRCA�_CN-� | �č���CY��EA`�W�\��ct��r;��b��qDAYy_����NTVAL��и��rU�Ӹ�SCA1`��CL�!�ѹ��ҏ@�}���sR,)�3�N_�pC5��Ҧ�y�~�v�h���j�����,��� ?2} o����@����j���LA�BFQ��& ��UNIr��X@ITY��q�s�QAIR�@� 3����T R_URLn[�$A�EN�0кy:�=�T,�T_}UrABKY_��RDIS��� ���JY�@��$$l�eJ	 Y�R�ō "d A�4�J��#FL@0I ��
��#�
�UJR�� ���FH0�W� W��] �J7a�tJ8B7u0��(7���	8?APHI�� Q\D20J�7J8�buL_K�E��  �K���LM� � �<�XR0�g�O�WATCH_VA�qx<`f�FIEL'�be�yi@�5� � b<QV)��`�CT ��1�@�LG߅� $I�LG_SIZ���0>%� X=&4�=&FDH(I<( S(�1J&;()@U'G(:  �sC#�&� �&4��&j @�&)@�&�a�5�@_0P_CM*S1G0:1AF�a 7:4: �t(9!�RE!_6R _64�_6j k7I^8u8�0`_6)@w7i8: RS��cP  Y3ZIPD9U��P�LNFr����ӠDED1E@��[*0�A`pLCnBDAU-EEA8�0���tCB9@GH�rl��@�BOO���g� CW��IT��wDs�S�REwЎHS#CRG0��X�D퐎�>o�MARGI��TЀ�LضKât�Bڤ@�S�{�?�W�D@�DK�J{GM"WMNCH;&@�FN�%VKKW9 �IYUFWX�PWXFW�DWXHL�YSTP�WZVWX��WX~@WXRES�YHps[H�C(t@�S�bK���G"iU/��kT�G�3U `�^RG;YV�PObg�Z�E�S�2ATc�YYEXG�TUIIUI� N�S��!@{��cS�cGP��� ^5��Fp�AN(�=��ANA@q��AIp@.���DCS��P��]s��]rOcxOow�SI�rzxS�x�HIGNS ��e#HQ w�nftDEV gLL�#eA��& ����Ta2$I'��b�M䴛�SAW�����m��:�S1
U�2U�3U��b^p�& � ���R�8t ʵ�E˴����}`�F�(��ST��RD@Y�	�� �$E��C�.���8!�c%!� LT�f� � {�<�߃��[�.�8��u���6��C_ � "�_ >���@ޣ� �MC�2�{ ���CLDP��>TRQLI��יŔFLh�����b��D���E�LD�����ORG��Q�~8RESERVu��X���X���
���� � 	��UԔL��� PTא�	<������RCLMC�ȤX�j�ک�����M�U /� ��$DEBUGMASi�(����2U�DTCp���E)+��MF�RQ��� � �.)HRS_RU���m�j�Ax�/eFgREQD0�A$P<'OVER��e#2�t���P`QEFI��%R�k�+���f���Ǒ \w ��($9U��h�?����SPST�� 	��CL@�ɣ��%�ڣU �0��?(t��pMISC��� dA��RQ��	U�TB�@�� 1���a��AX�|�ǵ�EXCES.�3�o�Mv�� ���t�o�SC�� O� He��_����ȋ�!۳�����M�K���@1�B�_ FLICM�B��@QUIREcM�O�O����?��MLo�M� @���A��"m�Ȣ GMNDA��eЗB�]/(�D*3[IN�AUT�A[RSM] %�pN��!!c�Ѽ����PSTLᘻ 4�LOC��R�I��EX��ANqG9r9�}�ODAh���|���� �MF"q%ʶ��n��`x�8���0/�SUP����FX� IGG�A � ���n��!Q� n�fn����@�� P��_�@�c;��%�3TI�N�����IN�� t��MD��IMA)��cp���ߡ��H����DIAD�� W�A��;�T�a��DKC)�O�ܲ eМ ��CU�S V ��9�<�A_�� �����L����u �P�h�P� P�KEb�T3-$BF0zH��ND2ᢹ�2_{TXw�XTRAcs4����LOE@e�1������2�N91��MR�R2sŠ 1�))AA�� d$OCALI���%GQq�u2�� �Q�RINQ1y<$R�SW0���wABC��D_J� ���9���_J3�
��1SP��) 9�P��-3-SD�9�B@%J�P%y��!O�qyI�Y�CSKP暐$&0Js$J6X�Q�,�%�%�%�'��_A1Z��L!�!EL�qK"�OCMP��Y���@RTP�3+1�M ��1�/8p=:Z;4SMG�P���;JG��SCL����SPH_�pX��0�3� 9��RTER$�y!pv_Pp�����A�@ڃX��4D�I�!n223U�"DgF  ���0LW�87VELבINv��`
@_BLcp9�D� ��DG0G(E� �N �ECH��TSAy_��0�IN�0���h�N�E�B9��tAA�__� ��E �B�5�Dң�I�6F��DH��g�D��$V�$�|3qa$Z0�����$�Q���RAh�H? �$BEL� x���1_ACCEA �PX�_PIRC_4�0|�K�NT�O$PS��ʒL�0���Tߓ�@uW��Rp@vV�UY�WkS�W3�R_���_R�R�Pa���C�UQ_MG��DDa�2��FW����[S�;ekSVR0hDEYkPoPABN�WRO�0EEbV��oא�!V����VQ{A$USE�_�sP/�CTR�tY{`1P�� G�YNr�A� �fo ���a!ME�YHr`O@�QtINC3��Xb?dp��8w���ENC�0�L��9QVR�ďPI�NʂI�Ru��l4N�TC)ENT23_�2���sLO�0���p��I��#��v�0#�/���0��du.�C�@�vMOSI$aG�f a���X�PERCH  �s���2 ,���7�w� �r�w�7 2�e�P`m#A�R��L�dm#B��l'�u��zˆ�vTRK�5]�AY-��� ���R
�����6!�Fr�MOM5���N�S "�Wcu��S�b�_DU��RS_BCKLSH_C�R ��E�����c8ì�_r��� q�%CLALM��tK�<��@�CHK�� ���GLRTY@{��t��@���_��N �_UM>�;�C>�p-aw1S���LMT �_LP�#l���w�E q�����p��U���X" 0D���Ӥp�PC=�p��H��#e;�CMC�	-`1gCN_�N�2�X#SFCQa�V �b��uw�1��Rv��7CATB�SH�� 1dgv,�v�vv*�Q*�00 `PAB�6r_PA�%�_� w0� ��!�$��JG�������0OG%��2TORQU�`%�s�g`p�0��1g`��_WT����91 Q��S��S��I*��I��ISF�����W"��f!)`VCUP0>�U��1#�!`7��!)�JRK#�h�[�G KDBu0MG M"��_DLQ��GRV��ħ�S��S��H_p0���P��COS��0��LNj��&�� P�Z0���C�1���b��Z ����MY��������ۢ�THE{T0�uNK23S���S�CB��CBSC�AS������0�S���SBS"�N��GTS�!�aC!���37�C7X�@�$DU���}�E���(EQl�_磿�NE
�$�QK"�9�8�@��A�����������чLPH����u��S &�>1�>@���O�h(R
o���VVP�'V6
VCVQV�_VmV{V�	H�(.&��ECH�QH_HmH{H*�	O OO�%UO6
OCOQO_UOmO{Oo�F�����M)1�R$SPBALANCE_��}#LE9�H_��S�P�A"�"1�"@�PFULC�(�"�'�"�@�J1�!1UTOy_��T1T29QR2N��\R�p14j1@5�� ��RLSP�T���O�@^Q��INSE9G\R�qREVV6�pΎqDIF具I1�l�7�B1��pOB�1ؑ��b�2s��p����?LCHWAR{b�bAB��d�bC�p��(qdEV�X�P��'F8���B0� 
(B���JQwuROB �CR��RjE�	
�C�HQ_�T � �x $WEIGHp��$ �C'��Iq�pIF�a9`LAG�bբS�b�0�b7BIL�EOD>��p&�BSTbP�BP�1ؐB�@�/P���A�@��@�
[pHR�a�  2y��t�FDEBU�C�L�PR|�MMY�9�U�0N޳kT��3$D�QG�$UP"����  �D�O_�PA�A� <@�@%V0���a��B�B�@N�s�X_�p�`S�O� �� E%Z�T~p�qY�T�1<MT�PTICK�C�0�T1�P%c��&`N � 0�S �R���a�2�8e�2De�PPROM�PsE�� $IRi��a�b���b�MAI��@�r�e_��@�c�0�	pRn��COD*SFU�`�FID_?��e0yb~� G_SUFF��G �C�a�a3b�DO;gv0<e�@;fGR�C�2tYc$t�2/u@�2;u��t�T4P��@�H�0_FI)Q9n�sORD�A �@�]R36���r�a�P�$ZDT�e  |Q�U�4 *�1L_NA�Q&`�r8eDEF_I�x�r^f �De�B7fT7f0�De>�^fIS��j��Q���7dw�Dc�}�[T4;�͢RD0����*S�Df�O� �RLOCKEޱs8oJo\gy�rpUMu�rt0� t>�t��$r�#u� $tN�$rVy�y�/s�0 �/u�r/u0�/s����x�PP�0g��Ps���PW������@��TE㑠T�( }�ALOMB_��-�0�BVIS��I�TY�BA"�O�CA�_FRI3U��0SIs�W��R#`~�.`R~�3CS�BWZ�Wf�Ș�\�l�_ɩ9qEAS�C9r3�T�ð���b��4|�5|�6�CORMULA_Iޱ��THR�B �EG�w��@��S\8cUCOEFF_O
a�m0��
aA�G���CS��@|RCA� �_�S$����C��QGR�� � � $�4D2�RX�PTM���`�b����SER�0qT؄�t�p�  �"�LL:t��S��_SAV��f�C���p�u��U��p� �SE;TUs�MEA�`�`�л@Q�r�@� �3 ̰[@ eP>�@������ǁ���r&`$ǁ�Ą����Dr�da������ۢ�:�0�`REC�q��=�MSK_� ��� P�A1_USER-1�2l��0q�l�-1VEL�l��0Ȕ҈��1I�p�0�M�T�QCFGbѰ � (`�0OBNGORE�@�P����0~��� 4 ��8G�BAXYZ�s�1�>0HS@���_ERR�A� � 8��Q�`A��/�0QXХ��PBUFINDX���p>0MORള H�@CU/��QA}��a�q�Ӑ2�q�$J@��M�� �*��GⲴ � $SI9����`�y1p�VO���t@O�BJE� ��ADJ1U�R����AY�?E��D�OU�p�}�\�a�r=|�T_0pL���K��RDIRP��X�0� x2g@DYNH������T0��R\���P�@���OPWO�RKbѵ,�PS�YSBU� �SO!P��R�B���U���01P�PAo���X	B�OP-pU�1����1'RdQ8�IM�AGB��@D RIM��^INɠ/]?RGOVRD����p�:P< \g@�0��(���BL�B,��0>��PMC_E�pR�YQN�M�dQ]R1�bR��SL� cж� � $OVSuL�6S�DEX��DL�2Be0��_�  6_p� 6_p@UP]RuCX@�p�5�R^� _ZER����$GA��Îbѷ @�С1EO&�`RI��B@
��`x�!�����1*��LbѸx�T@
P�ATUS��sQC_Tta�>#B��H&1!��ĝ�cQ#�pcй !D�Q8 �<!L��0B`<!�q]BѳXEB  �Ŗ"�"u$����@�A UPԏ�m�PX��`h&5[T3�q"��PG�ջ��$SUB0!1E[�0!#JMPWAIT� EH5LOW�a�RCVF�a)`BK1�Ri���$CCC�R���b�7IGNR_{PL#DBTB
PPq�ABW�`�4�ЙU�P�5IGh`I�CTNLN�6�2Rȩ�肰�Nh`PE�ED� 'HADO!W
P�����E&<D�51�SPDbѼ L�@AE �\@�jCUN�@;h@�!R�� �LY�p�0:!��QPH_PK�ս~��RETRIE#���<�гA�`FI��Ҿ ��p�@�D �2���DBGL�V�3LOGSIZ,�㩁KTh1U^�!T�D'C�0_T���MB9�CAѐGP0]RAS|���CHECK�0N��P��_A�6���It�LE�!�P�AրT�B�"�0I�P�2_A� h $ARR�b� �sK����O<p�7�ATT ���2K�VGP�¥��SƎCUX����PL��`��� $���S�WITCHC2��W���AS!� AdL�LB_A�� �$BAI�D���BCAM�y�i!�`#J5�Ѷb6�fka_KNOW�S�b���U�AD�h��g@D�o��iPAYLOA����s_b�w��w�ZsL[�A��<�L�CL_�� !@��Vr�a��ct�qvF{yC:�Qz��Tti��IQxR<�QwN�mtBdꠝ�J��q_J[q:����ANDM�(�x�t[roq���ա�PLz`AL_ ��O`g@��a�:�C��DsE��J3��"�� T�PPDcCK� ���CO���_ALPH2�x�BaE��&�2�D�����|�1�  � �@�D_1z2DtD��AR�!�����^��TIA4 �5 �6�MOM��,�L��9�L�F���B_0AD�,�p�9�p�F�PUB��RQ���9���F������"���`@�  ��PM>r� ��Bb_��� e$PI�Aуx�wP�~9y�I!�I/�I=�ݔ&n��!n�	1���n���u�� CHIG^c C`5YD��YD `5�0i��ƨ�1թ<�1`5SAMP� ���)���*�`5�`�s $�X���&��g��  q�Y@　��Ҳ��)�o��h�H�0q�IN������ۻ��`2����ش�!�GAM�M��SD!�ETȤ�^�D����
$N%�IBR�!BI�$HI�_yb����E���A������LW��������ֱ�л����0$�C�5CHyK� � g�I_�����Ј����k�d��䎖j�"� ��$T� 1�ĵ�I RCH_5D�1�0RNF'C��LEh���ػ�����@MSWFLܐ4̑SCR�(100NPg�3(RL掷���,���`�Y@o�PI�3A�METHO�����5��AX#� X#@��BERI���)�3U�R|@�u	D͡��FF�*�n�
�}����L��*�,�OOPn���B�}���'APP�F� �P0F�g�R���RT��!�O�Y@՘�"�ޔ�1��ޔ~��=�6��RA�PMGAŐ� �SV���P�*PCUR2�GRyO&@�S_SA�aX�$�#NO��C� �"��$ t�Ϗ%7C���
�i��bq���DOXAAq�SQh�b꛵ ���Q���Q�"��Zs �R3���� 7� p�YL��q
����S�r%�(Rt@:�>`s�Ԁ�q_��9C�є!M_WS �!2���.�M�0�vp�!�m4;�CA:���"�M��� ���Al��!W4 �$��L"aGq4 ��2"���2"��2"F��0��N��`v�Uc���X�@O����Z�%�j0���+ ���M��if x���#����ѭAt��_Ib� |e� �($ L�~69�~6F�$  %��7�6?�dan�Z1�!�b2��ͮ@Hpb4P��Q�PMON_Q}U.� � 8�P�QCOU���PQT�HN HOm)@HY�S`ES�b)@UE�@�POGd�  ��@P ��ERUNW_TO���O��N��� PprEC��{Q INDE��R�OGRA�9`�2>2�NE_NO�DrE�IT��@V@INFO�A� Qa�J�A����A�B� =(��SLEQ��Q0��P�F�OSD��T�� 4�PENA�B`"p@PTION<�S�0ERVEv�mW���@ESGCFNQԋ @@J��zB�z�R�Xn_�WQ�ѐEDIT�A� I�A � Kϑ�����E��NU�W�XAUyT@�UCOPYϑP��l��L M��N#`�'k<�PRUT� �*bN�POUC���$GwB�d��PR�GADJ�A� he�X_�I�ӷ �f� �fW�hP�h�f����`��N	�_CY�C`"/!RGNSrJU�b,�LGOI����NYQ_FRE�Q��Wǰ��?qSIZ]TJ�LA��6q�a8G�ǰ��CRE����fJ�IF/��CNA2��%}t_G��ST�ATUe0��hGMA�IL0�t��q��$DL�AST�qs�tEL;EMNQ� �K XXFEASI[Q"]� V�I��r��-(��⤰��I�@~�6r��,A�0L��]�ABDA��E�@rĠV�qu�BAS���v��µ�U⠤�9 �$����RMҐR W�����Ń�#᠑��qb�� Qr���m0�	4� 2�  糝$մ����� ������E����DO!U�C��a�tP���=�RGRID�ADCoBARS��TY\S��rOTO�0�A� cA_�t!�`�����O� KT� � �@�0POR�C铚�.�SRV�p)	��DIB T_w�#�5�P��?���?�4=�5=��6=�7=�8!�/!F�Q�NQ�a@$VA�LU����1�@F>JU�� !WUM!ĳAӓ�q��AN�Ǣ�q��Cr�TO�TAL_�t[�%�P�W,sI��:�REG#EN8�M��3X���C0,��1�@TR���r�8�_S ��M���V �a�T���Rv�E�s���.A�rB`�V_HƩ�DA3����S_�YH�"PvS' AR�02� zbIG�_SE%C����u_�v@ڴC_��$CMX\�U%f�DEW .��t�IL�Ze�?�>TF�T HANCAߊm0
WW�rSs��I#NT ��a�FlC�!�MASK�㧀OVR��@��+0�q�ѝ�OVCir�z�Q������SR��9�v����P�SLG7�ա� \  QuI�""��pqS��tx�UH� hG��γ��I�U�ar��TE� �� �(u���JQ�@`sI'L_M_t�Vc�����0TQ@���A��C��6�V=�CK�P_h�9 U�Ml�V1k�V1y�2��2y�3*��3y�4��4y��F�� +����IN�VIB E�2�T9�25�2A�35�3A�45�4A��@T� a2P� V��c����"��PL�pTOR@�IN���p�$�@�d�MC_YF2@G L	(���M� I��%�a� o02x��K�EEP_HNADED!`z�j	C�!�������ЁO A_-`Ű��ǁREM���q㒨���U�te�HPWD  `�SBM��ڐCOLLAB$蠃���r�PITp� 8bN=O1FCALW#��DON
ro��$� ,�FL] ��O$SYN �M�0�CR����UP_D�LY�A�DEL�A��q�rY�0AD�1$TABTP�_R��QSK;IP6%� ���t@aO� ��F��P_t@ �B'�@�"�`,'�Q:) �Q:)V�9*c�9*p�9*@}�9*��9*��9*9�aO�J2R�`�@�SSX��T9s�!�A��!��`\�!�A\TO��RDC���� ��PR�S��Rrq��,B���RGE�PF���j�FLG	A+��S9WjY�SPC�C�a�UM_� ��2TH�2Nd��0�  ?1� �� ��>JR � D�@��<t9~�2_PC�c�2�S��ف@pL10_�C^r  �6�� �`��9�� N5ꆀF�&�.A,4�`�Q)� =��1��eC�@�K�~�pˡ�5���0� P�0�DESIGB9�V�L1�91�6�C�G10� _DS�F�C�ھ0F2`11Q� �lQ ��ҍ XSDA�T� �do�Bw*RIND���!Q2`��!Q�R���HOMEKR �D2�B�__%_�7_I_[_ 	�D3�B�~_�_�_�_�_�_W ��D4�B��_�oo1oCoUo �
�D5�B�xo�o�o�oP�o�o��C6�B��o@+=O�g7�B�r�����aw8�B����%�7�vI� �1FPS$>�A�  ��C�b�p0C� E��� T�0���IO���!�I��G�O`_�OP-�E��o1ˠ��$��ASSp0����r�� �  �g��SI-�p��}�XK��IR�TUALo���AA�VM_WRK 2� �� �0  �5�y����� �	7�(�K�� ��!�9�v�]�{�'������6���������B�S�P1 1���? <ϯ@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0��B�T��C�AXL�M_�W��$�  di�INr���h�WPRE�0E����N��_UP<B�����~��IOCNV_�0֕� Ȁ�P��USص� �
�IO�V �1̛P $���`a�L��I��?�W� w�l~����� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ����
��.�@�R�i�LA�RMRECOV ���{��%LM_DG 5@ �Z�LM_IF 5��W����#�5πC��f�xϊϜϭ�, 
 ����Q�@]��� �2�C�$�� g�Nߋ�Jϯ����������¿NGTOL � �� 	 A�   5�G�i�PPINFO �� ��z����{�  �²���� 	���-��)�c�M���q������������� 1CUgy����ǺPPLI�CATION ?}$�����Handl�ingTool � 
V9.4�0P/17F��?
88340$sF0J7549�$+7DF5x�None��FRA� �6g�_ACT7IVE_�  �.��  �UTOM�OD���,��CHGAPONL/� /#OUPLE�D 1ܹ� �l p/�/�/�CUR�EQ 1	ܻ  UT�)�,�,	�/� 5� 4��Ξ"��$H��%o"�*HTTHKY?���/�/�/? m??�?�?�?�?�?�? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�_ �_�_�_�_�_oo+o =oOoaoso�o�o�o�o �o�o�o'9K ]o������ ���#�5�G�Y�k� }�׏����ŏ���� ��1�C�U�g�y�ӟ ������ߟ���	�� -�?�Q�c�u�ϯ���� ��ۯ����)�;� M�_�q�˿������׿ ݿ���%�7�I�[� m��ϑϣϵ�����<ư%TO��#DO?_CLEAN</��s�NM  $� �/��������	���.DSPDRYRLz��HI ��@�� u��������������)�;�M��MA�X� Z��1K'k�X�Z�jg"j�PLU�GGZ [�g#%PRUC,�B����d��V���O��5�G�SEGF3 K#.�� ��u������(LAPR�e'3# 5GYk}�������.#TOTA�L����.#USENUR _+ @�D/2�� RGDISPM+MC1 ��C9}�@@G�_$OP�r��=[#_STRIN�G 1
++
��M$ S�
~�!_ITEM1�&  n��/�/
?? .?@?R?d?v?�?�?�? �?�?�?�?OO*O<O�I/O SI�GNAL�%T�ryout Mo{de�%Inp|@�Simulate�d�!Out�L�OVERRO� �= 100�"I?n cycl�E�!�Prog Ab�or�C�!xDSt�atus�#	Heartbeat�'�MH Faul<WSAlerYOO =_O_a_s_�_�_�_�_�_�_ V��+V� �/�_0oBoTofoxo�o �o�o�o�o�o�o�,>Pbt�_WOR1 �+�q o��� �
��.�@�R�d�v� ��������Џ����*�PO�+ QP� �{9�s���������͟ ߟ���'�9�K�]��o���������ɯK�DEVS���g���-� ?�Q�c�u��������� Ͽ����)�;�M�|_�q�PALTm ���r���������� �,�>�P�b�t߆ߘ߀�߼���������GRIp��+<���d� v����������� ��*�<�N�`�r�������*�" Rm��T� ��,>Pbt ��������(:L��PREG�΅��^��� ��//*/</N/`/ r/�/�/�/�/�/�/�/~RM�$ARG_�p�D ?	����31� � 	$RF	[G8]G7�RGh9&0�SBN_CONF�IGa@3;�A�B��1�1CII_SAVE  RD�1�3�&0TCELLSE�TUP 3:%�  OME_IO�RMRL%MOV_qH�0 OOREP���QO:UTOBAC�K�139�2F�RA:\r X\Or�0'`�@rΥH� �K�0 �25/12�/01 20:2/1:02ri8r`_$_Q_H_�L��q_��_�_�_�_�_�_r� �_ o2oDoVohozoo �o�o�o�o�o�o
�o .@Rdv�������������  �A_tC_\A�TBCKCTL.TM?�W�i�{�����.fKINI���E�5��1q@MESSAG�0Ɓ�1;0ыODE�_D�0�6�5��Ox���nCPAUSd�� !�3; ,,		�i035h�v� \������������ڟ ����J�4�n�X�j�椯��;�E�TSK�  K��O��q@UgPDT��ćd���XWZD_ENqBĄ�:�STAÅ�31�%1WSM_C�FG 35��57b�GRP 2�l� F2B� s A�9XIS�0?UNT 235�1�0� 	ۯ��M1 �"��F�1�j�Uώ�pyϞ���ǴMET��2ֹ��P��߫ϼ,߿�SCRDf�1�l��@��5�2 !߅ߗߩ߻����ߞOrQ�9r�/�A�S�e� w���߭����������+�����7tAG�Rϰ	�)�j�:�NA�@2;	tDg�_�ED1l�
 ��%-@�EDT�-X�.J���LD�4@-tC��ri2�g_F���  ��t2}-K[�.� &�Xj �v3I����r� $6�Zv4/� b/��>/�/�/�/&/v5�/Q/.?u/��
?u?�/�/d?�/v6 �??�?A?��?AO�?�?0O�?v7yO�?�O O��O_TOfO�O�OBv8E_���_P��n_�_ _2_�_V_v9o�_^o�_S�:o�o`�_�_�o"ovCR| �O);�Mo�o�o�^�oj��NO_D�ELv�h�GE_U�NUSEt�f�IG�ALLOW 1���   (�*SYSTEM*��	$SERVp���)�E�REG2��$T��)�NUMxW�|�j�PMU�p>�LAY����PMPAL|J���CYC10�~�Ɏ�����ULS�U��k�˂à3�L��>�BOXORI�[�CUR_+�j��PMCNV���+�10ߎ��T4D�LI)�$�F�	*P�ROGRA1�PG_MI����AL�� ���B��)�$FLUI_RESUχW�a��{���MR@�O��| �0�ѯ�����+� =�O�a�s��������� Ϳ߿���'�9�K� ]�oρϓϥϷ���������rLAL_OU�T �S��W?D_ABORЀ��K�ITR_RTN�  rd���N�N�ONSTO��y�� �CE_RIA3_I�py��Ѕ����FCFG �����rn��_LI�M@�2�� �?  N 	P�1�}b<L�N����`��  ����rh
�p���\���PA8�G�P 1�����o�8�J�\��C�  C2���>��H���������Cf��z*��������x���\�������C�������rg?���HE�pO�NFI��X�.G_�Pq�1�  �u�x��������.KPAUSfH�1��� ߂ �>�,jPz� ������
/0/�/T/f/L/�/ P�A��y�ի�Mn�NFO� 1	��� ���/}b�/%?~b_ D��}bD��4  � 7?I;�ЍO����rgJ�COLLECT_��a	�B��ך7EN��py�`Ҷ2s1NDE�3� 	���r1�234567890
G}bC���OF�����~a)UOzOC|TO fO�OD{�O�O_�O�O �OK__(_:_�_^_p_ �_�_�_�_�_#o�_ o oko6oHoZo�o~o�o��o�o�o�6�!�;� �=�2IO #�9�1,7x�}�ء�KwTR �2$/}(��fy
�o�~9 �%Z}�z>Dy_M+OR�&� ��$ t�1t���z�����ԏPM����'[�,>A?'']0)���K1����*P��(/}�����>��ͯ=L����R��)`}?������K1A�,:5Ⱦ�x��A]0��Bː��B����@ֽ�����:d��<� <#ׁ
�1�$����IJ�3*��@�N�+[��k��d��T_DEFPROG ��%���~�SpNU�SE��/��KEY?_TBL  �����"�	
��� !"#$%&�'()*+,-.�/G:;<=>?�@ABC��GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~��������������������������������������������������������������������������������͓���������������������������������耇�������������������s��q��LCKϬ8�م�ϠSTAU�~�=X�1_ALM6�]���_AUTO_D�O����j�INDx�48Ι1R_T1t�f�T2�ϧՔӚϬ��TRL��LETE�w���_SCRE�EN ��kcsc��U��MMENU 1,�?  <���� ��,5gߑ���~#���� �����8��!�n�E� W�}���������� "����1�j�A�S��� w������������� T+=�as� �����> 'M�]o��� ���/://#/p/ G/Y/�/}/�/�/�/�/ �/$?�/?Z?1?C?i? �?y?�?�?�?�?O�? �?OVO-O?O�O|J�_MANUAL�φ��DB����DBG_ERRL��s-V�pq �O�!_3_E^�ANUM�J��~���?�DB�PXWORK 1.V�_�_�_�_�_|�_�DBTB_�G /�M��;q��uqDR�WAY�C�pqGCP ��=��>�AdS��J_�BY���Փ��H_�@ 10�{�
�_�o5���o�of_M��IS�5�Nk@*�sONT�IM������5v�i
ޥ�cMOT�NENDӯ�dRECORD 26V�� ���G�O��q���Nb�	�� -��x5�\������� ��ȏ_�u���m�"��� F�X�j�|�����ğ 3��������B��� f�՟��������/�� S��w�,�>�P�b�ѯ �������ο��� s�(ϗ�!ϻ�pςϔ� ����ϵ��� �o�p �8�J߹�n�Y�gߤ�o�MEN������]� ����H�o��Eu� �����,���P�� �)�;���_���������������L�wTO�LERENCLdB�ȕbZ`L���@C�SS_CNSTC�Y 27�Y��@���b�M[m� ������% 3EWm{��(�DEVICE 288'f�//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H?�Z?l?~?�?w+HN?DGD 98,`�Cz�:�q+LS ;2:8 �?O O,O>OPObOtO�?*�PARAM ;��i|bpe�D�5�5SL?AVE <�=�7_CFG =�O��CdMC:\�* L%04d.CSV�OePc-_�b��A ZSCHbP�1��o�Nm_�_�G��F��R�Q�_�_�_�H�`��JP�c�^�a��$m�DRC_OU�T >�=7a�O__NOCOD�@?�g��MSGN @��u�r�01-�DEC-25 20:22]P�o�c� [����i��a�N�`���s��M��Þ�,��\�EVERSION �j�V4.5.2���EFLOGIC� 1A� 	�h��ya�}srP�ROG_ENB � �U�6�sULS�E E d�Esr_�ACCLIM�v���C� �WRSTJNT�w�a�c�sqMO�|�Q�BA�I?NIT B��ev� ?�OPT�@� ?	~�W�
 ?	R575�C���74��6��7��50Ո1Ոft�y��mw>��TO  ��	tT�nvVe�DEX�w�d�b�l�PAT�H v�bA\�Z���˟��HCP_�CLNTID ?<Qv�C !k����IAG_GR�P 2G�I ��� 	 E�7� E?h D��� C� C ��B���!� U���!�}�� �����C��Cm��B�N�Bzo�OB�)�Bk��!�f383� 6789012�345��P�T�� � A��A����A�A��O�A��A�{+As�A�j�RAbJA�Y%!��3a@�bZTpZPY� A� Y ]PB4!��0�!���3a
��������Q�A����A���A����A�����hAx�~�Ao�7Af�9X~�Q�>��m@X�j�~���z�����_�AY�;A�S�TAM�^A�GdZA@�A�:bA3%A+�-A$Jz��Q���ϖ�@�;�d�ƀ��@{��@u�-@o��@i�7@cC��@\�j@V9{`�n��5?tφ����"�@_��@Z�^5@T��@O��@IG�@C�33@<��@6�+@/N�(�`@\�n�ߒ�0߶�s��nE�@h�@�b�!@\��Vf�f@P��Ihs@B��@;�t� �ߘߪ߼ߞ�H�p�� `���B���� ��� �6������~���n� ����P�����U�,����E���]���p�>8Q��0��R?� y <p�7�ŬX'Ŭ5AFd�p�@�p����@ѵ� � }@m�Ah�ZP�U�=+<���
=T��=��O�=��=��<���<�� ���^ �?�� �C�  <w(�U�R 4|9�V�)���4!�A@2b?x���j�� x��|�!�����/�@/R/��?#{�
t"�\>� ��%p���G��/G�p�8`�! �]T\Qp��8���!���$���CnB�Lo�Pq��A?/<�M'�uv?�4�?v��D�  D�  �CΟ?0<�?�? <`�?O-O�V�?PZO�?~O1;�H�H E��OgO�O�O__	_ B_-_f_Q_7�`/Z_�_�0�CT_CONF�IG H�o/c�eg�u2�ST�BF_TTS�w
@�ycHp�U�f}`�MAU'���RMS�W_CF�PI?� � q�8zOCVIE�W/`[�we{��� 	O�o�o�o�o	� �oDVhz��- ����
���@� R�d�v�������;�Џ ����*���N�`� r�������7�̟ޟ� ��&�8�ǟ\�n��� ������E�گ����X"�4��\RChcK��<b!ЯB�l�����ſി�ؿ�!dSBL�_FAULT �L_��h'�GPMS�Kg:��PTDIAOG M�Y{aD3��!aUD1�: 6789012345���R���WB�P�_������	�� -�?�Q�c�u߇ߙ߫� ��������R6��B�M�
��;��VTREC	Ppς�
�Ă��C� �Ͼ���������*� <�N�`�r����������������)�&�gU�MP_OPTIO1N`3�@TRhbc:7�aPMEeT�Y_TEMP  È�3B�"`� �A� �UNI�M`e�\fYN_B�RK N�o�fEDITORFL��_X�ENT 1�O_�  ,& ��V/D��Up� ����/�+// O/a/H/�/l/�/�/�/ �/�/?�/�/9? ?]? D?l?�?z?�?�?�?�? �?O�?5OGO.OkORO��OvOMGDI_�STA��Q��N�C_INFO 1yPok����P``�OW�C�B1Qok� ���I_<_/
/d�_�_�_�_�_ �_o!o3oEoWoio{o �o�o�o�o�o�o�o n4FXjxy�Q x������
� �.�@�R�d�v����� ����Џ����z- 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ ����%�/�A�S�e� ���������ѿ��� ��+�=�O�a�sυ� �ϩϻ��������� �9�K�]�w�mߓߥ� �����������#�5� G�Y�k�}������ �������'�1�C�U� ��ߋ����������� ��	-?Qcu �������� �);M_y��� �����//%/ 7/I/[/m//�/�/�/ �/�/�/�/!?3?E? W?q{?�?�?�?�?�? �?�?OO/OAOSOeO wO�O�O�O�O�O�O�O ?_+_=_O_i?[_�_ �_�_�_�_�_�_oo 'o9oKo]ooo�o�o�o �o�o�o�o_�o#5 Ga_s_}���� �����1�C�U� g�y���������ӏ� �o�-�?�Q�ku� ��������ϟ��� �)�;�M�_�q����� ����˯ݯW�	��%� 7�I�c�m�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� �����/�A�[�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ������������� '�9�S�I�o������� ����������#5 GYk}���� ����1�]� gy������ �	//-/?/Q/c/u/ �/�/�/�/�/��? ?)?;?U_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�/�O_!_3_M? W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�O�o +E_7as� �������� '�9�K�]�o������� ��ɏ�oՏ���#�= OY�k�}�������ş ן�����1�C�U� g�y���������ۏ� ��	��-�G�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ�3������%� ?�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������7�A�S�e� w��������������� +=Oas� ������� /�%K]o��� �����/#/5/ G/Y/k/}/�/�/�/� ��/�/?�/9C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�/�/�O�O_ _1?;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo[omoo�o�o�o �O�o�o�o)_3E Wi{����� ����/�A�S�e� w��������oя��� �!�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ����ۯ����+�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝϷ�ɯ���� ��	�#�-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E Wi{������ ���/ASe w������� //+/=/O/a/s/�/ �/��/�/�/�/? '?9?K?]?o?�?�?�? �?�?�?�?�?O#O5O�GOYOkO}O�O�/ ��$ENETMOD�E 1R5��  � ¹ �%�O�K�@OATCFG S5/�AT�B�C�UDATA �1T�I!P��A*W_*�Hu_�_�_D�_�[d�_�[1�& �_	oo-o?oQocouo �_o�o�o�o�o�o o,�oM_q�� �!3����%� 7�I���������� ǏُS� �w�!�3�E� W�i�{������ß՟�������@RPO_ST_LOPV@[��
%V_�q������ARROR_PR;��%�J%��ׯ��TABLE  �K�?�,�>�'�RSEV_NUM �B  ��A�n�1�_AUTO_?ENB  �E�C_NO�� W��K�Am�  *U�ư�ư�ư�ư�y�+Ű߿�ϟ�F�LTR����HIS�j����@��_ALMw 1X�K ���Ƽ� +ϟϱ� ���������_c���  �Kı�B>���@TCP_VER� !�J!Ư	�$�EXT:�_REQ�?�薹��SIZ\�ߋ�STK�������TOL  ���DzG��A= ��_BWD��а#���B�DI� �YWJ��A��$�S�TEP5�G�@a�O�P_DO�߶AFA�CTORY_TU�N?�d��DR_G�RP 1Z�I)�d� 	9����@���x����� �n��So �k� ���+���=�N�8�q� \������������������7"
@R�Z�@���?Ơs�?*�>
 E����[>�H8�����E7� E?�p D��� D}��Й  C���	B�  � � A@C@UU�U7UUC�>�?]�>П�| �EͰF@ F��5U�OL����M��Jk��K�v�H�,�/Hk�O?} ��%9tQv�8�?��6h�%%O�(/}�FEATUROE [5��A�Handl�ingTool �v%��Engl�ish Dict�ionary|'4�D Stk ard�v&~%Analog� I/O�'�'gle Shift�/�uto Soft�ware Upd�ate�)mati�c Backup�z)1ground� Edito |'C_amera� F�/�CnrRndIm�!3X<ommon �calib UI�S3{6n:1�0Monoitor�;trt ?Reliab� {(�DHCPo9�:at�a Acquis��3�9iagnos�1�!�;ispla�y=1Licens��1�5ocument Viewe�2��7ual Che�ck Safet�y�1&hance�d�6{*�EsS@Fr�K0}'xt. DI�O �0fiD�Ge�nd�@Err�0L(B�M�Gs�Ir� �@� �y*FCTN /Menul@v�3W�TP InPfayc3U~%GigEE^�WU30p Mask� Exc�@g�GH�TCPProxy �SvTD�Vigh-wSpe�@Skin4��U@�@mmuni�c0ons�Xur�*PP�?�!FRcon�nect 2�Xn{crEPstru�"$�Z#`eJAd@JE$�KAREL Cmod. L�Pua�X~ZcRun-Ti�@�EnvPhPel u+0s0S/W|'�5EgBSL�@Book�(System)�y*MACROs,~�R/Offse� ��eH�@0�?�`MR��0�2NMechStop�Qt`�2�ei�B�+Ovx�@� 0�~od� witc�h}#sA.v�{O�ptm�#s�Pfi�lSL"wg�W�eul�ti-T�P=3z)P?CM fun-g+��o�4gB$�K�Regei�`r�P.�riL@�F;���� Num �SelGu���@ Adju�P��Ɓ�*׍tatu��NJ~%�RDM Robo}t� scove�!�+�ea��@Fre�q Anly�WRemEp�An�'+�7�Servo�@�p{(?SNPX b�b�.;SNCPCliKA���"Libr�#Οk Q Vt����o�`t*P�ssag$�$R� 0�#�ax+R�/ID]'��MILIBP�*�P� Firm�":�P�*SAcc40<;TPsTX�?(�eln�`�m�+�s!�e;�orq}u� imula�14Q1�u�pPa�a:��30�1�s&�Pev.�'�� rid@ïU�SB port ��0iP�@aL@w�R� EVNTj�|�n?except�@l��Y�w��H�MVC�1r�R�RKxV�0����	�4���S��SC��;�gSGEP�F�UIx+?Web Pl��΀���_�ĢP~DJAVZDT Appl�T<y*��EOAT6� 4�}&����!�Gridp;�-A��iR��.�*o�AϺ"RC|P0120iC�,�larm Cau�se/j�ed�(A�scii�QłLosadS@��Upl��2r?l� �1Gu�&�2)�P0B6yc� �b0��e�q@VRA/��@��$Jain1��r{(�NRTL���#On>n e Heln8/�`E_.�}�z�`�tr�KROS Eth�a�tI�e��j�"�$6�4MB DRAM���Q�FROZ�� r_cWeld�Pcg��"tC5ell�,y=sh�����c�{��� Yp1���ty� s��A7W�R��p.�;k��A�2w-maie@ěwMh6����0qglu�pHj�CP�hR�/��L��Sup���q�� �@Pcro�6���c�x�6@�uest�#rtcA6�x*�9/� dv������ ///2/</i/`/r/ �/�/�/�/�/�/?? ?.?8?e?\?n?�?�? �?�?�?�?O�?O*O 4OaOXOjO�O�O�O�O �O�O_�O_&_0_]_ T_f_�_�_�_�_�_�_ �_�_o"o,oYoPobo �o�o�o�o�o�o�o�o (UL^�� ������ �� $�Q�H�Z���~����� ��Ə����� �M� D�V���z������� ������I�@�R� �v����������� ����E�<�N�{�r� ���������޿�
� �A�8�J�w�nπϭ� �϶���������=� 4�F�s�j�|ߩߠ߲� ��������9�0�B� o�f�x�������� �����5�,�>�k�b� t��������������� 1(:g^p� ������ - $6cZl��� �����)/ /2/ _/V/h/�/�/�/�/�/ �/�/�/%??.?[?R? d?�?�?�?�?�?�?�? �?!OO*OWONO`O�O �O�O�O�O�O�O�O_ _&_S_J_\_�_�_�_ �_�_�_�_�_oo"o OoFoXo�o|o�o�o�o �o�o�oKB T�x����� ����G�>�P�}� t���������֏��� ��C�:�L�y�p��� ������ҟܟ	� �� ?�6�H�u�l�~����� ��ίد����;�2� D�q�h�z�������ʿ Կ���
�7�.�@�m� d�vϣϚϬ������� ���3�*�<�i�`�r� �ߖߨ���������� /�&�8�e�\�n��� �����������+�"� 4�a�X�j��������� ��������'0] Tf������ ��#,YPb �������� //(/U/L/^/�/�/ �/�/�/�/�/�/?? $?Q?H?Z?�?~?�?�? �?�?�?�?OO OMO DOVO�OzO�O�O�O�O �O�O_
__I_@_R_ _v_�_�_�_�_�_�_ oooEo<oNo{oro �o�o�o�o�o�o A8Jwn�� �������=� 4�F�s�j�|�����͏ ď֏����9�0�B� o�f�x�����ɟ��ҟ������5�,�V� � H552�F�l�21r�R78�q�50r�J614�r�ATUP��54�5��6r�VCAM�r�CRIѧUIFv��28ҦNRE~��52ŦR63}�S�CHr�LIC�DwOCV2�CSU~��869��0��EI�OC�4q�R69�ŦESET��ħJ�7ħR68}�MA{SKr�PRXY�]7r�OCO��3��hq�����3ٶJ6���53U�H�LCH^��OPLG��0�MHCR¶SP�MkCS��0��55���MDSW���OP��MPR���0n��PCM�R0�ǰ����Z��51��5u1�0��PRS���69ٶFRDѦFwREQ~�MCNr�{93��SNBA�^�SHLB~�M��t���2��HTC���TMIL~�U�TP�Am�TPTX��ELq�Z�U�8����}�wJ95��TUT巻95ٶUEV��U�EC��UFRѦV�CCy�Oi�VIP���CSC�CSGt�G�Ir�WEB��7HTT��R6�#�l����CG��IG��oIPGS
�RC�ֻDG�H84��R[66��R7��RطR53�68�2��RȂ��4i�6u6E�4}�NVD���R6\�R84�Du0��F��AWSѧsLI�ȸ�CMSm��2 ��STY��TO���7T�NNٶOR�Si�J�?�OL�@END~�L��S{FVRm�M��� � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z#�  H5�52V'p!21v)R�78u,50v)J6{14v)ATUP�*�545�,6v)VC�AMv)CRI�+U�IF�+28�*NR�E�*52�*R63�+SCHv)LIC�5:DOCVv:CS]U�*869�+0�*�EIOC6;4u*R{69�*ESET�+v�+J7�+R68�*�MASKv)PRXuY<7v*OCO�<�3�,u*@�,3UJJ�6�,53�:H�LL{CH5JOPLG�+�0uJMHCR6JS��KMCS�,0K5=5�*MDSWV[dK;OPdKMPReJR0��L0�*PCM:R�0�[@�*P�K51��+51�\0�*PR�S�;69UJFRD��*FREQ�*MC�Nv*93�*SNByAF;�KSHLB�j�M�kR0E\2�*HT=C�*TMIL�,�:�TPA�:TPTXF�jELujP�;8�+ܒ �*J95%:TU�TeK95UJUEV��:UEC5JUFR��*VCC�|OZV�IPzCSC5zC�SG5:�0Iv)WE�B�*HTT�*R6�D<c|� 5�CGT�I�G4�IPGS��R�CzDGdKH84n�*R66�*R7�;�R�\R53�[68��\2uJR�L�0�\4��66�4�*NV�D�:R6[R84�uJD0��FӜAW�S�+LI�\�+CMqS�:"��*STY�kTOU�7�<NNUJORSZJ��&J3l�OL4�END�*L:�{S��FVR�9U( ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���������*� <�N�`�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�o�o �o�o�o&8J \n������ ���"�4�F�X�j� |�������ď֏��� ��0�B�T�f�x��� ������ҟ����� ,�>�P�b�t������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��� �2�D�V�h�z� �ߞ߰���������
� �.�@�R�d�v��� �����������*� <�N�`�r��������� ������&8J \n������ ��"4FXj |��������//0/B/R)^ �STDY$LANGz$u)�/�/�/ �/�/�/�/??/?A? S?e?w?�?�?�?�?�? �?�?OO+O=OOOaO sO�O�O�O�O�O�O�O __'_9_K_]_o_�_ �_�_�_�_�_�_�_o #o5oGoYoko}o�o�o �o�o�o�o�o1z�RBTy&OPTN N`r�����>�DPNx$� � �2�D�V�h�z�������Q(���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\�n���� �����������"�4� F�X�j�|��������� ������0BT fx������ �,>Pbt �������/ /(/:/L/^/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n��� ������"�4� F�X�j�|�������ď ֏�����0�B�T��f�x���������қ��՟���)�;�M��99T��$FEA�T_ADD ?	��������  	Q����� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto�t�DEMO [~��   Q� �m�o�o�o�o�o& /\Se��� ����"��+�X� O�a�{���������� ߏ���'�T�K�]� w����������۟� ��#�P�G�Y�s�}� �������ׯ��� �L�C�U�o�y����� ��ܿӿ��	��H� ?�Q�k�uϢϙϫ��� �������D�;�M� g�qߞߕߧ������� 
���@�7�I�c�m� ������������� �<�3�E�_�i����� ����������8 /A[e���� ����4+= Wa������ ��/0/'/9/S/]/ �/�/�/�/�/�/�/�/ �/,?#?5?O?Y?�?}? �?�?�?�?�?�?�?(O O1OKOUO�OyO�O�O �O�O�O�O�O$__-_ G_Q_~_u_�_�_�_�_ �_�_�_ oo)oCoMo zoqo�o�o�o�o�o�o �o%?Ivm ������� �!�;�E�r�i�{��� ����ޏՏ���� 7�A�n�e�w������� ڟџ����3�=� j�a�s�������֯ͯ ߯���/�9�f�]� o�������ҿɿۿ� ���+�5�b�Y�kϘ� �ϡ����������� '�1�^�U�gߔߋߝ� ������ ���	�#�-� Z�Q�c������� ��������)�V�M� _��������������� ��%RI[� ������� !NEW�{� ������// J/A/S/�/w/�/�/�/ �/�/�/�/??F?=? O?|?s?�?�?�?�?�? �?�?OOBO9OKOxO oO�O�O�O�O�O�O�O __>_5_G_t_k_}_ �_�_�_�_�_�_oo :o1oCopogoyo�o�o �o�o�o�o�o	6- ?lcu���� ����2�)�;�h� _�q�������ԏˏݏ ���.�%�7�d�[�m� ������Пǟٟ��� *�!�3�`�W�i����� ��̯ïկ���&�� /�\�S�e�������ȿ ��ѿ���"��+�X� O�aώυϗ��ϻ��� ������'�T�K�]� �߁ߓ��߷������� ��#�P�G�Y��}� ������������ �L�C�U���y����� ��������	H ?Q~u���� ��D;M zq������ 
///@/7/I/v/m/ /�/�/�/�/�/?�/ ?<?3?E?r?i?{?�? �?�?�?�?O�?O8O /OAOnOeOwO�O�O�O �O�O�O�O_4_+_=_ j_a_s_�_�_�_�_�_ �_�_o0o'o9ofo]o oo�o�o�o�o�o�o�o �o,#5bYk� �������(� �1�^�U�g������� ��������$��-� Z�Q�c����������� ��� ��)�V�M� _������������ݯ ���%�R�I�[��� ��������ٿ�� �!�N�E�Wτ�{ύ� �ϱ���������� J�A�S߀�w߉ߣ߭� ���������F�=��O�|�s��  ������������ !�3�E�W�i�{����� ����������/ ASew���� ���+=O as������ �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?}?�? �?�?�?�?�?�?OO 1OCOUOgOyO�O�O�O �O�O�O�O	__-_?_ Q_c_u_�_�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m �������� !�3�E�W�i�{����� ��ÏՏ�����/� A�S�e�w��������� џ�����+�=�O� a�s���������ͯ߯ ���'�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߯� ��������	��-�?� Q�c�u������� ������)�;�M�_� q��������������� %7I[m ������� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo�1oCoUogoyo�o�i  �h�a�o�o �o�o%7I[ m������ ��!�3�E�W�i�{� ������ÏՏ���� �/�A�S�e�w����� ����џ�����+� =�O�a�s��������� ͯ߯���'�9�K� ]�o���������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ��������� ��1�C�U�g�yߋ� �߯���������	�� -�?�Q�c�u���� ����������)�;� M�_�q����������� ����%7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qcu��� ������)�;� M�_�q���������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����+� =�O�a�sυϗϩϻ� ��������'�9�K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }������������ ��1�C�U�g�y��� ������������	 -?Qcu��� ����); M_q����� ��//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo�]ooo�o�o�a�` �h�o�o�o�o) ;M_q���� �����%�7�I� [�m��������Ǐُ ����!�3�E�W�i� {�������ß՟��� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9� K�]�oρϓϥϷ��� �������#�5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u����� ����������) ;M_q���� ���%7I [m����� ��/!/3/E/W/i/ {/�/�/�/�/�/�/�/ ??/?A?S?e?w?�? �?�?�?�?�?�?OO +O=OOOaOsO�O�O�O �O�O�O�O__'_9_ K_]_o_�_�_�_�_�_ �_�_�_o#o5oGoYo ko}o�o�o�o�o�o�o �o1CUgy �������	� �-�?�Q�c�u����� ����Ϗ����)� ;�M�_�q��������� ˟ݟ���%�7�I� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�s߅ߗߩ� ����������'�9��K�]�o�����$�FEAT_DEM�OIN  ����������INWDEX���ኽ��ILECOMP �\���������SET�UP2 ]����  N �@���_AP2BC�K 1^� G �)��t���%j�����������i� ����"��/X��| ��A�e� �0�Tf�� �=��s/�,/ >/�b/��/�/'/�/ K/�/�/�/?�/:?�/ G?p?�/�?#?�?�?Y? �?}?O$O�?HO�?lO ~OO�O1O�OUO�O�O �O _�OD_V_�Oz_	_ �_�_?_�_c_�_
o�_ .o�_Ro�__o�oo�o ;o�o�oqo�o*< �o`�o��%�I �m���8��\� n����!���ȏW�� {��"���F�Տj����w����N�PR� }2g�*.VR���_�*���\� �D�.�ېPCL�u�_��FR6:`���0�ůT�T���������%��දK�-�*#.Fޟ|�^�	��j�⩼8�Ϳ\�STM@ؿω����-���Q�\�Hτ��r�/�8A���]�GIF��
����ϳ���Z�]�JPGdߎ��z�7�I���FU�JS���_�����߼�%
Java?Script=�h߃CS.��Ƃ�?� �%Cascad�ing Styl�e Sheets���3�
ARGNA�ME.DT��S��\���$�4�E���}4�DISP*;�Q�0��I�[�����u�
TPEINS�.XML�� �:\���,�Custo�m Toolba�rM|�PASSW�ORD��Q�FR�S:\�O��Pa�ssword Config�,� �P��t�� 9�]�/�(/� L/���//�/5/�/ �/k/ ?�/$?6?�/Z? �/~?�??�?C?�?g? y?O�?2O�?+OhO�? �OO�O�OQO�OuO
_ _�O@_�Od_�O_�_ )_�_M_�_�_�_o�_ <oNo�_roo�o�o7o �o[o�oo�o&�oJ �oC��3�� i��"�4��X�� |�����A�֏e�Ϗ ���0���T�f����� �����O��s���� ��>�͟b��[���'� ��K��򯁯���:� L�ۯp�����#�5�ʿ Y��}��$ϳ�H�׿ l�~�Ϣ�1�����g� �ϋ� ߯���V���z� 	�s߰�?���c���
� ��.��R�d��߈�� ��;�M���q������ <���`������%��� I��������8�� ��n���!��W �{"�F�j |�/�Se� �/�/T/�x// �/�/=/�/a/�/?�/�,?�/P?�/�/�?i6��$FILE_DG�BCK 1^���s0��� < �)
S�UMMARY.DyG�?<<MD:�?�OH0Diag� Summary�O:
CONSLOG�?�?�1HO�OA�Console� log�O;	T�PACCN~O�O%��O_ETP A�ccountin��O:FR6:I�PKDMP.ZI	P<_@8
T_�_E$P�Exceptio�n�_B[�0MEMCHECK�OeO�?o��AMemory� Dataoi6�4n )�QRIP�E{O�_�_�o#c%�[a Packe�t L�Oj4L�$y��R[aSTAT�o�uo�o %~�bStatus�k	FTP_ot�xg�Ammen�t TBD��g �>I)ETHERNE�oy�Q�$��AEthern��`�@figura��_4�qDCSVRAF�{���-sk�� verify �all��j3M4=f�DIFF�����+��c��diff�-���Qk�CHG01"�	����/qC�؟�2�n�2������ 4�?�՟�u�3*��#��� J�߯n��VTRNDIAG.LS䯕���<�z'a�� OpeL���a Anosti�cIg��)VwDEV �DAT=���,�>�0pVis~_�Devicef�s�IMG ��_�����BϩcشImag��q�UP��ES����FRS:\����AUpda�tes List���:0�FLEXEVEN�!�3�L��/q� UIF �Ev�q�oj2-v�Z)
PSRBW�LD.CMx�<<���ϝ@PS_R?OBOWEL�X�:GIG^o+�6�O�>"fGigEh�r�~j2N�@�)@�HADOWJ�/�A����%cShado�w Change�>Ke(dt��RCMERR�����Z��%c�CFG E�rrorްtai}l�� a��cCMSGLIBR��9�K���g��8r��iyc�����)���ZD�:��^!g�ZD{�ad ��= ��NOTIp�=�O�#eNoti�ficM��j5,�AG?;B?_f?l �?�H��~/ �7/I/�m/��/�/ 2/�/V/�/z/�/!?�/ E?�/i?{?
?�?.?�? �?d?�?�?O/O�?SO �?wOO�O�O<O�O`O �O_�O+_�OO_a_�O �__�_�_J_�_n_o �_o9o�_]o�_�o�o "o�oFo�o�o|o�o 5G�ok�o�� �T�x���C� �g�y����,���ӏ b��������(�Q��� u������:�ϟ^�� ���)���M�_�� ���6���ݯl���� %�7�Ư[����� � ��D�ٿ�z�Ϟ�3� ¿@�i�����ϱ��� R���v��߬�A��� e�w�ߛ�*߿�N��� �߄���=�O���s� ���8���\���� ��'���K���X���� ��4�����j�����# 5��Y��}�� B�f��1� Ug����P �t	//�?/�c/��p/�/z#�$FI�LE_FRSPRT  ��� ����(�MDONLY 1�^�%z  
 ��)MD:_V�DAEXTP.Z�ZZ�/Q/(?7;�6%NO Ba�ck file <?z$S�6P./�? ?�?v/�?�?(/O�? +O=O�?aO�?�O�O&O �OJO�O�O�O_�O9_ �OF_o_�O�_"_�_�_ X_�_|_o#o�_Go�_ ko}oo�o0o�oTo�o �o�o�oCU�oy ��>�b�	�~�$VISBCK�(|�!�#*.VD
�|T��pFR:\#��ION\DATA�\?��r�pVision VDU2 ���ȏڏ����"� ��3�X��|������ A�֟e�������0��� T�f�!������=��� �s����,�>�ͯb� 񯆿�'���K��� ��ϥ�:�ɿK�p��� ��#ϸ���Y���}���ϳ�Hߨ*LUI_�CONFIG �_�%6�S� $ 1��#�߰����������
��$$ |x:�<�N�`�r��� *������������ 5�G�Y�k�}������ ����������1C Ugy���� ���-?Qc u������ �/)/;/M/_/q// �/�/�/�/�/�/�/? %?7?I?[?�/l?�?�? �?�?�?p?�?O!O3O EOWO�?{O�O�O�O�O �OlO�O__/_A_S_ �Ow_�_�_�_�_�_h_ �_oo+o=oOo�_so �o�o�o�o�odo�o '9K�oo�� ��N����#� 5��Y�k�}������� J�׏�����1�ȏ U�g�y�������F�ӟ ���	��-�ğQ�c� u�������B�ϯ�� ��)���M�_�q��� ����>�˿ݿ��� ��$�I�[�m�ϑ�(� ����������ߦ�3� E�W�i�{ߍ�$߱��� ��������/�A�S� e�w�� ������� �����+�=�O�a�s� �������������>��  x��$FLUI_D�ATA `����L���>RESULT� 2aLu  �T��+�� �����!3 EWi��~��� ����/!/3/E/�W/i/{/�-?��0����L�/�+� ���/�/??,?>?P? b?t?�?�?�?�?{�/ �?�?
OO.O@OROdO@vO�O�O�O�O��O  �/�G�/_�/+_=_O_ a_s_�_�_�_�_�_�_ �_oo&_9oKo]ooo �o�o�o�o�o�o�o�o �O2�OV_}� �������� 1�C�U�g�&o������ ��ӏ���	��-�?� Q�c�"��F��jl� ����)�;�M�_� q���������x�ݯ� ��%�7�I�[�m�� ������t�ֿ����� Я3�E�W�i�{ύϟ� �����������ʯ/� A�S�e�w߉ߛ߭߿� �������ƿ��4� ^� υ�������� ����'�9�K�]�� ���������������� #5GY�b�<� ��r���� 1CUgy��� n����	//-/?/ Q/c/u/�/�/�/j| ��?�)?;?M?_? q?�?�?�?�?�?�?�? O�%O7OIO[OmOO �O�O�O�O�O�O�O_ �/�/�/T_?{_�_�_ �_�_�_�_�_oo/o AoSoOwo�o�o�o�o �o�o�o+=O a _2_D_�h_�� ���'�9�K�]�o� ������do��ۏ��� �#�5�G�Y�k�}��� ����rԟ����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ���ğ&��J�� qσϕϧϹ������� ��%�7�I�[��� �ߣߵ���������� !�3�E�W��x�:Ϝ� ^�`���������/� A�S�e�w�������l� ������+=O as���h���� � ��'9K]o �������� ��#/5/G/Y/k/}/�/ �/�/�/�/�/�/� �(?R?y?�?�?�? �?�?�?�?	OO-O?O QO/uO�O�O�O�O�O �O�O__)_;_M_? V?0?z_�_f?�_�_�_ oo%o7oIo[omoo �o�obO�o�o�o�o !3EWi{�� ^_p_�_�_��_�/� A�S�e�w��������� я����o�+�=�O� a�s���������͟ߟ �����H�
�o� ��������ɯۯ��� �#�5�G��k�}��� ����ſ׿����� 1�C�U��&�8���\� ��������	��-�?� Q�c�u߇ߙ�X����� ������)�;�M�_� q����f������ ���%�7�I�[�m�� ��������������� !3EWi{�� ��������� > �ew���� ���//+/=/O/ s/�/�/�/�/�/�/ �/??'?9?K?
l? .�?RT?�?�?�?�? O#O5OGOYOkO}O�O �O`/�O�O�O�O__ 1_C_U_g_y_�_�_\? �_�?�_�_�Oo-o?o Qocouo�o�o�o�o�o �o�o�O);M_ q������� �_�_�_�F�om�� ������Ǐُ���� !�3�E�i�{����� ��ß՟�����/� A� �J�$�n���Z��� ѯ�����+�=�O� a�s�����V���Ϳ߿ ���'�9�K�]�o� �ϓ�R�d�v����Ϭ� �#�5�G�Y�k�}ߏ� �߳������ߨ��� 1�C�U�g�y���� �������������<� ��c�u����������� ����);��_ q������� %7I��,� �P������/ !/3/E/W/i/{/�/L �/�/�/�/�/??/? A?S?e?w?�?�?Z�? ~�?�OO+O=OOO aOsO�O�O�O�O�O�O �OO_'_9_K_]_o_ �_�_�_�_�_�_�_�? o�?2o�?Yoko}o�o �o�o�o�o�o�o 1C_gy��� ����	��-�?� �_`�"o��FoH���Ϗ ����)�;�M�_� q�����T��˟ݟ� ��%�7�I�[�m�� ��P���t�֯诬�� !�3�E�W�i�{����� ��ÿտ翦���/� A�S�e�wωϛϭϿ� ���Ϣ��Ư�:��� a�s߅ߗߩ߻����� ����'�9���]�o� ������������� �#�5���>��b��� N߳��������� 1CUgy�J� ����	-? Qcu�F�X�j�|� ���//)/;/M/_/ q/�/�/�/�/�/�/� ??%?7?I?[?m?? �?�?�?�?�?�?�� �0O�WOiO{O�O�O �O�O�O�O�O__/_ �/S_e_w_�_�_�_�_ �_�_�_oo+o=o�? O O�oDO�o�o�o�o �o'9K]o �@_������ �#�5�G�Y�k�}��� No��roԏ�o���� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ᯠ��ď&��M�_� q���������˿ݿ� ��%�7���[�m�� �ϣϵ���������� !�3��T��x�:�<� ������������/� A�S�e�w��Hϭ�� ��������+�=�O� a�s���Dߦ�h����� ��'9K]o ��������� #5GYk}� ����������/ ./��U/g/y/�/�/�/ �/�/�/�/	??-?� Q?c?u?�?�?�?�?�? �?�?OO)O�2// VO�OB/�O�O�O�O�O __%_7_I_[_m__ >?�_�_�_�_�_�_o !o3oEoWoio{o:OLO ^OpO�o�O�o/ ASew���� ��_���+�=�O� a�s���������͏ߏ �o�o�o$��oK�]�o� ��������ɟ۟��� �#��G�Y�k�}��� ����ůׯ����� 1�����v�8����� ��ӿ���	��-�?� Q�c�u�4��ϫϽ��� ������)�;�M�_� q߃�B���f��ߊ��� ��%�7�I�[�m�� ������������� !�3�E�W�i�{����� �������������� ASew���� ���+��O as������ �//'/��H/
l/ .0/�/�/�/�/�/�/ ?#?5?G?Y?k?}?< �?�?�?�?�?�?OO 1OCOUOgOyO8/�O\/ �O�O�?�O	__-_?_ Q_c_u_�_�_�_�_�_ �?�_oo)o;oMo_o qo�o�o�o�o�o�O�O �O�o"�OI[m �������� !��_E�W�i�{����� ��ÏՏ������o & J�t�6������ џ�����+�=�O� a�s�2�������ͯ߯ ���'�9�K�]�o� .�@�R�d�ƿ����� �#�5�G�Y�k�}Ϗ� �ϳ��τ������� 1�C�U�g�yߋߝ߯� ���ߒ������ڿ?� Q�c�u������� ��������;�M�_� q��������������� %�����j,� ������� !3EWi(�z� �����//// A/S/e/w/6�/Z�/ ~�/�/??+?=?O? a?s?�?�?�?�?�?�/ �?OO'O9OKO]OoO �O�O�O�O�O�/�O�/ _�/5_G_Y_k_}_�_ �_�_�_�_�_�_oo �?CoUogoyo�o�o�o �o�o�o�o	�O< �O`"_$���� ����)�;�M�_� q�0o������ˏݏ� ��%�7�I�[�m�, ��P��ğ������ !�3�E�W�i�{����� ��ï�������/� A�S�e�w��������� ~�ȟ����؟=�O� a�sυϗϩϻ����� ����ԯ9�K�]�o� �ߓߥ߷��������� �п���>�h�*Ϗ� ������������� 1�C�U�g�&ߋ����� ��������	-? Qc"�4�F�X�|� ��);M_ q����x��� //%/7/I/[/m// �/�/�/�/���? �3?E?W?i?{?�?�? �?�?�?�?�?O�/O AOSOeOwO�O�O�O�O �O�O�O__�/�/�/ ^_ ?�_�_�_�_�_�_ �_oo'o9oKo]oO no�o�o�o�o�o�o�o #5GYk*_� N_�r_����� 1�C�U�g�y������� ������	��-�?� Q�c�u���������| ޟ���)�;�M�_� q���������˯ݯ� ��ҏ7�I�[�m�� ������ǿٿ���� Ο0��T��ύϟ� ������������/� A�S�e�$��ߛ߭߿� ��������+�=�O� a� ς�DϦ��|��� ����'�9�K�]�o� ��������v������� #5GYk}� ��r����
�� 1CUgy��� ����	/��-/?/ Q/c/u/�/�/�/�/�/ �/�/?��2?\? �?�?�?�?�?�?�? OO%O7OIO[O/O �O�O�O�O�O�O�O_ !_3_E_W_?(?:?L? �_p?�_�_�_oo/o AoSoeowo�o�o�olO �o�o�o+=O as����z_�_ �_ ��_'�9�K�]�o� ��������ɏۏ��� �o#�5�G�Y�k�}��� ����şן����� ��R��y������� ��ӯ���	��-�?� Q��b���������Ͽ ����)�;�M�_� ���B���f������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ��p��������/� A�S�e�w��������� ��������+=O as������ ���$��H
� �������� /#/5/G/Y/}/�/ �/�/�/�/�/�/?? 1?C?U?v?8�?�? p/�?�?�?	OO-O?O QOcOuO�O�O�Oj/�O �O�O__)_;_M___ q_�_�_�_f?�?�?�_ �_�?%o7oIo[omoo �o�o�o�o�o�o�o�O !3EWi{�� ������_o�_ &�P�ow��������� я�����+�=�O� s���������͟ߟ ���'�9�K�
�� .�@���d�ɯۯ��� �#�5�G�Y�k�}��� ��`�ſ׿����� 1�C�U�g�yϋϝϯ� n������϶��-�?� Q�c�u߇ߙ߽߫��� ���߲��)�;�M�_� q����������� �������F��m�� �������������� !3E�V{�� �����/ AS�t6��Z�� ���//+/=/O/ a/s/�/�/�/��/�/ �/??'?9?K?]?o? �?�?�?d�?��?� O#O5OGOYOkO}O�O �O�O�O�O�O�O�/_ 1_C_U_g_y_�_�_�_ �_�_�_�_�?o�?<o �? ouo�o�o�o�o�o �o�o);M_ q������� ��%�7�I�oj�,o ����dǏُ���� !�3�E�W�i�{����� ^ß՟�����/� A�S�e�w�����Z��� ~�ȯ򯴏�+�=�O� a�s���������Ϳ߿ 񿰟�'�9�K�]�o� �ϓϥϷ������Ϭ� ��Я�D��k�}ߏ� �߳����������� 1�C��g�y���� ��������	��-�?� ���"�4ߖ�X߽��� ����);M_ q��T���� %7I[m ��b�t������/ !/3/E/W/i/{/�/�/ �/�/�/�/�??/? A?S?e?w?�?�?�?�? �?�?�?���:O� aOsO�O�O�O�O�O�O �O__'_9_�/J_o_ �_�_�_�_�_�_�_�_ o#o5oGoOho*O�o NO�o�o�o�o�o 1CUgy���o ����	��-�?� Q�c�u�����Xo��|o ޏ�o��)�;�M�_� q���������˟ݟ� ��%�7�I�[�m�� ������ǯٯ믪�� Ώ0����i�{����� ��ÿտ�����/� A� �e�wωϛϭϿ� ��������+�=��� ^� ��ߔ�Xϻ����� ����'�9�K�]�o� ���RϷ��������� �#�5�G�Y�k�}��� Nߘ�r߼����� 1CUgy��� �����	-? Qcu����� �������/8/��_/ q/�/�/�/�/�/�/�/ ??%?7?�[?m?? �?�?�?�?�?�?�?O !O3O�//(/�OL/ �O�O�O�O�O__/_ A_S_e_w_�_H?�_�_ �_�_�_oo+o=oOo aoso�o�oVOhOzO�o �O'9K]o �������_� �#�5�G�Y�k�}��� ����ŏ׏鏨o�o�o .��oU�g�y������� ��ӟ���	��-�� >�c�u���������ϯ ����)�;���\� ���B�����˿ݿ� ��%�7�I�[�m�� �Ϣ������������ !�3�E�W�i�{ߍ�L� ��p��ߔ�����/� A�S�e�w����� �������+�=�O� a�s������������� �� ��$����]o �������� #5��Yk}� ������// 1/��R/v/�/L�/ �/�/�/�/	??-??? Q?c?u?�?F�?�?�? �?�?OO)O;OMO_O qO�OB/�/f/�O�O�/ __%_7_I_[_m__ �_�_�_�_�_�?�_o !o3oEoWoio{o�o�o �o�o�o�O�O�O, �OSew���� �����+��_O� a�s���������͏ߏ ���'��o�o
 ~�@����ɟ۟��� �#�5�G�Y�k�}�<� ����ůׯ����� 1�C�U�g�y���J�\� n�п����	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹����ߜ� ����"��I�[�m�� ������������� !���2�W�i�{����� ����������/ ��P�t6��� ���+=O as������ �//'/9/K/]/o/ �/@�/d�/��/�/ ?#?5?G?Y?k?}?�? �?�?�?�?��?OO 1OCOUOgOyO�O�O�O �O�O�/�O�/_�/�O Q_c_u_�_�_�_�_�_ �_�_oo)o�?Mo_o qo�o�o�o�o�o�o�o %�OF_j| @o������� !�3�E�W�i�{�:o�� ��ÏՏ�����/� A�S�e�w�6�Z�� Ο�����+�=�O� a�s���������ͯ�� ���'�9�K�]�o� ��������ɿ��ҟ�� �� ��G�Y�k�}Ϗ� �ϳ����������� ޯC�U�g�yߋߝ߯� ��������	��ڿ� ���r�4ϙ����� ������)�;�M�_� q�0ߕ����������� %7I[m >�P�b������ !3EWi{�� ������//// A/S/e/w/�/�/�/�/ �/���?�=?O? a?s?�?�?�?�?�?�? �?OO�&OKO]OoO �O�O�O�O�O�O�O�O _#_�/D_?h_*?�_ �_�_�_�_�_�_oo 1oCoUogoyo�_�o�o �o�o�o�o	-? Qcu4_�X_�|_ ����)�;�M�_� q���������ˏ�o� ��%�7�I�[�m�� ������ǟ�蟪� �ПE�W�i�{����� ��ïկ�����܏ A�S�e�w��������� ѿ�����؟:��� ^�p�4��ϩϻ����� ����'�9�K�]�o� .��ߥ߷��������� �#�5�G�Y�k�*�t� NϘ���������� 1�C�U�g�y������� ��������	-? Qcu����|� ������;M_ q������� //��7/I/[/m// �/�/�/�/�/�/�/? ���f?(�?�? �?�?�?�?�?OO/O AOSOeO$/�O�O�O�O �O�O�O__+_=_O_ a_s_2?D?V?�_z?�_ �_oo'o9oKo]ooo �o�o�o�ovO�o�o�o #5GYk}� ����_�_�_
��_ 1�C�U�g�y������� ��ӏ���	��o�?� Q�c�u���������ϟ �����8��\��j��$FMR2_�GRP 1bj��� ��C4  B�#�	� #�������E��� E�  F@ F�5Uܥ����L���M���Jk�K��v�H�,�Hk{��?�   �����9tQvH�8���6h�%T���A�  p���BMH��B��������	@�����ʿ۽��/@UUU�U�۽�>�]�>П���;r8	=�==E��<D��><�ɳ<�����:�b�:/�'79�W�9
�@�8�8�9�ϑ�ܿ���Ϣ��E7� E?p �D������D�  D�  C����#�~�_CFG =c��T �[��m��!�NO ^��
F0�� ��� �RM_CHKTYP  {�#������K�}�ROM��_�MIN��#��������X~�SSB�1�dj� ��/�#�&�O�a��'�TP_DEF__OW  #���>v�IRCOM�Ї���$GENOVR/D_DO��-���THR�� d��d޺�_ENB�� ^��RAVC��e��#� �ȥFn�H E�� Ga� H�� H�?@Jh`��K��|�������� ���OU��k�������⸥< ��2���&T#�+C�������j)� �#�����������h��SMT��l�(���%�y�$HO7STC1�1m��$��-� 	O&OO#� �e����/* �3/E/W/i/��/  �	anonymous�/�/�/�/�/? N`rO?�/�"/ �?�?�?�?/�?OO 'O9O\?�/�/�O�O�O �O�O?"?4?F?HO5_ |?Y_k_}_�_�_�?�_ �_�_�_o0_fOxOUo goyo�o�o�O�O_�o o	P_-?Qc�_ t�����o�:o �)�;�M�_��o�o�o �o������%� 7�~[�m������Ə ������!�3�z� ����L������ïկ ������/�A�S�e� ����П����ѿ��� <�N�`�r�Oφ����� �ϩϻ�������� '�9�\ϒ����ߓߥ� �����"�4�F�H�5� |�Y�k�}������� ��������f�C�U��g�y����1ENT� 1n�� P!\���  � �� ��,��Pt7 �[����� �:�^!3�W �{�� /��6/ �Z//~/A/�/e/�/ �/�/�/�/ ?�/D?? P?+?y?�?a?�?�?�? �?
O�?.O�?OdO'O��OKO�OoJQUICC0�O�O�O_�DA1	_�O�OX_�D2Y_�5_G_�_!ROU�TER�_�_�_�_!?PCJOG�_�_�!192.168.0.10�O~�CCAMPRTIo%o!9e1B`poWf�RT�_to�o�o !�Softwar�e Operat�or Panel��o6o7��NAME� !��!RO�BObo?S_CF�G 1m�� ��Auto�-started^��FTP���q ���H��1�C�U� g���������ҏ�x�	��-�?�Q��#��֩������ �����(��L�^� p�������9�ʯܯ�  ��$������� ��ן��ƿؿ���ï  �2�D�V�hϋ�Ϟ� ����������?�Q�c� @�w�d߫��ߚ߬߾� ��������*�M��� I�r������� %�7�9�&�m�J�\�n� ����Y���������� !���4FXj|� ��������A� 0BT��� ���w//,/>/ P/������/ �/�/??(?�L?^? p?�?�?�/9?�?�?�?  OO$Ok/}/�/=O�? �O�/�O�O�O�O�O�?  _2_D_V_yOz__�_��_�_�_�_zNp_ERR oXz�_f�PDUSIZ  ��P^�@�d>~6eWRD ?�u�hA�  guest�Vvo�o��o�o�o�oGtSCD�MNGRP 2p�u `��hA�P���VKt 	�P01.05 �8MA   
��  3  ͬMpLpٝ�CK ����U��������3uptp�'����]}$o�h���wDp���U�Mp�Z@Z@U]������t�p�up���Hp�}��5�li@6i@I=��zdASew�k__GROU pqi�p�b	�a8q4���QUPD  ddEe���TY���m`TTP_AUTH 1rk� <!iPeOndan�gR��_���!KAREL�:*R�[�m�KC ������z�ݟ˟���q �@��)�v�M�_������������˯ݤ!�C?TRL smq�>��Q
�QFF�F9Eh�\�hBF�RS:DEFAU�LT`�FAN�UC Web Server`�N�>� !�^opd	�ֿ������0�dWR_CONFIG t{� `�aIDL_CPU_PC���QB�i@�� BH��MIN��Na��?GNR_IOaDb��Ph��NPT_S_IM_DO�����STAL_SCR�N�� ���INT�PMODNTOL8��˻�RTY�Ȣ����VIS%�ENB������OLNK 1ukr`�߼�����������MA�STE���SL?AVE voE��RAMCACHE�4�,�O'�O_CF1Gv�ӎ�UO���~��CMT_OP�8��j��YCLu���y�_ASG 1wwPa
 �;�M� _�q����������������% ��NU�MCci
��IP�s��RTRY_C�N�����Cc���be �����xT��j`�j`��P�?�T� ��	�*< N`r���� ���/�,/>/P/ b/t/�//�/�/�/�/ �/?�/�/:?L?^?p? �?�?#?�?�?�?�? O O�?6OHOZOlO~O�O O1O�O�O�O�O_ _ �OD_V_h_z_�_�_-_ �_�_�_�_
oo�_�_ Rodovo�o�o�o;o�o �o�o*�oN` r���7I�� ��&�8��\�n��� ������E�ڏ���� "�4�ÏՏj�|����� ��ğS������0� B�џf�x��������� O�a�����,�>�P� ߯t���������ο]� ���(�:�L�ۿ� �ϔϦϸ�����k� � �$�6�H�Z���~ߐ� �ߴ�����g�y�� � 2�D�V�h��ߌ��� ������u�
��.�@� R�d������������ ������*<N`�r�_MEMB�ERS 2y��   $:��������	� RCA_A�CC 2z��   [��� Sȴw6O�"    '!+�C�BUF00�1 2{= ��u0  u0��(�N�s��j������U2�X�}��������$8�$`$�$�$��IP  IP��V���9$�9$���� Q$FQ$kQ$�jQ$�Q$ݙ��$������ %[� � �%�$J�$Up�$��$��$���	�$.�$S�$y��$��$��$ $��474]4�4�j4�4���I4UEI4jI4�I4�I4	ۙv2���� �2��2��2��2� �2����2��2� �2��2��2��2   �!B B B   B( B0 1!7!�?! DBH DBP �W!\B`  \Bh \Bp \Bx \B�  ��!�B�4�!�B�4�! �!�!�B� �B� �B�  �B� �B� ��!�B�  �B� �B� �B 0�B0 �B	D1R 0R(0R 00R80R@0RH0� O1TRX0TR`0TRh0TR p0TRx0�v3�?� �3�R��3�R��3�R ��3�R��3�R��3 �R�C#Cb" &Cb("6C7#FCEb H"VCW#fCebh"vC ebx"�C�#�C�b�T �#�C�b�"�C�b�"�C �b�"�C�#�C�b�" �C�b 2S�bd3&S %r(26S%r82FS%rH2 VS]rX2fS]rh2vS]r�x2�VCFG 2| 4 � �z� < �t�q��xHIS�~� � 202�5-12-� ~1�C�U�g�y�苏�����7  �A;�Aʃ˂��� ��	��-�?� Q�c�u��������� ����)�;�M�_� q�����̟��˯ݯ� ��%�7�I�[����� ������ǿٿ���� !�3�j�|���{ύϟ� ������������T� f�S�e�w߉ߛ߭߿� �������y�0��� L�^�p�������J��6 dI݁dЀ ����,�>�(�:�L� ^�p�����������(� � $6HZl ~���������  2DVhz� ������
// ./@/R/d/���/�/ �/�/�/�/??*?<? s/�/r?�?�?�?�?�? �?�?OO�P�)� ;�qO�O�O�O�O�O�O �O��K0Ȃ�bK3؂N? `?J_\_n_�_�_�_�_ �_�_�_J?5_"o4oFo Xojo|o�o�o�o�o�_ oo0BTf x����o�o�� ��,�>�P�b�t��� ����Ώ����� (�:�L�^��������� ��ʟܟ� ��$�6��$MI_CFG 2�=K H
C�ycle Tim}ev�Busyp��Idl}�t�m�in@���U�py�w�Read>��Dow����� ��t�Cou�ntw�	Num Dt�u��l�#�p�����PROGZ��=EG@�3�x����������ҿ��E�SD�T_ISOLC ; =I� ���J23_DSP_?ENB  ˳�~.�INC �>��p��A   ?��  =���<#��
�u�:�o ���ϫ�p�����'�+OBN�C7���`����G_GROUPw 1��<��<��s�n�9���E?o�g�x�p�Q�� �����ߖ�����1��p�����G_IN�_AUTO��B�P�OSRE���KA�NJI_MASK���^ȫ�RELMO�N �=K+�p�y ���!�3�E�W����JR��Y�I�p�y�|��J�KCL_Lo��NUM;���$KE�YLOGGINGī�B@�-�F�I�LA�NGUAGE �=E �DEFAULT #6+ALG[��Y�����p�xl�P8n��H  #Q'0o��� 
�p��p��޿�;��
�(?UT1:\g�� ����� 0GTfx�p��(�����  N_D?ISP �Xϯ���ߋ�)CLOCTOL$ p�DzC��q��:!GBOOK �4d�����r X��/�/�/�/�/��+ =@��9�&	@X%�	5��^?{V"�_BUFF 2�N� z�p�2�� �?q"�?���?�?O O!ONOEOWO�O{O�O �O�O�O�O�O___�J_�P�DCS �Y�d�y�<N?o�a��_�_�_�_aTIO ;2�m[ ��o5��!o1oCoUoio yo�o�o�o�o�o�o�o 	-AQcu�������UER_ITM
�dO�*�<� N�`�r���������̏ ޏ����&�8�J�\��n�����4'�rSEVt��>��vTYP
΁���������R�ST��_USCRN�_FL 2�
mC���_������ȯگ���/�TP��
��}.-NGNAM7���%�UPS_A�CRG���m�DIG�Iw�F�m�_L�OAD��G %�+�%REQME�NU�-,MAXU�ALRM��z�.0e�F�
񲒱_Pv��z� L#1�C���4�/�?�83��Pw 2�b+ ر6�	:���]  �Z�D���ϻ��� ߐX��5� �Y�<�N� ��z߳ߞ�������� ��1��&�g�R��v� ���������	����� ?�*�c�N�����|��� ��������;& _qT����� ���7I,m X�t����� /!//E/0/i/L/^/ �/�/�/�/�/�/�/?�?A?�DBGDEF �<�I�H�J?�\0_LDXDIS�AX�*��SMEMO�_APR�E ?+�
 n1UX�? �?�? OO$O6OHO��FRQ_CFG k�<�r3A VW�@��CVP<I�d%�KL�O\On@�<�{��* P=/R **:RVT �OX�O�6_H_u_l_ ~_�_�_�_�_-?<�
o��p�_1ol*o@j,( �_�o�vo�o�o�o�o �o�o1UgN��r�����I�SC 1�+��@ �3?-���s?C�.?|��g�����_MST�R ���ÅSC/D 1��=���� ��6�!�Z�E�~�i�{� ����؟ß��� �� 0�V�A�z�e�����¯ ���ѯ���@�+� d�O���s�������� Ϳ��*��N�9�K� ��oϨϓ��Ϸ�����  �&��J�5�n�Yߒ� }߶ߡ߳�������� 4��X�C�h��y�������������M�KqA�ҍ�A0�$�MLTARMpBu��G[� $c�l0����[0METP�U�0����ډN�DSP_ADCO�L��p0��CMNT6�� ��FN����>��FSTLIˀ �Ҏq��A�����POSCFz?PRPM����	ST��1�ҋ; 4�B#�
"a +	+-?� cu������ #///Y/;/M/�/y!���SING_CH�K  !$MODAoC��Y�[�~�%DEV 	�:�	MC:�,HS�IZE�=����%T�ASK %�:%�$1234567�89 j?|5�'TR�IG 1�ҋ l[5�O�?Vi�?�?VmFL6YP71Ve�$�#�EM_INF 1���K`)AT&FV0E0�?�uM)]AE0V1�&A3&B1&D�2&S0&C1S�0=dM)ATZuO�O�DH�O�O�A�?_�HA%_M__q_X_�_�_ [O�_O�O�O �O&o�OJo�_no�o3_ �o_o�o�o�o�o�_�_ 4�_�_o|�oAo� �o���o��0�� T�f���=Oas 䏗�?��>��b� ��������o���� ����ɏ:�L���p��� ��O�Y�ʯ���կ� $�ןH�����1��� U�ƿؿ����� �ۿ�1�V�=�z��/NIT�ORZ G ?; �  	EXESC1��2��3��E4��5�ȍ0��7��8��9���D�(� ��(���(���(���(� ��(���(�
�(��(�T"�(�2/�2;�2G�U2S�2_�2k�2w�U2��2��2��3/��3;�3���!R_G�RP_SV 1�JK (�m��%T1�_D�:>��ION�_DB� ��-A/  �@G�(��������'p�N� �,���)-u�d1#59�K�]���P�L_NAME �![5���!D�efault P�ersonali�ty (from� FD)���RM�K_ENONLY�/��R2A� 1��L�XL�<����l d^� %7I[m� ������! 3EWiH2��� �����//)/;/���e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogoyo|<T/�o�o�o�o�o�o 1CUgy��D�o�}
��|P� ���'�9�K�]�o� ��������ɏۏ��� ��5�G�Y�k�}��� ����şן����� 1�C��$�y������� ��ӯ���	��-�?��Q�c�u����� �FnH F�� gG=�|]��ƿؽ|d\����� +�9ǫ���z]�|�g��ϣ� �ȿϵ� ���������=ߓ���h`�p�|��	`���ߵ��߆�:�o�A��� ��| �A�  2��,��� ||���0������  �h  3�=���S���Ϫ�����������(�S�d�R�R��~������ | ����|� @D�  ��?����{�?|��|A��Ǐ�K%H�  �;�	l��	 �X8  ���������� � _� � l����K(��K(��K ��J�n��J�^J&u������Wa��@Y�,@Cz?@I�@Ɂ���:I�=�N���f��N���_�� a������?�*  �� W �9� H� � ���|?s8y��
�/|�x�	�� �M�!|���:���D
�  �Y��w�s�7  ~Ї���H	'� �� �I� ��  �?�F:��È�È=��������]����� F��9/�ہ��)�/HN�Б/  '��&t� @2��_@���@� @� �@�C� C��C���\C� C� Cz����@@1	�	�	� -_ EB3��?6��K5"�1g5��Dz��?��?�?�?�?��2�l� ���E1E  R�Һ55��p7A?�ffJ�EOWO�?C �ЌO�K�18��<�O�J?��7��C
(���EP�HI������Y#?L	 8D�1�;�Cd;�pf�<߈<��.<p��<�?�J�3��@��ۗ������/�?fff?�0?&�PH@��׳R�N�@T���U��2�Q��C	�� �_��o�V��vOKo6o ooZo�o~o�o�o�o�o0�o���UF��  M�oq�_�id��`xC��E����Gd G;�\��  �9�$�]�H���l�~� ����ۏƉn/�̏-� �N��u�菙�����dϟ�����dOA�� !����W�B�{�F��!A|P��;���Ck�Яg�U����$���|H�3�  �P������.40DE� C x5��B������� �S�B�/B�"�}A��#A���9@�dZ?�vȴS��~���<)�+� �=�G��������q���
AC
�=C��������� ��p��Cc�¥��B=���ff��{S�I����HD-�H�d�@I�^�F8$� D;q�oʭ̠�Jj��I�G�FP<���x�QpJnPH��?�I�q�F.� D�|\8�� ��%��I�4�m�X�j� �ߎ��߲�������� 3�E�0�i�T��x�� �����������/�� S�>�w�b��������� ������=(: s^������  9$]H� l������� #//G/2/k/}/h/�/ �/�/�/�/�/?�/
?�C?.?g?"�('���33:n?'Q���5W5�3�V��?�?�2���?�?�4M���?�?��=��O%O4Ue'��T9?M?IOmO�O�O(�O�L�P_RP�N���"_u?._X_C_|_gY���(�_�_�_`�_�_�_�_�B��_ oFo1ojoUo�o5_�0�o�o�o�k/�o�o�+;aO��{f gy�������  2 FnHn�F���G=�1B�0����C9��"`��@��m�����E��� F�5��H C፰��ɏ���M�E�h�1�a�o�0�B��?q�c��@*��d���9i���
 Q��� Ɵ؟���� �2�D��V�h�z������l�����;�~Y��$�MR_CABLE� 2��H �x�QTP@@�Y�`��������u��`�C��O8�tBx�@����+�`�M��O��1��H�>Q��c�
P�
PCQ�6'�~ȅ��������2�1�C�)�HE�ٿ�7��T�K o�G�YϾ�}��Ϲϳ� ������N�I��k�C�@Uߺ�y���1��A�� �"�4�yh��c�u���yh*��** �ףOM ������%ybST=�%% 23456�78901���� �����y`�y`\��y`ya
����not sent� ��9�W�E�TESTFECS�ALGR  egDwj\�d��@�
��P�Pydl�yg�������
 9U�D1:\main�tenances�.xmlY  ����DEF�AULT܌עGR�P 2���  �E�ye  �%�1st mech�anical c�heck�ya�B�d����@ �1CUgyyb��controll�er������"�	//-/?/�1M�g/yb"8}#ʰ�"�/���/�/�/�/�/J*C�-?|/Q?��/?�?�?�?�?ڎC� ge�. battery�?A?O�	n?COUOgOpyO�O�9�dui�Oable�O��p�C��O'G2O__�+_=_O_��4grgeas�Oygf��S!-y`�Q�_��O�_��_�_oo�
�4oaiG�_�_�_�_@�o�o�o�o�o��:,�O����s<��q&�
~oSew����Lt�?�B�)�;�M�_��Overhau`/6�|��� x��������ۏ����#���$̏K�����z� ʏ����ß՟�6� �Z�l�~�4�e�w��� ������ѯ �2�D�� +�=�O�a������� ��
�߿���'�v� K�]Ϭ���п�Ϸ��� ����<��`�r�Gߖ� k�}ߏߡ߳����&� 8��\�1�C�U�g�y� �ߝ�������"���	� �-�?���c������ ���������T�) x���_������ ��>PbI [m��� (�/!/3/E/�� {/�j/��/�/�/�/ ?Z//?A?�/e?�/�? �?�?�?�? ?�?D?V? +Oz?OOaOsO�O�O�? �O
OO�O@O_'_9_ K_]_�O�_�O�O�__ �_�_�_o#or_Go�_ �_}o�_�o�o�o�o�o 8o\onoC�ogy ����o�"4F �-�?�Q�c�u���� �������)�8;���҂	 X=�j�|���҉B ����ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ�����!�3�E�WϽ� о݁?�  @ҁ ���ϨϺ�҆��p�����҈*+�** F�@ �� ����]�c�u߇�I߫�8������������ E���5�G�Y��}�� ������q����� e���U�g�y������� ����������-? Q�����������]>���ҁ�$MR_HI_ST 2���q�� 
 \��$ �23456789C01��?%��9~�����|�:/ L/^//'/�/�/�/o/ �/�/ ??�/6?�/Z? l?#?�?G?�?�?}?�? �?O O�?DO�?hOzO 1O�OUO�O�O�O�O҄�]SKCFMAPw  ��t)��XҀ _U�ONREL  �҄q)QVREXC/FENB[W
'SU�tQFNC{_mTJO�GOVLIM[Wd�q�PRKEY[Wz�U�U_PANZX��R�RRRUN�\��[SFSPDTY�P�XfUSSIGN|[_mTT1MOT�_�jQR_CE_G�RP 1��� )SyU����o҃�o�o \d�o�o>Pt +��a���� �(�:�!�^������ {���o��Տ�ɏ��H���l�#�QQZ_EDITXd#WLc�TCOM_CFG 1�]~U˟ݟ�� 
��_ARC�_xR[e�YT_M�N_MODEXf=磚_SPL��VUAP_CPLT���TNOCHECK� ?[ �O ����ͯ߯�� �'�9�K�]�o����������D[NO_WA�IT_LWg���`N�T���[.�DS�	�_ERR�a2�YV���`�rτ��̠7Q�ϻ��.�O7ó>>�| S��a��2DQ<`S?�B[&���:P��0�PARAuM8´[�6R�X�ϩ�^�X���� = �������1� C��O�y��g������]�������)�~LbODRDSPS��Zf�XOFFSET�_CAR��z�_�DsISl�]�S_A.��ARKXg��OPE?N_FILE��Za�򑢖
�OPTIO�N_IO�_�Q��M_PRG %Z�%$*.��WO�����g���S_J6R��y �y	 �DXyJ�DS�?�RG_D?SBL  i)Q�"��<�RIEN�TTOZPDQC��9P(QA =�UN�IM_D��&R��?��VC�LCT �@͞�r�dDUdj	;_PEX6�����RAT6� d�U|�d�UP �H
��R ����!/�/)�$s�2�c�L�XL�2l{�w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�?�?�?DW2e/O O2O DOVOhOzO�O�O�O^b�?�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p����� ����ʏ܏���O� (�:�L�^�p������� ��ʟܟ�:��� �<�:�P)�f�x� ��������ү���� �,�>�P�b�t�C�U� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����������������;�M�w�k�}�b� ��� � ���������z 
�4�*�<�N� l�r������R ������	�	`�*<<��:�oZ�l~���A� � �	�,������������0��}��  h�~� =�  GS�A �����CU@y�d�����C$K OU�N �)��)��HZ$� |� ��� �@D�  !?��#�?��"��D	�"!�E�  ;��	l"	 X8  �b!�Y  � �/ � lx"�~"��H<zH<W��H3k7G�C�G���G9|���>/5��/�$�C_C  C/� 4� ��#(!?�#�*  ��  �9&0H&0&0�? ?2?��BY����}���^�H�� `?� �?��!�3�|�*�  � ���0��0�  �0� F�O�%	'� � <B�I� �  ����&=���`OrKC!��   �(��O���D�I�O�&NX 
_  '� V�!I0CX C�W�\CU0CY0C]?�/_A_����@@~�)	�	� �-� �'B � �VX �U��Q�U$"z�ob?'oo7o]o�HbIAl� ��LB�e}Q�e  �����R�A�!��p�a?�ff��o�o�bo ��{Ia8x��-;z?���1$!�*(��iuPrx�i0o!h#h$�C?L�@�d�Ha;�Cd;�p�f<߈<���.<p��<�?�Xz�/�g@���!���"� ?fff�?�P?&��$@���,��N�@T�8����R�=I` %p�(���vT$�oď ���ӏ���0��T� f�Q�����s������@[�}��ݟ>�٘C	 �E��D"Gd G;��-���y����� ֯�������0��T� ?��O��E����ǿ%���a��$�6�H��j�	�oAϚ����� �ϻ��Ͽ&WA�p��	B+C��I����?X�?��w�~߷ߢ�D)�P�D"L1H^�PDE� C�Uﻳ�Կ�А�4�@I��8=B�/B"��}A��#A���9@�dZ?v�ȅ;���~���<)�+� =��G��v䀽q����
AC
=�C��������� ��p�C�c�¥�B�=���ff��{8=I����HD-�H�d@�I�^�F8$ �D;����̠J�j��I�G?�FP<����QpJnPH��?�I�q�F.� D��|��z�e� �������������� @+dO�s� �����* N9K�o��� ���/&//J/5/ n/Y/�/}/�/�/�/�/ �/?�/4??X?C?|? �?y?�?�?�?�?�?�? O	OOTO?OxOcO�O �O�O�O�O�O�O__ >_)_b_M_�_q_�_�_�_�_��(���3�:�_�q��e�U3��V�oo(b��4oFo��4M��x`oro��=ӌo��o4Ue'��T9�m�i�o�o
@�.|i�P�rPr~�� ����_�����y���(��;�&�0K�q�\���B�t��� �����Ώ����:�(�^�L�/d�n���`����ڟȟn�{f����(��L�:�p�~�  2 FnH��F�Е�G=��B/`��C95Л����@!����
���E��� F����H �C���B���o����{�������ÿ��?P��ܱpp���������k��o�
 ʿ-�?�Q�c�uχ� �ϫϽ��������������\k�~Y���$PARAM�_MENU ?��e� � DEFP�ULSE��	W�AITTMOUT�{�RCV�� �SHELL_W�RK.$CUR_oSTYLy����OPTС��PTB�����C��R_DECSN��cu�0�B� T�}�x��������������,�U�P�S�SREL_ID � �e�q�d�US�E_PROG �%_�%Q���e�CC�R��v�qg���_H�OST !_�!����T�p��'��� )c��_TGIME��v���P�?GDEBUGt�_��e�GINP_FLgMSK��	TR���PGA�  ��j��CH��TY+PE\�h�P�J� �������� /9/4/F/X/�/|/�/ �/�/�/�/�/??? 0?Y?T?f?x?�?�?�?��?�?�?�?O1O�W�ORD ?	_�
? 	PR� ��MAI-�	�SU��lCTEJ �-Hs	��yBCOL�h�I�O.L�� �`՜����d�TR�ACECTL 1�ei� �pp�p"_!S�FD/T Q��eMPP�D � bsZ_l_~_�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�o�o�o�o �o
.@Rdv �������� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ����"�4�F� X�j�|�������į֯ �����0�B�T�f� x���V_����ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� ^�p������������� �� $6HZl ~�������  2DVhz� �������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o �o�o�o�o�o, >Pbt���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п�����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶�����������"�4�F�P��$�PGTRACEL�EN  Q�  ��Q���f�_UP �/����������  ��f�_CFG7 ����P������������|x���  ������DEFSPD ����O�x���f�H_CONFI�G ���}� UQ�Q�d\��u� O�_�P����{�Q��f�IN��T�RL �����8l���PEA��K������[���f�WLID�����	���LLB 1�K�� �|�Bk�B94;�� |�T�N��� <<=��  ?�~� ~����� 3Q7Ik����g/�/9/��2/o/b/t/�/��G�RP 1� �zQ�A��333P��A��D�@ �D�� D@ A@O-T`���9"9[�[�� �/v�>>´u3W?@;B x0�1?i?{?�?�?�?��
��?�����?0OBN,O =o=	7LGO�OCO }O�O�O�O�O_O�O"_��O2_X_C_  Dz}S�_Q�
m_�_]_�_ �_�_o�_,ooPo;o to_oqo�o�o�o�o�o� z!P�
V7.10beta1�� A��/q�B1��@�!,p>�y�#Cq;3���+q@�
=Sq>a�G�+rm8cq>��z�!�!�!;q;t�  ������Ap���2k��	��-� ���o�5�oI��>l�V�@��z�ۏ��,p\��"��u0�����N���F���Pq�!�p�r� �B�B�m�_�BHT���Q�Q��&|�����ǒ�x˔x7��3����t�S����`=��_�;�k�\�o�u�_�A𘯺����KNOW_M  ������SV �K� r���_/�A�S���w�@b�t���P�=��M�#]�K� �;r	��?	�	� �������� ���"Pqx{b�g�c�,����MR�#��1�Ώ�X�5���˱-OADBANFWD����ST�!1 1����4��;�;r Q���9�K�]ߎ߁ߓ� �������� ����V� 5�G��k�}����� ���������2%��8���<b�6�!�A3L�^�p����4���������5��(�6EWi{�A7�����8���!�MA��4I��OVLD  Aϭ/��PARNUM  �(����SCH� �
''�5)�G%UPD��R5|�/��_CMP_ذ��)��'թ$E�R_CHK�%�������&�/�+RS8���ס_MO�(8�_?��_RES_G$��A
���? �?�?�?�?�?OOO FO9OjO]O�O�O�Of7K�s<�?�Oh5���O �O�Oj3��_0_5_j3 D P_o_t_j3� �_�_ �_j3� �_�_�_j3=�o,o1oj2V 1��+���@k�p�+2THR_INRФ�����d�fMA�SS�o Z�gMN��o�cMON_QU?EUE �(��T��q��N� U�!qN�fx/sEND4qR?NyEXE]Nus �BE\p>/sOPT�IO;w[;2pPROGRAM %z�%1pko/0rTA�SK_I��~OCFG �/�^9�DATA۳�B�"�2������̏ ޏ�����&�8�J�\�����������i�IN+FO۳ц��!tr� �!�3�E�W�i�{��� ����ïկ������/�A�S�e�w�җޔ�Ɔ� �I8�. K_�<��B�����EN!B�Ƚ@��2���G<�2�Ȼ X�,		�!=��=�Oϸ�@��hā$3��!g�gɏd��_EDIT �B������5�WERFL�~x�c�RGADJ� ֬�A�  �?X &սa��2qñ����?��  Bz�X <g�X ��%S���ȡM�:Ֆ�2�H��	H�)pl�&�bBP���UT@V����*
�/� **A:���7�$��]`A��8���zߠo����iX"R���`�������(��A]`������� ~�(�z�d�^�p����� ��������V R< 6H�l���� .�* �D ��z�/�/� ��r//n/X/R/d/ �/�/�/�/�/�/J?�/ F?0?*?<?�?`?�?�? �?�?"O�?OOOO �O8O�OtOnO�O�O�O �O�O�O�Of__b_L_ F_X_�_|_�_�_�_�_��	U�_o��Mo�oqd�t$ �o�kto�o�po�o8�PREF� �H�����
~��IORITY�w��ƀ�MPDSP0�q��p�fwUT$��Ӿ��ODUCT!�e����OG���_TG��&��ʥrHIBIT_DO����{TOENT 1�۬� (!AF_INE�pC�N�?!tcpN�v��!ude���!icm��;�rkXYA�ܬ�����)� "��������=� �,�i�P��� t���ß���Ο�� �A�(�e�w�*�sAӁ�H�p�yߺ�̯��>W��J �"�/,�H�������ܬ�Aj�?,  �>p��@g�y�������C���Z�ݿ��������ENHANCE� ߘ���A��dx�s�Z�  ʡv�'t�/As���PORT_NUM�s���]u�_C_ARTRE���>ׂSKSTA�w�oSLGS@�����j�xpUnothing{�\�n� �ߐ�B߳�������TEMP �y���e��_a_seiban�oK��o [��l�������� ������G�2�k�V� ��z����������� ��1U@ydv ������ +Q<u`��� ����//;/&/ _/J/�/n/�/�/�/�/ �/?�/%??I?��џVERSIop�w��0 disa�ble��`=SAV�E �z	2670H844Z8	F?�?!c��?�?���O 	<H�ronKeOtse�O�O�O�O�O��J�LO"_���7_��p 1���0�iP9b�Us_�_�W pURGE2�B�p	�؁�WF�P��tH��vW�<��T{q��WRUP�_DELAY ����wvb_HOT %�u�rb�Vo�U�R_NORMAL�5h�rEo�oigSEM�Iyo�o�oqQSKKIPQS��bSxD? #@?GYk.}�u� �w������� �>�P�b�(���t��� ��Ώ��ޏ��(�:� L��p�^�������ʟ ���ܟ�$�6���F��l�Z��������5�$RBTIF�TjҠ�CVTMOU�v���ҠDCRQS}�y �:u�CL�CL	��A7�fy8s�F���@���~%��a5.~�A� �;�Cd;�pf�<߈<��.�>�]�>П������z����  ���,�>�P�b�tφ���Ϫϼ������eRD�IO_TYPE � X]Կ��EDP�ROT_CFG ��w#�9TBHf�SE6��a2�H�7 �ѱB�[Џ� ��ѿ��u�������� ��<��oc���v��� ����������&�4� R�W�ܥ���n����� ����������"D�I h�jz���� ��.3Rf  �x����� /*//N/�P/�/ t/�/�/�/�/�//? +?�/L?�/p?^?�?�? �?�?�?�??O4?�? HO6OlOZO�O~O�O�O��O�? O_ޣ8�INOT 2�8i�р�G;� O_a[��ο<�_J�f�0 �_�[ �O�_�O�_�_�_3o!o Wo=ogo�o{o�o�o�o �o�o�o/Se K�w����� ��+��O�a�G��� s�������ߏŏ���'�ĮEFPOS1� 1��  x�Ou�T�|_���� Θh�z���� �9� ԟ]������~���R� ۯv�����#�5�Я� �}�h���<�ſ`�� ���Ϻ�C�޿g�� �ϝ�8�Jτ�����	� ��-���Q���N߇�"� ��F���j����߲� ��M�8�q���0�� T��������7��� [�m���T������� t�����!��W�� {�:��p� �A�e � $��Z�~/� +/=/��$/�/p/�/ D/�/h/�/�/�/'?�/ K?�/o?
?�?�?@?R? �?�?�?O�?5O�?YO �?VO�O*O�ONO�OrO �O_�O�O�OU_@_y_ _�_8_�_\_�_�_�_ o�_?o�_couoo"o \o�o�o�o|o�o)��o&_�cK�2 1�W�M��� �o��7��4�m�� ��,���P�ُt����� ҏ3��W��{���� :���՟p�������� A�ܟ� �:������� Z��~�����=�د a����� ���D�V�h� ����'�¿K��o� 
�lϥ�@���d��ψ� ߬Ͼ���
�k�Vߏ� *߳�N���r����� 1���U���y��&�8� r����������?� ��<�u����4���X� ��|�������;&_ ����B��x �%�I�� B���b��/ �/E/�i//�/(/ �/L/^/p/�/?�//? �/S?�/w??t?�?H? �?l?�?�?O�?�?�? OsO^O�O2O�OVO�O zO�O_�O9_�O]_�Ox�_gyt3 1� ._@_z_�_�_o"_@o �_do�_ao�o5o�oYo �o}o�o�o�o�o` K��C�g� ��&��J��n�	� �-�g�ȏ��쏇�� ��4�Ϗ1�j����)� ��M�֟q�����ϟ0� �T��x����7��� үm��������>�ٯ ���7�������W�� {�ϟ��:�տ^��� ��Ϧ�A�S�eϟ� � ��$߿�H���l��i� ��=���a��߅��� �����h�S��'�� K���o���
���.��� R���v��#�5�o��� ��������<��9 r�1�U�y ���8#\�� �?��u�� "/�F/��/?/�/ �/�/_/�/�/?�/	? B?�/f??�?%?�?�_�T4 1�_[?m? �?%OOIOO?mOO�O ,O�O�ObO�O�O_�O 3_�O�O�O,_�_x_�_ L_�_p_�_�_�_/o�_ So�_woo�o6oHoZo �o�o�o�o=�oa �o^�2�V�z �����]�H��� ���@�ɏd�Ə���� #���G��k���*� d�ş��韄����1� ̟.�g����&���J� ӯn�����̯-��Q� �u����4���Ͽj� 󿎿ϲ�;�ֿ��� 4ϕπϹ�T���x�� ����7���[����� ��>�P�bߜ�����!� ��E���i��f��:� ��^���������� �e�P���$���H��� l�����+��O�� s 2l��� ��9�6o
��.�R��?�45 1��?���R/ =/v/|�/5/�/Y/�/ �/�/?�/<?�/`?�/ ??Y?�?�?�?y?O �?&O�?#O\O�?�OO �O?O�OcOuO�O�O"_ _F_�Oj__�_)_�_ �___�_�_o�_0o�_ �_�_)o�ouo�oIo�o mo�o�o�o,�oP�o t�3EW�� ���:��^��[� ��/���S�܏w� ��� ������Z�E�~���� =�Ɵa�ß���� ��� D�ߟh���'�a�¯ ��毁�
���.�ɯ+� d�����#���G�пk� }���ɿ*��N��r� ϖ�1ϓ���g��ϋ� ߯�8�������1ߒ� }߶�Q���u��ߙ��� 4���X���|���;� M�_���������B� ��f��c���7���[������ $6 1�/����j� ���b���!� E�i�(:L ���/�//�S/ �P/�/$/�/H/�/l/ �/�/�/�/�/O?:?s? ?�?2?�?V?�?�?�? O�?9O�?]O�?
OO VO�O�O�OvO�O�O#_ �O _Y_�O}__�_<_ �_`_r_�_�_o
oCo �_goo�o&o�o�o\o �o�o	�o-�o�o�o &�r�F�j� ��)��M��q�� ��0�B�T����ڏ� ��7�ҏ[���X���,� ��P�ٟt��������� ��W�B�{����:�ï ^����������A�ܯ e� ��$�^������ ~�Ϣ�+�ƿ(�a��� �� ϩ�D���h�zό� ��'��K���o�
ߓ� .ߐ���d��߈���x5�-7 1�8 ����.��������� ������N���r�� ��1���U�g�y��� ��8��\���} �Q�u��"� ��|g�;� _���/�B/� f//�/%/7/I/�/�/ �/?�/,?�/P?�/M? �?!?�?E?�?i?�?�? �?�?�?LO7OpOO�O /O�OSO�O�O�O_�O 6_�OZ_�O__S_�_ �_�_s_�_�_ o�_o Vo�_zoo�o9o�o]o oo�o�o@�od �o�#��Y�} ��*����#��� o���C�̏g������ &���J��n�	���-� ?�Q����ן���4� ϟX��U���)���M� ֯q����������T� ?�x����7���[��� ����ϵ�>�ٿb�H�Z�8 1�e��!� [��������!߼�E� ��B�{�ߟ�:���^� �߂ߔߦ���A�,�e�  ��$��H����~� ���+���O������ H�������h����� ��K��o
�. �Rdv��5 �Y�}z�N �r��/��� /y/d/�/8/�/\/�/ �/�/?�/??�/c?�/ �?"?4?F?�?�?�?O �?)O�?MO�?JO�OO �OBO�OfO�O�O�O�O �OI_4_m__�_,_�_ P_�_�_�_o�_3o�_ Wo�_ooPo�o�o�o po�o�o�oS�o w�6�Zl~ ���=��a����  �����V�ߏz���� '�ԏ� ���l��� @�ɟd�퟈��#����G��k����uχ�M�ASK 1���≢ӯ᧳�XNO�  ¯��MO�TE  ���8�_?CFG �?������A��*SY�STEM*7�V9.40107 ���7/23/202?1 A �q����z�REPOWE�R_T    $FLAGr��  ��STAR}T�� , ɶ�$DSB_SIG�NALr�$ײU�P_CND��7���RS232X���� � $COM�MENT �$DEVICEU�SE��PEE�$�PARITY��O�PBITS��FL�OWCONTRO~��TIMEOU*����CUS�M��AU�XT����INTE�RFAC8�TAT}UZ����CH�� t �$OLD_>�C�_SW �FR�EEFROMSI�Z��n�ARGET�_DIR 	�$UPDT_MA�P�¹�TSK_E;NB��EXP���ý!/�FAUL��E�V���RV_DA�TA��  �$3�Ep�  � 	�$VALUH� �	/�GRP_ �Ų3�  2 ��SC��
  �$ITP_E� $NUMc��OUPr���TOT�_AXZ���DSP���JOGLI��F?INE_PC)�y��OND��$��U�M��K��_MIR�����P6�TN�AsPL���_EX'��ԕф�������PG�<�BRKH�� �N�C��IS K� �c�TYP��n��P���D8��� �BSO�C��8�N��DUM�MY166��SV�_CODE_OP�v�SFSPD_O�VRDl�#�LDl����OR��TP ЋLE��Fd����O�V��SF�RUN����SF5�����U�FRAK�TOi�L�CHDLY��RE�COV�����WS0��������ROvæ����_5�   �@��SD�NVER]T��OFS��CP���FWD�������ENAB���TR�����_%�FDO> �MB_CM�� =B��BL_M����-32=�V�������BЋ��G.A�AM�?�! ��o��_M�E ��M��x��T$SCA�е Dj�� �HBK�����IOvv� �IDX�PPA�
�	������DVC_DBG��E ��F��@��]��g�]3e^��ATIOr��������UL�иy�A	B��۰Y���З�F��h����_����SU�BCPU���SICN_հW��1,�FWʲm�$HW_C1��"!� K&F�$AT��K��$/UNITw�q j ATTRI�~"���CYCL��NEC�A��FLTR_2_FI��������LP��CHK_n��SCT�F_j'cF_t,�"�*FS�Oo"CHA �(>18Nx�=2RSD��첰��
��� _TlP�RO�n�EMP�����k�T+2" K�x+2F �6DIAG �?RAILACS��M|�LO�����7&��PS��w� � �֮PRGS�� ���AC9+�	��F�UNCl���RINS_T����0<DFm�RAM@��l�� peC���eCWAR�~�CBLCURzHDA�K�!�H�HDA`u�fA�H�C�ELD�� ����C��oA�1�C�TI	BU��K�$?CE_RIA����+AF	 P�CS��IUT2�0C��f@�OIu DF_LaEc1����p�LMQ�FA��HRDYO,���RG�@H_0����@�UMULSE�P�'3nB$J���J����FAN?_ALMLV��a�WRNeHARDHw���$�P��p@2a�S���O�_����AU��R04��TO_SBR;�e�Ћjj ;|DA�cMPINF����!�d�A�cREG��C�V�����d�DgAL_��!�FLL%l�$M�@� ��fd� K�%h,uCM93NF�!�ON j!�e0�b/r8F�3�q� ���� ���$Y�r����z�d���$ ��4�EG7������qAR�й��2�3�u�@�A�AXE��ROBn��RED��WR��2h�_"���SYe��qtj�D�SN�WRI���vJ STڰ�Ӆ�i�J��El!M��t8��Dca��B����9�3.� OTO�aMЦ�ARY��̂�1�W����FIJ���$LwINK�QGTH�M�T_������s30���XYZ��8�"!/�OFF���)��ЀB��1B�q�������r�FI@� ��������1B��_J)�K������X`4����3F$6�|0��R��Cٰ0�DU����3�P�3TURB`XS3�ځ�bX]�� �FL�i���p�Q�5���34���� W1M�K��M�Ă!�5�5%	B'��ORQ�6��kC蘹��0
G�O@�N	B�ӵќ�a�OVE��rM ����s7��s7��r6����5���5���4�AN B!�7�IQ�q���v� fW�/��;����s��L[���ER��oA	�2!E��3�	C��A��o ��]E�2؇�A��AAX��K��A�S!� XŹ1d��Qdɋ�cʱ� cʹ�c��0cʞ�cʼ�c�1+�cƗP`ɗPp� �P�ɗP�ɗP�ɗP�� �P�ɗP�ɗP������x� �RC�DEBUB#$=AIc�2�����CAB�7����V� A" 
��n�q�� F �*� 狡 籡 � �� ��1 瞁 缁OTp��IR��r�LAB��q�> KGRO� 4�Bl� B_�1� z��3���`�������va��AND���� ����va"� �Jq���6��AE�� �NT8)`��h�VEL�1���r��1z���VP?Rr�NA`|�-�CS1�%���3񤞂  �SE�RVEh�p	 $�^�i@��!��P�O�BP_�0T �!	�򜱱p
 � $TRQ"�b
-� IR�2
0'P�0_ � l'@�Q�&ER	R���"I� v𒴃'TOQ����L�b�(j���0G��%�A���� �@  ,h��4N ��RA�? 2 d�+��'  �pa$+��2yPR� �OC�A=   }uCOUNT��� ΨpFZN_wCFG 4G �f�"TA�?#��ӡ�����e�s ���M �R�q����4� �FA6P��DV�X�����r����� �P?b�pH�ELpj� 5��B_BASNA�RSR�f%@��S1Q^ 1�^ 2��*3�*4�*5�*6ʁ*7�*8�Q!RO0�����NL�q��AB���0_ ACK���IN#T_uUpX`�Pya9_PU�,Cb*ROU��PM@�h�>#�z`|�>�TPF?WD_KAR��a&w RE���PP��Ab@QUE�i+���k�C`VaI`��>#�po3w��f�SEM���F
��PA�STYf 4SO�0ldDI,1�`���1=�wQ_TM>�cMANRQ]F��ENDjd$KEYSWITCHo3؄1?A�4HE�BE�ATM�3PE�pL�E��1��HU�3F��4�2SDDDO_H�OMGPO?a0EF��PRw��/�{�u�C�@O�Qt �OV�_MԒ��Ev�OC�M ��7
��q>$HK�q D��g�	Uo�2M�p�4W���FORC�cWARޚ���=%OM>�p  @�ԧ�*u`U��P�p1�V,p��T3�V4��(Oʔ0L�R��hUN�LOJ0mdEDZ[a 2NPZpSkw 0pADD���$SIZ�a�$VA���MUL�TIP2?c�PA��Q � $ Y9@`R���rS���yC� �fFRIFY"�#S�0�YT�`NF`DODBU]�G��e`�c�i��Fqw@IA��A����������P|_ �p � ]`ƠTEl�񢞃SG%LoqT��]�&��sx��F�ppSTMTj�ޡsPSEGn�BW<�qtSHOW�uZ!7BAN�pTPT���༄��+��J��SmV�_G� ���$PC��$�T�F�B�QP-�SP�0A�+0/��PVD���� �hA00��p��Pw��Pw��P�w��Pw�5u�6u�7�u�8u�9u�Au�B�u��Pw�|�x��pw�Fu���9���1��Gp9����1��11ω1�܉1�1��1�1��1�1*�17�2�t�2��2��2��2���2��22ω2�܉2�2��2�2��2�2*�27�3�t�3��3��3��3
��3��3��٨܉U3�3��3�3�U3�3*�37�4t�U4��4��4��4��U4��44ω4܉U4�4��4�4�U4�4*�47�5t�U5��5��5��5��U5��55ω5܉U5�5��5�5�U5�5*�57�6t�U6��6��6��6��U6��66ω6܉U6�6��6�6�U6�6*�67�7t�U7��7��7��7��U7��7��7ω7܉U7��7��7�7��7�7*�77��V�P�@U �! ��v"
���b��� x $TOR��1%p  ��M	 RXJ 1 +�Q_<R��P���P�SD�C�AY�s�_U�`~�R�YSL� �� � ]er{�dRg�@����@��4rVALU�{60�6F���F��IgD_L`CHI
�I�R$FILE_]36'$$S� ��{SA h�~b E_BLCK�3�o�qxD_CPU �	^`�	R`�9K3�YopW3R  � PW>� �`6�LA�qS�\��RUN8pG ���@6�6��HW0X�XqT�2�1_LI�R  w � G_O�2}�0P_EDI�Rf�T2�x!��i	0��`�`oABsUI���" $��91LINE�sIAG%_Njp�`�Q�{SC�P# �CLLS �PT�R!	�TBC2a�$ �fp{@8p9`��1xFTDH$CT#DC8u�c M�]&Ls!\'TH�`�Q�$�8�'R�!-`vPER�VEC�$C�$Hq�(!0�  %Xw -$�!LENC0�$C� :0RA�0+b&��W_T�1�!#M2)7MO�(eS�`ERTIAm�/Q9�!�� f;DEv5�aLgACE=RO�CC'co��@_MAC`u6�5�7�1TCV�<�1�7TiA�:�5�:M�t34��E�34�JPA0�MD@D�@J��_�t5aA
�5�!2P�pW�zAls3-`JK�FVK� �AOQ�AHq�@J��A��CJJ�CJJ�CAAL�C�@�C�@�FTq2�B5�#
@N1�<
P�;�0m��_�qp�@v(!CFGb& `�GROU���qr9��N? C�cePREQ�UIR�"`@EBU��c�!AF$Tv02�%�Q� �V(!F`.$'� \��APPR��PCLm�
$�NN�XCLO��YS%��Yt5
(!�f( �3 Mq �0	@R8d_MG.qB`Ca�c Lh�A@�0MgBRKKiN�OLDKf�pRTM!Ow�j{m<eJ�3P�D�0�C�0�C�0�C(�0 S�06�e7�e}q����!.$)� �R	2�(w�A6sPATH2wKqAsKq�8Gs(`�P(q��S�CA��g�RAaINF�"UCU0<1�pCO�KUM�xY+0� J@ �q�!�z�@�z�`�p�PAYLOA�gJ;2L��R_A���L� ���#�LeR_F2LSHR�$P�LO��qQ��s_�>�sACRL_!1�u����w�tRH��m��$HLb��FLEX��S�!J,&* P �R=/O/�/�/V܀�%+ :�/ 6�0 Q�h�?Q�0??0<F1h���ʗ??Q?c?u?�?�?��E�?�?�? �?�?�?O!O3OѨ� 5GLC�Dސ �TOfOxO$g�JT��ϡX{�ء �E=�%��E��x��O�O �O�@�E�E�E�E __�$_6YnBJIT, ��8 V_h_z_� ��A1T㖍Q?@ELQ��ԶXJ�P+�PJE�x`CTR�qޑTN��ƅWHAND_�VBm�ہ��t-��20Lf�$��S�Wۑ%#&f.� $$M5�9i6�hab�@warܔ�eնb��A  �<f��EmAVl��
hjAvkA�k��Wk� �hjDvkD�kPepGN�STjgV�wiV�N�hDY�PLf�� ���� G�h�G�b�� �G%���r��eP�e�e��e�e�e�eurrJ�-%/ X�=�0r ��T�
a`�ASYIMuu���Puv.K��}b��_W���p�t �m��)������J��`$�D:	C��_VI��
c� V_UN�� �ȳO�J�E���b�� y�����?@���`����G��̄ԃ "0 3HR��0"�uL�j"DI�`�SO�8 "vIS1 ذ��I��A�ay��������" p�w �2 � :�MEB9���D��T�PT' F�Rp!N�R�A�	 (2!&)T( �;Q $DUM�MY1�a$PS�_�RF��n$�m&2`FLAKPY�Pw��"#$GLB_T[Њ�% ��p;� ����3 X뀬�WqSTDA�PS�BR6M21_V��RT$SV_ERb5�O���# 3CL� ��"AR�O�qGLv� EWLQ4 4SP�!$Y�Z�WK3�@L�6�A��r%0�+3U155 C�N�e0- $GI���}$11 4�8+3d0LQ6 LSP�6���}$F��E�6NWEAR3�N�F�9�0�TANC�  ��JOG���` �79�$JOI�NT��J�Ο4MS�ETLQ8  �7E�5��S�5��LQ_9�  ��U9��?��PLOCK_�FOa�AѐBGL�V��GLHTES�T_XM�P>AEM�P@�R�B�"j@c$U1�02��25�P�d3�A6�B=�o@�A4��!CE8P�3�@ $�KAR��M�TP�DRA40T�1VE�Cy�V@IU�A7��AHEq@TOOL���=SV��REPI�S3)�]R6�a�ASCH$@�P8JQO�p�#\$3Oq�0SI��R  @$RAIL_BOXE���0ROBO�D?��1HOWWAR�Q�Qj �QROLM u"�UE��T�Ru��PҐnpO_Fv�!0�HTML5��q���" ���P+2wQq:T
NoR"POC�;
BȢ�A`�-1OUN&B< t0�E4���j@�bPOsa.��PIP�FN1�SR��RwQ��AJ`.�CORDEDo@{pi`�0SXT�`�1)F�Pq��O� = D � OB�ѿ�o@w�qV#� r����SYSqADR�q �TCH� > M,C�ENz��AvAE_�4ttN�7�
q�VWVA�? Ǥ P12�PR�EV_RT��$�EDIT�vVSHWRv��&�p1�E1%� D����tȱ?$HEADA4	��sKEE1P �CPSPD �JM%P$pL�@�R5���@p�lvI�@S��C�NEFP����OTICK��"M���:�J�HN�!A� @pg�R�(�_GqP���V��STYnr�QLO�!�J���E��B�`
�pGzu%$ԙq�4=� S��!�$���!�%��&P��SQUP���"��TERC ���{TS`�C �0�� s�1�r��4Q��O 
#�IZ�$�1�%i!PR�`v!Ւc��`PU��_DO��2spXS"@K�A�XI�c�AUR ��R����P��2v1я�Y_4PDrETE�PxB@ pz��p`{��A��V}�]$9�W2ر�nSR�Dl��[ْ�j���}�ҩ ��������������� ���������2�(��V�f�6�C��D�C�U���*�!SS}C�  E h0cDSŀQ\ SP�&2�AT�Б�摤��s�Y"ADDRESzGSB�pSHIFIB^�A_2CH�.q�I� ���TU� I�o� F
BCUSSTOf���VTBI�AGer�HF�ɓ_�
�J�
 0����H \Y��h���̣�Z��C'㦒i��˜e2���TXSCREE�	rI��TIN!A#3�0dԆ4zaF�F�J�J TY�0ɒ Dq1� ���Cr����pRRO���0������  �UE�O�K �r�]q{ S�$1DqRSM���U`�`o���uS_^3�;��+�>�Y��F�CxdB�� 2J�pUEF�L�2~�ՐWGMTL�!��� �aXa��BBL_r�PWC �M ��j��OX1��LEv����P����RIGH���BRD4l�CKGRC #�T�`"��WIDTH�S�p���Q�!GQ��UI�`EY-`�N d�<0"`�P炧PёB�ACK�u"��1��FO�a��LAB��?(�I�PhBg$UR�Q��MEn���H�� O 8�V�0_������R@E0jB���X����O}�J�P�� 7�U�rGRxB�QLUMG)�f�ERV�a)0o�P�0v�Q�z�G�E���1d��b�LP$�o�El���)������qP�	5�6
�7�8�j���АP�0%�[&qQbASZ��Pn�USR14'R <Y��U�2���2FO���2PRI₡m�P���TRI�P�Qm�UND-ON�S�0(���
��Q	�. �AC�=� �T��cԑG ��T`居��OS:!&RI����CQ��U:?L3S>+"Ǆ�U���V4/F/T�ƅN�OFF�@60W)�%\#O� �@U�`�$Z�$V�`GU>qP�!�Vb�#��'��SUB�ǂ �E_EXeENpVb��WOۡ� X{ ��WQA�pc&1�@b�V_DBE3]0Ac	T- ��Y���1`��sOR�P�5RAU��"�4T�9jws1_�pO��Z | jxOWN|�{t$SRC���c�&�D�@�5��MP�FIބ�E�ESP ᑬ�|�UUv�QrcRp��2�p��[ `} �32{t��J�COP&�!$:��_@��0�A�a�EO2CT5�31AC31OC ��p�R��� \��SHAD�OW&�GS�A_UN�SCA&S�C[��CD�GD|QqEGAC��C���@C�Ct#]�� �R=q4�$5PER��J\H��S� C�`JUDRIVǖP�_V��mT����PDDMY_UBYCRT
�+#4���I��|��q�XOA�RP_h�@ބ�RL�BM��$r�DEYosE�X�`�ӒEMU>�X��=d0�USB�0��_Rzч"����҈!}Gw�PACIN��1�RGAvd�b�#�b0Q#�bc�AREz��+!�"/S�b�p^ )��y@G�PPG��`$��0SR �p_~�@ ���d�2	�B�RE6IcSW�`_A�a� I>cӐOYl�A~�Es��E��U�� �!Y��0SHK��`= �]z]���Bp�ЎsEA���w30�0Eu��0R�MRCV��a ��� O�M�0CH�	p�r�#�c�rREF�� �v�v�q4p� s�ph �z-��z-��{O��v�A_�0�z���{@�S1�5g�S�����v��b ��!`��ri�t�U��OU0�N��bL�RS� ]�e�2^`��e�'�Ԑ��_Eð���f�UL���`F@CO� a/`,�NTACn�OBm� (y�Py�8�L�S����S��(��P�V�IA26c ���HyD����$JO/����$Z_USPL���Z�W�pڑ7���_LI�$EP,�#��� ڑX�_�t_�mِDR���d 5E�P�AP� E�CACHSLO!�����0`Х�k�@CC0�MIw�F/�ѥT�Ц���$HO�0�2��C'OMMhS�O����d�A��@V�P�b+pT�_SIZS^�Zp`Y��Z�O1v6�MP~�FAI�5G�t��AD���B�MRE�βc�GP��%`@�FASYN�BUF�FVRTD� ��c�6�OL�D�_�#(�WQ#PC_��PUc��Qbp�EwCCU�hVEM�`x��p�ϧVIRC��� ����_DEL�A�cA���TAG:�R2aXYZ]�E�2aWq����ă��T5PbIM��ƨ�|k ĥGRABB(!�YIcNpLERW`C!���F_D�PY�A5��b֪�c�n�r��e�Ѣ�LASx�\Yqn�_GEu�f�A��"���T�A5QG@Q�eI�Կb�ƀP�BG��V��QPK��`��v��GI��N��Gr~ �Ѡ�۱��Ig���Sа��Ne���L"1v�h�B�3{"PB5�J�I&`�A ���@��d�sH��@��@�"io����!TP�YiAD���a�T��j $>1IT�0n��U�-C�"VSF|@�3k�  �B[y���URl�s�`SM�l���8ADJ0�5eؐZ�Di�m D��)�A�L�Ͱ� (�PER�I^�$MSG_Q �$d����pO2���n�M��1��#^��XVR�o�Ҿ�T_OVR��
_�ZABCz5p�b�f���
֑��AC�TVS:� q �� $����CgTIVB�IO�R���QIT(S�bD�V'@
�av��04��A� PS�B� ǳB����L�STR�̐ �/_�S�Ak���DCwSCH�2r L�1 S���@#P��c�GNA�'5c�R�_FUN��	 '�Z� Js[�$W�$L�R�I�Z/MPCFz5ts��phA��QLNK�"�
 ���{4u� $��p�CM+CM~`C�CCzA-!��P� $	JK#E$DI�Q"b"[' O@g%O@E'�p�t`"�'sUX���UXEDa �&��V%�%l%�!�!�)8�!�'J FTFZ�Q#�4Yq	�Z�vC ���ˁ$2Y1�}D:� w 8�p�R��U�A$HEgIGHwcM�?(4��:��`%0քx g� ,G�$B8�x_@UjBSHIF��58RV0�F����2[ C�F"zAK�-@bb �1 ��C>�DH5�CEhV��$1S�PHER�P y� ,4�`8v?�9��`�PLc`N���A � ������A�BOWER� �B�A�@�FS�M_DRY>�%�E�B%��A�O�M�Bd�`��N�JUM<�O�O�OY_�D����i�G�]S�IGSPD=�}�|X�X��_�ZR��_�Fې[��CփQ�C�QNG�e�z� :Y�H_�II_AIRP�U�`  :Z  :oa^r����@\k�  �@�ISO�LC  �lkb@�ala�A�!k�0o�JOB�Tf�g�Cjc�@;Cts#���?�HhaH844  t�~��y�@E����Oxރ@S232u� 1��E�S L�TE�� PEND�AN�ps�a�a��|�oB@Ma�intenanc�e Cons0���0�"*�<�No Use�Z� �~�@������Ə�B�rN���r�a
e�qCH�O� �m�A		�I��!UD1�:o��RSMAV���? e�EaSR  \kt �A���̐��TVv� e���I���^��V  �2dv�Q� D�P ���q�\��� ���E��§���Я� ��*��:�<�N���r� ����̿���޿ �&� �J�8�n�\ϒπϢ� �϶��������4�"� X�F�hߎ�|߲ߠ��� ������
���T�B� x�f���������� ����>�,�b�P�r� t��������������(8^L��A��$SAF_DO_PULS�pCq�C�QsSCAN� e�F�@SC�@)��*ШQ�
@�a�d�qY�Y���� ��4FXj|� �����/�+��25$�@)d5$P!���) @�b{/�/�/�/�d)x/ Z��$�/_ @�#T`�/�?!?3?@9T D��@?i?{?�?�?�? �?�?�?�?OO/OAO�SOeOwO�O��v)��O�O�O�G { 
�;�o�D�Q�ap�U
�u��Di�~�J0 � ��j �w_�_�_�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o �������� �#�5�G����/p� ��������ʏ܏� � O�#%,�>�P�b�t����������Οӑ��0 ]RZS(Ud]�1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ�������Z��%� 7�I�[�m�ߑߣߵ�  ��������!�3�E� W�i�ԟ��3"��� ��������'�9�K� ]�o�}����������� ���� 2DVh z������� 
.@Rdv��OO3���� �//*/</N/`/r/��/�/�/�/�/�/�*p��/"?,6��iR�?�M	123�45678ARh�!B!�� )���P�? �?�?�?�?�?�?O"O (A�KO]OoO�O�O�O �O�O�O�O�O_#_5_ G_Y_k_|]:O�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o~_�_ �o+=Oas �������� ��o9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�*������� şן�����1�C� U�g�y����������� ���	��-�?�Q�c� u���������Ͽ�� ��֯;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�,ϑߣ� �����������!�3� E�W�i�{������"���6��������.�@�\:Cz  �B\�   ��M�2� }��M�
���  	�������������
��� ��Pbt���� ���(:L ^p���5�� � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?a5:2��:K2<]4 S5��?  �m;�?�q�s�j2���t C t�9�?��(�3 `:2j2�? Og�s��.�$SCR_G�RP 1*+�*4� �� ��� �F5	 ^A�fBwBpD�1L3��OG�G�O�O�OP������BDE� DP� }CW�K.�ARC Ma�te 120iC� 67890���M-VPA 8���M2IAZQ�C
�12345[T�FfO2  x0�� �VfA�FUA�CUA.\1"�AtJ�A�Y	�Ro�o(o:oLo\l�G�H�f@�TjGUB �o�O�o�o�o�F��с�o�o=C8/{hjGxxl`X�IB�c�!ƈ�r�t�AAt��  @ �u�A@���p� ?��w�rH�c���z�AF@ F�`)�1�(U�@� y�d�������ӏ���� z}�q�r"���1�C�B�Q�揗������� ߟʟܟ� �9�$�]� H�����-�C�O��دF7��կ
���q�qO6����G@�p4J�c��`��W�\�C���A�p��õ$�o�eа.Ĳ��A ���-���BȸN�`�/� P��( �Ϥ϶�y������ς�J_�T�;��S��5@ECLVL  ������RѰQ�@N�L_DEFA�ULTV�J��� j�HOT�STRv�ѱ��MI�POWERFU��X�����WFDO�w� ��4AERV?ENT 1	]�]���� L!DU�M_EIP����j!AF_IN�Ev�;�C�!FT$�j�1��!�o��� �}���!RPC_MAIN������&���VIS�����r�!O�PCUAs����a���!TP��P�U��$�d��
!
�PMON_PROXY'�e��V���$ �fE�!R?DM_SRV�$�9g��!R�T
�%�h�:!
��M�m!�i)�!R�LSYNC���8u�!ROS����4�/!
�CE��MTCOMd/'�k/j/!	3"OCONSk/&�lY/��/!3"WASR�C�'�m�/?!N3"USB?%�n�/>N?!STM��h?#�o=?�?��?��?��=��ICE_KL� ?%�� (%�SVCPRG1��?/JE2/O4O@3�WO\O@4O�O@5��O�O@6�O�O@7@�O�O@wT?_:L9G_L[Dt_A!O�_ AIO�_AqO�_A�O oA�O<oA�OdoA _�oA9_�oAa_�o FA�_FA�_,FA�_ TFAo|FA*o�FA Ro�FAzo�FA�o� FA�oD�FA�ol�nA �?�2@O@����>A  �$��H�3�l�W��� {���Ɵ���՟��� 2��V�A�h���w��� ��ԯ������.�� R�=�v�a��������� п��߿��<�'�`� KτϖρϺϥ����� ���&��8�\�G߀���:_DEV ~���MC:���4����GRP� 2�Ֆ�@b�x 	� 
 ,�����	���,� �P�7�I��m��� ���������(�:�!� ^�E������߸�o��� ������6H/l S�w�����  D��9z1 �������/ .//R/9/v/�/o/�/ �/�/�/�/?]*?<? #?`?G?�?k?}?�?�? �?�?OO�?8OO\O nOUO�OyO�O�O?�O �O_"_	_F_-_j_|_ c_�_�_�_�_�_�_�_ ooBoTo;oxo�Omo �oeo�o�o�o�o, PbI�m�� ������:��o ^�p�W���{������� �Տ���6�H�/�l� S�������Ɵ����� S� �ןD�V�=�z�a� ������ԯ����߯� .��R�9�v���o��� ���⿙���*�<� #�`�Gτϖ�}Ϻϡ� ���������8��1�\n�u�d �u�	\� �ߐ��ߴ������ ��%� �E�L����^�
�^�n�|�f�� ���������2��Z� ��D�2�h�V�x�z��� �����(���
@ .dRt�����  ���<*` ���P�L�� �//8/z_/�(/ �/�/�/�/�/�/�/? R/7?v/ ?j?X?�?|? �?�?�?�?*?ON?�? BO0OfOTO�OxO�O�? �O�O�O�O�O_>_,_ b_P_�_�O�_�Ov_�_ �_�_�_o:o(o^o�_ �o�_No�o�o�o�o�o �o 6xo]�o&� ~�����>d 5�t�h�V���z��� ��ԏ���:�ď.��� >�d�R���v����ӟ ������*��:�`� N���Ɵ���t�ޯ̯ ��&��6�\����� ¯L�����ڿȿ��� "�d�I�[��4��|� �Ϡ�������<�!�`� ��T�B�d�f�x߮ߜ� �����8���,��P� >�`�b�t������� �����(��L�:�\� ������������  ��$H��o��8 �4�����  bG�zh�� ����:/^� R/@/v/d/�/�/�/�/ /�/6/�/*??N?<? r?`?�?�/�?�?�?�? �?�?&OOJO8OnO�? �O�?^O�O�O�O�O�O "__F_�Om_�O6_�_ �_�_�_�_�_�_o`_ Eo�_oxofo�o�o�o �o�o&oLo\o�oP >tb����o� "���&�L�:�p� ^����������܏ � �"�H�6�l����� ҏ\�Ɵ���؟��� �D���k���4����� ¯���ԯ
�L�1�C� �����d��������� �$�	�H�ҿ<�*�L� N�`ϖτϺ����� � ����8�&�H�J�\� ���Ϲ��ς������ ��4�"�D���ߑ��� j�����������0� r�W��� �������� ������J�/n��� bP�t���� "F�:(^L �p����� / /6/$/Z/H/~/� �/�/n/�/j/�/?�/ 2? ?V?�/}?�/F?�? �?�?�?�?
O�?.Op? UO�?O�OvO�O�O�O �O�O_HO-_lO�O`_ N_�_r_�_�_�__4_ oD_�_8o&o\oJo�o no�o�_�o
o�o�o�o 4"XF|�o� �ol����
�0� �T��{��D����� ҏ������,�n�S� �����t�����Ο�� �4��+���ޟL� ��p�����ʯ��0� ��$��4�6�H�~�l� ���ɿ������ � �0�2�D�zϼ���� j����������
�,� �Ϩ�y߸�R߬ߚ��� �������Z�?�~�� r���������� 2��V���J�8�n�\� ~�������
���.��� "F4jXz� ������ B0f���Vx R���//>/� e/�./�/�/�/�/�/ �/�/?X/=?|/?p? ^?�?�?�?�?�?�?0? OT?�?HO6OlOZO�O ~O�O�?O�O,O�O _ _D_2_h_V_�_�O�_ �O|_�_x_�_o
o@o .odo�_�o�_To�o�o �o�o�o<~oc �o,������ ��V;�z�n�\� ��������ڏ��� ʏ�Ə4�j�X���|� ���ٟ������� �0�f�T���̟��� z��ү�����,� b�����ȯR������ ο���j���aϠ� :ϔςϸϦ����� � B�'�f���Z���jߐ� ~ߴߢ������>��� 2� �V�D�f��z�� ������
���.�� R�@�b��������x� ������*N�� u�>`:��� �&hM�� n������@ %/d�X/F/|/j/�/ �/�/�//�/</�/0? ?T?B?x?f?�?�/? �??�?O�?,OOPO >OtO�?�O�?dO�O`O �O_�O(__L_�Os_ �O<_�_�_�_�_�_ o �_$of_Ko�_o~olo �o�o�o�o�o�o>o# bo�oVDzh�� ������� R�@�v�d������ � �������N�<� r�����؏b�̟��� ޟ ���J���q��� :�����ȯ���گ�� R�x�I���"�|�j��� ��Ŀ���*��N�ؿ B�ԿR�x�fϜϊ��� ���&ϰ���>�,� N�t�bߘ��Ͽ��ψ� ������:�(�J�p� �ߗ���`�������� � �6�x�]�o�&�H� "�����������P��5t�}��$SER�V_MAIL  �~�t �ZOU�TPUTi��@^RV �2��  w  �(D�^SAV�E�x	TOP10� 2�	 d z�0BTfx� ������// ,/>/P/b/t/�/�/�/ �/�/�/�/??(?:? L?^?p?�?�?�?�?�?��?�? OO$O��Y�P�[FZN_C�FG ���w���dAGR�P 2nG� ?,B   A�@}�D;� B�@��  B4�R�B21�HELL�gB���� ���G_&[%RSR &_'_9_r_]_�_�_�_ �_�_�_�_o�_8o#o�\oGo�o�o�n�  �tb�o�o�o�b�o ��orpS��g�b2�d�l��mOr�FHK 1�K ��� �����(�#�5� G�p�k�}�������ŏ�׏�LOMM ��O'��BFTOV_�ENBi��grO�W_REG_UI�G�\IMIOFW�DL���E|�WAITD�Hy�B��� h����TIMnh���۟VAh |��|�_UNITC����	LCa�TRY�h��^ MON�_ALIAS ?5e�� he/�� ����̯ڪ�����!� 3�ޯW�i�{�����J� ÿտ���϶�/�A� S�e�w�"ϛϭϿ��� |�����+�=���a� s߅ߗߩ�T������� ����9�K�]�o�� ,����������� #�5�G���k�}����� ��^��������� CUgy$��� ���	-?Q �u����h� �//)/�M/_/q/ �/./�/�/�/�/�/�/ ?%?7?I?[???�? �?�?�?r?�?�?O!O �?2OWOiO{O�O8O�O �O�O�O�O�O_/_A_ S_e__�_�_�_�_�_ |_�_oo+o�_Ooao so�o�oBo�o�o�o�o �o'9K]o ����t��� #�5��Y�k�}����� L�ŏ׏������1� C�U�g�y�$������� ӟ~���	��-�?���c�u����������$�SMON_DEF�PROG &����ա� &*SYST�EM*����$SP�D_LĤRECA�LL ?}թ ( �}��A�S�e�w����� /���ҿ� ���ϭ�>�P�b�t� �Ϙ�+ϼ�������� ߩ�:�L�^�p߂ߔ� '߸������� ����+copy mc�:diocfgs�v.io md:�=>192.16�8.56.1:24292�m������51�frs:o�rderfil.�dat virt:\temp\H�Z�������-��*.d������p��������xyzrate 11J�\�Q�c������8����mpbackI���w܉� }/1�db9�*FXa�6��3x1:\�;��� �v����41a9K�f�	/ /.@��u/�/�/ �G/�b/�/??* ��`q?�?�?�9? K?��?OO&/8/�/ \/mOO�O�/�/QO�/ �O�O_"?4?�?X?i_ {_�_�?�?C_�?h_�_ o�_0OBO�O�_wo�o �o�OIo�Odo�o ,_�_�ob_s���_ ;M�_���(o:o �o^oo������o�oS� �o����$6�Z k�}�����E��� ��� �2�D�ҟ�y� �����K�ԏf���	� �.���ίd�u����� ��=�O�����*� <�ů`�qσϕϨ��� U�ޯ����&�8�˿ \�m�ߑߤ���G�ڿ �����"�4Ͻ���i� {��ϲ�M���h�������$SNPX�_ASG 2����<���  0+�%���d�  ?�-�PARAM <�{F� �	R��Pg�+�g����� ��/�OF�T_KB_CFG�  )�B�,�OP�IN_SIM  <���#5�?/�RVNORDY_DO  �����QQSTP_DSB����$��SR <� G� &������=�/�TOP_ON�_ERR^-�P_TN <�6��A RIN�G_PRMpV�CNT_GP 2�<���I�x 	 ��+�~���(��VDeRP 1�����<�/(/ :/L/^/�/�/�/�/�/ �/�/�/ ??$?K?H? Z?l?~?�?�?�?�?�? �?OO O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oco`oro�o�o�o �o�o�o�o)&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�{�x� ��������ҟ���� �A�>�P�b�t����� ����ί����(� :�L�^�p�������Ϳ ʿܿ� ��$�6�H� Z�lϓϐϢϴ���������PRG_CO7UNT���6�'ENBK�M;����H�_UPD 1>�T  
��)� �ߤ߶���������'� "�4�F�o�j�|��� ������������G� B�T�f����������� ������,>g bt������ �?:L^� �������/ /$/6/_/Z/l/~/�/ �/�/�/�/�/�/?7? 2?D?V??z?�?�?�? �?�?�?O
OO.OWO ROdOvO�O�O�O�O�O��O�O_/_*_<_�_INFO 1���fЈP	 �__�_�_�_�Y@(���@^.D??�¾q��_�_�oo=oEd D���TRD�  C4  ´Pobm�YSDEBUG �ʁ��VPdiّ`SP�_PASS �B�?�kLOG �}V��  VP�Eh\_  �e�VQ?UD1:\�dc^�b_MPC�m��Q$c��q� ��1v?SAV �i/Ѱ1a�ar�uxS�V({TEM_TI_ME 1�g�� 0VP��t	���&}TMEMBK  ��e��`�oe��w���X|f��3 @��TSЩ�Ώ�ތ������a 1k@�G�Y�k�}� 0o����şן���TS xc�+�=�O�a�s�����������eů��� � �2�D�V�h�z��� ����¿Կ���
��.�@��uSK<�A�+�`P��ϒϤϘ�=VP"C���b�A�����  ��&�8�h�zߌ߀���VQ� ������� ����5��ʀB�g� y����VP$���� ˯����1�C�U�g� y����������������	-?QE�T1�SVGUNSPD��e '�e�t 2�MODE_LIMG  �y�bp2} �!�moABU�I_EDIT �"��SCRN �#�m�SK_?OPTION�`D���a�_DI�`ENB  �ţe>�BC2_GRP 2$cţc���Qx`�C��hBCCF�G &m�| ���`�$o!/ /1/W/B/{/f/�/�/ �/�/�/�/�/??A? ,?e?P?�?t?�?�?�? �?�?O�?+OOOOaOiDLL{OMO�O�O;O �O�O�O__>_�~^_ F�3Pf_�_z_�_�_�_ �_�_�_o
ooRo@o vodo�o�o�o�o�o�o �o<*`Np r���x�@��� �"��F�4�V�|�j� ����ď���֏��� 0��@�B�T���x��� ��ҟ������,�� P�>�t�b��������� ������.�@�^� p��� �������ܿʿ  ��$��H�6�l�Z� ��~ϠϢϴ������ ��2� �V�D�fߌ�z� �ߞ����������
� �R�@�v�,����� ����`�����<�*� `�r���R��������� ���� J8n \������� �4"XFhj |������ // 0/B/�f/T/v/�/�/ �/�/�/�/?�/,?? P?>?`?b?t?�?�?�? �?�?�?OO&OLO:O pO^O�O�O�O�O�O�O �O_ _6_�N_`_~_ �_�_ _�_�_�_�_�_  o2oDoohoVo�ozo �o�o�o�o�o
�o. R@vd��� ������(�*� <�r�`���L_����ޏ �����&��6�\�J� ������r�ȟ���ڟ ��� �"�4�j�X��� |�����֯į���� 0��T�B�x�f����� ��ҿ������� �>� P�b�࿆�tϖϼϪ���������$TBC�SG_GRP 2�'��� � ��� 
 ?�  )�;�%�_� I߃�m�߹ߣ�������	�)�d �� |�?��	 H�C���>���n:��ff��C�L���!�X�d�.�33���C�L�d�f�x0�&�&�>���F�e\L�Ȭ���BL���B$��9���(����L�^�p���  @ ������������0�M*x��?3�33~�	V�3.00!�	mw2ia�	*� �������� ��(��z	 &�'_   nB �X\n�J2	�*����CFG -,��� Ц���<���!//*��//U/@/ y/d/�/�/�/�/�/�/ �/????*?c?N?�? r?�?�?�?�?�?O�? )OOMO8OJO�OnO�O �O�O�O!�;��O�O_ �O?_*_O_u_`_�_�_ �_�_�_�_oo�_;o &o_oJooo�o���Ϻo ���o�o�o8& \J�n���� ���"��2�4�F� |�j�����ď���֏ ����B�0�f�x�8� ����L��ҟ��� ,��P�>�`������� h�����ί��(�:� L�^����p������� ��ʿ ��$��H�6� l�Z�|Ϣϐ��ϴ��� ������ �2�h�V� ��z߰ߞ�������
� ��"�4�F���v�d�� �����������*� <�N��r�`������� �������� &J 8n\����� ���4"XF h�|����� �
///T/B/x/f/ �/�/X��/�/�/�/? ?>?,?b?P?r?t?�? �?�?�?�?�?OO:O (O^OpO�O�ONO�O�O �O�O�O_ _6_$_Z_ H_~_l_�_�_�_�_�_ �_�_ ooDo2oTozo ho�o�o�o�o�o�o�o �o
@�/Xj|& �������*� �N�`�r���B����� ̏��܏��&���� \�J���n�����ȟ�� ؟���"��F�4�j� X�z�|���į���֯ ���0��@�f�T��� x�����ҿ俎��� �ʿP�>�t�bϘφ� ���ϼ��������� L�:�p�^ߔߦ߸��� �������� ��H�6� l�Z��~������� �����2� �V�D�f� h�z������������� 
,R@v�"� ��\��� <*`N���� x����/8/J/ \/n/(/�/�/�/�/�/ �/�/�/�/4?"?X?F? |?j?�?�?�?�?�?�? �?OOBO0OROTOfO �O�O�O�O�O�O__ �2_D_V_ _�_t_�_ �_�_�_�_o�_(o:o Lo^oo�opo�o�o�oδn  �`�c ��f�b�$TB�JOP_GRP �2-�e��  ?��f	� r's/.|��`�X8  ��rrDt  � �� � l�r�c �@�`?r	 �C�� �vf  Cq�w?q�rL���vp�q�q�u�qz��q�>�=�Z�C��p�p��p���C�  B��w�"��~�@w�v��X�333T��x�p=_�7LC�f��Z��D�p	����C��pŅA��r>�33����s��y<��G�C\�t��pC�#CH��?�
�LR�ԁD�qڌ��x�t��x~@p<X��B$�s@�q�����ßF�X�pڌ���� �������p?�ffC���[�ޟ�r�����'g�Ҩ���@Y�@pB�֣߯񯔝4�� "��>�H�y�T�f��� ����οؿ	����(�@B�,�^�hϙ�,���f����u	V3.�00Esm2iaDt*��Dt�a����� E�'E��i�FT�F�"wqF>��F�Z� Fv�RF��~MF��F����F��=F����F�ъF���3F���F��{G
G�dG�G�#
�D���E'
EMK�E���E�ɑ�E�ۘE���E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F��v�F�u�<#�
/<t�����0�Q�o�����f���?逘v�}ESTPARS���h9ps�HRO�ABLE �10.y���dD*�� hP��*�*�*��g�a*�	*�
�*�*���a*��*�*���i�RDIq�8q���������J�OR�d�n�����H����j�SP�6s � w������� +=Oas� ����}O S7r ��)��	-��������!�3�j��NUoM  �e8q�p�` ����j�_CFG 1�+�#�q@ pIMEBF_TTU�%6sb��6VER�� !56�3R 12y� �8���b�`�1 �`/  z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O_ �O�O=__*_@_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o5 "8FXj|�J�Rb1_�!L6@V5L�MI_CHAN+7� V5 �sDBGL�Vu�-5V5K��pE�THERAD ?UY�O������h�z�D��pROUmTI0!��!���̏��SNMASK�D�V3U�255.�
�����,���L�O�OLOFS_DI�U��u.�ORQC?TRL 3i;���ߪ�T��Ο���� �(�:�L�^�p����� ����ʯܯ�����!���E�I�PE_DE�TAI"�o�PGL�_CONFIG �9�)�!��/�cell/$CID$/grp1I�@��ѿ���Ͻ󀕏 2�D�V�h�zό�ϰ� ��������
ߙ�.�@� R�d�v߈��)߾��� �������<�N�`� r���%�������� �����J�\�n�������.}9��������"4�!6�\;� 8�������2� !3EWi�� �������/ //A/S/e/w//�/�/ �/�/�/�/�/?+?=? O?a?s?�??�?�?�? �?�?O�?'O9OKO]O oO�OO�O�O�O�O�O �O_�O5_G_Y_k_}_ �__�_�_�_�_�_o �_1oCoUogoyo�o�o����User� View ��}�}1234567890�o�o�o`(0t�p��P���i2�i-o������K]�b3u:�L��^�p��������c~4 )�� ��$�6�H���i�c~5ݏ����Ɵ؟ ���[��c~6��V� h�z��������ѯc~7E�
��.�@�R�d�ï��c~8����п������w�9�?� �lCamera�j��~ϐϢϴ����϶�Eq���&� �o@�R�d�v߈ߚߐ�  X�tym������  �2�D���h�z���߀����������
�1�� X�(���V�h�z����� ��W�������C�. @Rdv�/�܉ ����
��@ Rd������ ��/���{0/B/T/ f/x/�/1�/�/�// �/??,?>?P?�Y� D��/�?�?�?�?�?�? �/O*O<O�?`OrO�O �O�O�Oa?/���QO_ _*_<_N_`_O�_�_ �_�O�_�_�_oo&o �O/����_ro�o�o�o �o�os_�o_o8�J\n��9oKg9 ���	��-��o >�c�u�������ϏP�����	Z�0�� @�R�d�v�����A��� П⟉���*�<�N� `���_�a����˯ ݯ�����7�I�[� ���������ǿٿ�� Z���p�%�7�I�[�m� �&��ϵ�������� �!�3�E��&�9��� �ߣߵ������ߒ�� !�3�~�W�i�{��� ��X�jեH����!� 3�E�W���{������� ����������j� +��i{���� j���V/AS ew�0j�}; � ��////�S/e/ w/��/�/�/�/�/�/�  �$?6? H?Z?l?~?�?�?�?�?<�?�;   �/?  O2ODOVOhOzO�O�O �O�O�O�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\�<�  
�(  }�0( 	 l �������� � �2�h�V���z���:vz
J �D/�� ���/=�O�a�s��� ������ӟ�,�	� �-�?�Q�c������� ���ϯ����)� p�M�_�q��������� ˿ݿ�6�H�%�7�I� ��m�ϑϣϵ���� �����V�3�E�W�i� {ߍ��ϱ�������� ��/�A�S�߬߉� ������������� +�r�O�a�s������ ��������8�'9 ��]o������ ��X5GY k}����� �//1/C/U/�y/ �/�/��/�/�/�/	? ?b/t/Q?c?u?�/�? �?�?�?�?�?:?O)O ;O�?_OqO�O�O�O�O  O�O�O_HO%_7_I_�[_m__�O��@  �R�_�_�_�S�W�p���)frh:\�tpgl\rob�ots\m20i�a\arc_ma�te_1`c.xml�_6oHoZolo~o��o�o�o�o�o�h�� �o	-?Qcu ������o�� �)�;�M�_�q����� ����ˏ�܏��%� 7�I�[�m�������� ǟޏ؟���!�3�E� W�i�{�������ïڟ ԯ����/�A�S�e� w���������֯п�� ��+�=�O�a�sυ� �ϩϻ�ҿ������ '�9�K�]�o߁ߓߥ������X!Q |�_�P<< �P ?�������&� T�:�\��p����� ��������>�$�V�@t�Z�l������F�@�(�$TPGL_�OUTPUT �<�A�A�� ��#5GY k}������ �1CUgy�������Є��2�345678901���
//./6# �B�]/o/�/�/�/�/ O/�/�/�/?#?5?�*}??g?y?�?�?�?G? Y?�?�?	OO-O?O�? MOuO�O�O�O�OUO�O �O__)_;_�O�Oq_ �_�_�_�_�_c_�_o o%o7oIo�_Woo�o �o�o�o_oqo�o! 3EW�oe��� ��m���/�A� S�����������я �{���+�=�O�a� ��o�������͟ߟw�~�� $$�� �'��G�9�k�]��� ������ׯɯ���� �C�5�g�Y���}��� ��ӿſ�����?�}��Y�k�}Ϗϡϳ����@�������� ( 	 A�/�� S�A�w�eߛ߉߫߭� ��������=�+�a� O�q��������� �����'�]�K������  <<4϶��� ���� ��%7���hz ������V� .�dvP�� 
��|�/*// N/`/�H/�/�/B/�/ �/�/�/?r/�/J?\? �/d?�?l?~?�?�?8? �?O�?�?FO O2O|O �O�?�O�O^O�O�O_ �O0_B_�O*_x_�_$_ �_�_�_�_�_T_�_,o >o�_botoNo`o�oo o�o�o�o�o( ^p�ot�@�� ���$���Z�� F�����|�Ə؏6��� � ���D�V�0�b��� ���ԟn�ܟ
�� ��@�R���v���"�t�������������)�WGL1.XML���;��$TPOF?F_LIM ��������I�Nw_SVQ�  ���c�P_MON �=��e������2E�STRTC�HK >��c��V�L�VTCOMP�ATx��g�VWV_AR ?��%�.|� ٿ =������M�_DEFPROG %ǹ�%Tϛ�J�_DISPLAYX�Ǿm��INST_MSK�  �� ��I�NUSER����L�CK���QUIC�KMEN%߯�SC�RED����tpsc���_�hd�c�u�_y�ST���c�RACE_CF�G @��%����	F�
?���HNL 2A|�u���,� R��*�<�N�`��r������ITE�M 2B� ��%$123456�7890����  �=<���-�5�  #!;�C�O���� F���������C��� g�y�B��]��m� 	-GQ�u !GY�}�� )��/q/� ��=/�/��/�/%/ �/I/[/$?/??�/c? u?�/�?�/O?�?3?�? W?O)O;O�?GO�?�? �?aOO�O�O�OSO_ wO�O�O_7_�O�_�_ _�_+_=_oa_!o�_ EoWo�_mo�_�_�oo �o9o�o�o�o�o�o �o�oC�o���5 �Yk}��M�s� �������1���� g�'�9���E���ӏ�� �����۟�Q��u� ǟP���k�ϟ{����� ���;�M�_�ٯ��/� U�g�˯������� ��I�	���'ϣ��� ~�ٿ��������3���PW�i�2߾�S��C��>7��  ��7�� �ю߅�
 ����ߨ���f�UD�1:\����I�R_GRP 1D���� 	 @ ��=�O�9�o�]������������������:�%�?�   U�g�Q���u������� ��������)M;�q_����	����G�SCB ;2ES� @�= Oas������=�UTORIAL� FS���/B�V�_CONFIG GS��ы���w/'-�OUTPUT yHS�h ���/ �/�/�/�/?!?3?E? W?i?{?�?�?e!�/�? �?�?�?O!O3OEOWO iO{O�O�O�?�O�O�O �O__/_A_S_e_w_ �_�_�O�_�_�_�_o o+o=oOoaoso�o�o �o�_�o�o�o' 9K]o����o �����#�5�G� Y�k�}������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ�Q/ c%�/����)�;�M� _�q߃ߕߧ߹��߾� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������ /ASew��� �����+= Oas����� ��//'/9/K/]/ o/�/�/�/�/�/�/� �/?#?5?G?Y?k?}? �?�?�?�?�?�/�?O O1OCOUOgOyO�O�O �O�O�O�?�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�Ooo)o;oMo _oqo�o�o�o�o�o�o>������o �a�o9��]o�� �������#� 5��_Y�k�}������� ŏ׏�����1�C� T�g�y���������ӟ ���	��-�?�P�c� u���������ϯ�� ��)�;�L�_�q��� ������˿ݿ��� %�7�I�Z�m�ϑϣ� �����������!�3� E�V�i�{ߍߟ߱��� ��������/�A�R� e�w��������� ����+�=�O�`�s� �������������� '9K\�o�� ������#�5GV�$TX_�SCREEN 1}Iu�`�}�V�������Ev�4/F/ X/j/|/�///�/�/ �/�/??�/B?�/f? x?�?�?�?�?7?�?[? OO,O>OPObO�?�? �O�O�O�O�O�OiO_ �O:_L_^_p_�_�__ �_/_�_�_ oo$o6o �_�_lo~o�o�o�o�o =o�oao 2DV�h�o��$UAL�RM_MSG ?5v�� �Y
 ����%��I�<� N�l�r�����Ǐ���~�uSEV  �}���rECFG� Kv� � Y@�  A�M�   B�Y
 �`v������ ��ȟڟ����"�4��B�)�GRP 2L�3� 0Y	 �j����pI_BBL�_NOTE M�3�T���l`{b?���D_EFPRO�p%�{ (%ߏ�b �� -��Q�<�u�`��������Ͽ���޿ϕ�F�KEYDATA �1Nvv�p B�Y @�{ύ�`ʠjϴ��Ϡ�,("� ��Y��"�	�F�-�j� |�cߠ߇����߽��� ���0��T�;�x�� q�����������,�[΄�<�c�u��� ������`Q�����
 .@��dv�� ��M��* <N�r���� �[�//&/8/J/ �n/�/�/�/�/�/�/ i/�/?"?4?F?X?�/ |?�?�?�?�?�?e?�? OO0OBOTOfO�?�O �O�O�O�O�OsO__ ,_>_P_b_�O�_�_�_ �_�_�_�_�_o(o:o Lo^opoG��o�o�o�o �o�o�_$6HZ l~����� �� �2�D�V�h�z� 	�����ԏ���
� ��.�@�R�d�v���� ����П������*� <�N�`�r�����%��� ̯ޯ�����8�J� \�n�����!���ȿڿ ����"ϱ�F�X�j� |ώϠ�/��������� �߭�B�T�f�xߊ�h�߮߅d����`����������#�5��,!�f�� ��q���������� ��>�%�b�t�[��� ������������� :L3pW���o ��� $3�H Zl~���C� ��/ /2/�V/h/ z/�/�/�/?/�/�/�/ 
??.?@?�/d?v?�? �?�?�?M?�?�?OO *O<O�?`OrO�O�O�O �O�O[O�O__&_8_ J_�On_�_�_�_�_�_ W_�_�_o"o4oFoXo �_|o�o�o�o�o�oeo �o0BT�ox �������� �,�>�P�b�i���� ����Ώ��򏁏�(� :�L�^�p��������� ʟܟ�}��$�6�H� Z�l�~������Ưد ����� �2�D�V�h� z�	�����¿Կ��� 
ϙ�.�@�R�d�vψ� ϬϾ�������ߕ� *�<�N�`�r߄ߖ�%� �����������8� J�\�n���!����@�������"��p$����p����M�_�q�I������, ��������0 T;x�q��� ���,>%b I�m����� //�:/L/^/p/�/ �/��/�/�/�/ ?? $?�/H?Z?l?~?�?�? 1?�?�?�?�?O O�? DOVOhOzO�O�O�O?O �O�O�O
__._�OR_ d_v_�_�_�_;_�_�_ �_oo*o<o�_`oro �o�o�o�oIo�o�o &8�o\n�� ���W���"� 4�F��j�|������� ďS������0�B� T�+/x���������ҟ ُ����,�>�P�b� 񟆯������ί�o� ��(�:�L�^��� ������ʿܿ�}�� $�6�H�Z�l����Ϣ� ��������y�� �2� D�V�h�z�	ߞ߰��� �����߇��.�@�R� d�v��������� �����*�<�N�`�r� ������������� ��&8J\n���i���i���������,/F�jQ �������� //B/T/;/x/_/�/ �/�/�/�/�/�/?,? ?P?7?t?�?e��?�? �?�?�?O(O:OLO ^OpO�O�O#O�O�O�O �O __�O6_H_Z_l_ ~_�__�_�_�_�_�_ o o�_DoVohozo�o �o-o�o�o�o�o
 �o@Rdv��� ;�����*�� N�`�r�������7�̏ ޏ����&�8�Ǐ\� n���������E�ڟ� ���"�4�ßX�j�|� ������į�?���� �0�B�I�f�x����� ����ҿa�����,� >�P�߿tφϘϪϼ� ��]�����(�:�L� ^��ςߔߦ߸����� k� ��$�6�H�Z��� ~����������y� � �2�D�V�h���� ����������u�
 .@Rdv�� �����*< N`r�������/٠+�>٠���-/?/ Q-)/s/�/_&,q?�/ i?�/�/�/?�/4?? X?j?Q?�?u?�?�?�? �?�?OOOBO)OfO MO�O�O�O�O�O�O�O կ_,_>_P_b_t_� �_�_�_�_�_�_o�_ (o:oLo^opo�oo�o �o�o�o�o �o$6 HZl~��� �����2�D�V� h�z������ԏ� ��
����@�R�d�v� ����)���П���� ���<�N�`�r����� ��7�̯ޯ���&� ��J�\�n�������3� ȿڿ����"�4�_ X�j�|ώϠϲϹ��� ������0�B���f� xߊߜ߮���O����� ��,�>���b�t�� ������]����� (�:�L���p������� ����Y��� $6 HZ��~���� �g� 2DV �z������ u
//./@/R/d/� �/�/�/�/�/�/q/?�?*?<?N?`?r?I��t;�I�����?�?�=�?�?�?�6,�O&O�OJO1OnO�O gO�O�O�O�O�O�O�O "_4__X_?_|_�_u_ �_�_�_�_�_o�_0o oTofoEϊo�o�o�o �o�o�/,>P bt����� ���(�:�L�^�p� �������ʏ܏� � ��$�6�H�Z�l�~�� ����Ɵ؟����� � 2�D�V�h�z������ ¯ԯ���
���.�@� R�d�v��������п ����ϧ�<�N�`� rτϖ�%Ϻ������� �ߣ�8�J�\�n߀� �ߤ�{o��������� "�)�F�X�j�|��� ��A���������0� ��T�f�x�������=� ������,>�� bt����K� �(:�^p �����Y� / /$/6/H/�l/~/�/ �/�/�/U/�/�/? ? 2?D?V?�/z?�?�?�? �?�?c?�?
OO.O@O RO�?vO�O�O�O�O�O��O���K������__1]	_S_e_?V,Qo�_Io�_ �_�_�_�_o�_8oJo 1onoUo�o�o�o�o�o �o�o�o"	F-j |c������� ��0�B�T�cOx��� ������ҏ�s��� ,�>�P�b�񏆟���� ��Ο��o���(�:� L�^�p���������ʯ ܯ�}��$�6�H�Z� l���������ƿؿ� ���� �2�D�V�h�z� 	Ϟϰ��������χ� �.�@�R�d�v߈�� �߾���������*� <�N�`�r����� ���������8�J� \�n������������ ����"��FXj |��/���� �BTfx� ��=���// ,/�P/b/t/�/�/�/ 9/�/�/�/??(?:? �/^?p?�?�?�?�?G? �?�? OO$O6O�?ZO lO~O�O�O�O�OUO�O �O_ _2_D_�Oh_z_ �_�_�_�_Q_�_�_
o�o.o@oRo)�Tk}�)����}o@�o�myo�o�o�f,� �*N`G� k������� �8��\�n�U���y� ����ڏ�ӏ���4� F�%�j�|�������ğ �_�����0�B�T� �x���������үa� ����,�>�P�߯t� ��������ο�o�� �(�:�L�^��ϔ� �ϸ�����k� ��$� 6�H�Z�l��ϐߢߴ� ������y�� �2�D� V�h��ߌ������� ������.�@�R�d� v�������������� ��*<N`r� [������	 &8J\n��! �����/�4/ F/X/j/|/�//�/�/ �/�/�/??�/B?T? f?x?�?�?+?�?�?�? �?OO�?>OPObOtO �O�O�O9O�O�O�O_ _(_�OL_^_p_�_�_ �_5_�_�_�_ oo$o 6o�_Zolo~o�o�o�o Co�o�o�o 2�o Vhz����� ��{�� �������3�E��,1�v�)������� Џ���ۏ�*��N� 5�r���k�����̟ޟ ş��&��J�\�C� ��g������گ��� �"�4�CX�j�|��� ����ĿS������ 0�B�ѿf�xϊϜϮ� ��O�������,�>� P���t߆ߘߪ߼��� ]�����(�:�L��� p���������k�  ��$�6�H�Z���~� ����������g���  2DVh���� ����u
. @Rd����� ���˯/*/</N/ `/r/y�/�/�/�/�/ �/?�/&?8?J?\?n? �??�?�?�?�?�?�? �?"O4OFOXOjO|O�O O�O�O�O�O�O_�O 0_B_T_f_x_�__�_ �_�_�_�_oo�_>o Poboto�o�o'o�o�o �o�o�o:L^ p���5���  ��$��H�Z�l�~� ����1�Ə؏����� �2��$UI_I�NUSER  ����S�?�  3�7��_MENHIST� 1OS�  ( `����(/SOFT�PART/GEN�LINK?cur�rent=men�upage,153,1r����	���� ����936 ҟg�y�����,���Ư د���� ���D�V� h�z�����-�¿Կ� ��
�ϫ�@�R�d�v� �ϚϬ�;�������� �*߹�N�`�r߄ߖ��߸��Gѧ�G����� ��,�>�A�b�t�� ����K������� (�:�����p������� ����Y��� $6 H��l~���� Ug� 2DV �z������� ��
//./@/R/d/g �/�/�/�/�/�/q/? ?*?<?N?`?r??�? �?�?�?�?�??O&O 8OJO\OnO�?�O�O�O �O�O�O�O�O"_4_F_ X_j_|__�_�_�_�_ �_�_��0oBoTofo xo�o�_�o�o�o�o�o �o,>Pbt� �'������ �:�L�^�p�����#� ��ʏ܏� ��$��� H�Z�l�~�����1�Ɵ ؟���� �ooV� h�z���������ԯ� ��
��.���ϯd�v� ��������M����� �*�<�˿`�rτϖ� �Ϻ�I�[�����&� 8�J���n߀ߒߤ߶� ��W������"�4�F��1���$UI_P�ANEDATA �1Q���|��  	�}X����������� )���;���J�\� n�������������� ����"	F-j| c������4�� C�2�7 I[m���(� ���/!/3/E/� i/P/�/t/�/�/�/�/ �/???A?(?e?w?^?�?�6~���? �?OO&O8O�?\O� �O�O�O�O�O�OAO�O _�O4__X_j_Q_�_ u_�_�_�_�_�_o�_ 0oBo�?�?xo�o�o�o �o�o%o�oiO,> Pbt��o��� ����(��L�^� E���i�������܏Oo ao�$�6�H�Z�l��� ����Ɵ؟����  ���D�+�h�z�a��� ��¯ԯ����߯�.� �R�9�v�������� п�����k�<ϯ� `�rτϖϨϺ�!��� �������8�J�1�n� Uߒ�y߶��߯����� �"��X�j�|�� ������I����� 0�B�T�f����q��� ����������,> %bI���/� A��(:L� p�������  /g$//H/Z/A/~/ e/�/�/�/�/�/�/?��/2??V?��}��g?�?�?�?�?�?�?) �?O�OKO]OoO�O �O�OO�O�O�O�O�O #_
_G_._k_}_d_�_ �_�_�_�_�_�����$UI_POSTYPE  ��� 	 �o^o-bQUICKMEN  <k�Koao/`REST�ORE 1R��  �	�_��o�c�o�m,>Pbt �������� (�:�L��oY�k�}�� ��ʏ܏� ���$�6� H�Z�l�~�!�����Ɵ ؟ꟕ���	����V� h�z�����A�¯ԯ� ��
���.�@�R�d�v� !�+������˿��� �*�<�߿`�rτϖ� ��K��������߿� !�3�E߷πߒߤ߶� ��k������"�4�F���j�|����lgS�CRE|`?�m�u1sc�`�u2��3��4��5*��6��7��8����wTAT8m� �c<�%jUSER����2��T����ks���U4��5��6��7���8��-`NDO_CFG S<kw0v1�-`PD0�j��?Noneoba��_INFO 2Tj� �`0%�� /�^A��w �����$�HZ=~elOFFSET W<i�S��`[��� �/2/)/;/h/_/q/ �u/�/�/�/�/�/? .?%?7?I?�+�o�=�?��?
�?�?L���W�ORK X��?�?O+O�`�UFRAME  �5�����RTOL_A�BRT|O��BEN�B�O�HGRP 1�Y�i�aCz  A��C�A���O__�'_9_K_]_o[�F{`U��H��KMSK  ��5�KNyA%�	�%e?o�E_EVN�@�T��f��2Z�
 h���UEV�@!t�d:\event?_user\o``#C7eo�?U�F�=Y`�SP^acgspo�tweld�m!�C6�o�o�o���T! �_to2gw�Q V D��z���)� ���q����@�R� ��ݏ̏������I� 8�m��*���N�ǟٟ �������3�ޟ�5f�W@2[k��18.����� ��ί௻� ���:�L�'�p��� ]�������ܿ�ɿ� $���H�Z�5�kϐϢ���$VARS_C�ONFI��\� �FPS����CM�R�B2b��YU�	��B%1�: SC130E�F2 *.�2�S䙲�(��P�5U�V��?�P@PpsP�ȣ� OO�� ��L����������Z��mUA�U���U�h B���p�ht��ߕ��߹� ���������%��"� [���<���|�����z�X������IA DcM��,		d1DeF>TG�P �g �8~RTSYNC�� Di�HazWINURL ?�
Ђ����'SIONTwMOU o �?�=bdS۳�S�۵P�A F�R:\A\DAT�A  �� wMC�LOG�   UD1��EX�(�' ?B@ �����~�/�6/| �� n6  �������VO'��  =��͌!&�� ���TRAIN��T"�"rd�#p�%�(��4�d��eDk (���),= ��,?6?H?Z?l?�?�? �?�?�?�?�?�?O O�9_GEhfDk�`(��
�@(��B,\G�REkg�I�.��LEXgDh����1-e/VMPH?ASE  De��l��RTD_F�ILTER 2i.Dk �O��}�G_ Y_k_}_�_�_�_�_�_ �_�2_o)o;oMo_o�qo�o�o�o�o6SH�IFTMENU {1j;
 <),1%)/R���o T+=�as�� �����>��'��t�K�	LIVE�/SNA��%v�sfliv�N���+A � U����menu��ď^�#��5�A�ehk��hM�Ohl�N�z��Z%DT�m�O(�<� }@��$WAITDINENDL�h���OK  �؜Jr�S�ڙTIML��2�GğT�柀w��W�%�W�D�ؘRELE�A��d���G<Y��_ACT����t)ؘ_� n!	��%7�����;�RD�IS����$X�VR�Ao�N�$oZABC��1p��' ,� ��2��1���@�VSPT qq�M�!$
"��"�a��nτ�#�D/CSCH�@r!Eζ۲IP��s���� �2�D��MPC?F_G 1t�ɶa0������R�MP�iu���!p������߲�`  ��!$?���#!D�� D����H� ��	��-��Q�>��{����
�f���C4  ´!�3� �w� k�e�w�������_�q���#"6��$ٴe��@�v��8_CYLI�NDQwm� ��& ,(  * ��!#����� 0B�e ��p���� /J+/��a/H/�/@l/��/�/03xES� Ă�?(<K� Q?<?u?��?�?��喿1A��ZSPH�ERE 2yj� /�?o/�?1OOUO�/ �?�O�O/�O`OFO�O �O__tOQ_c_�O�O �__�_�_�_�_:_o�)o;oݰZZ%� � d�