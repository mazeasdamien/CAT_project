��   g�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����BIN_CF�G_TX 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG���DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST��NSS�* 8�D�FACE_NUM? �$DBG_LE�VEL�OM_N�AM� !� FTޒ @� LOsG_8	,CMO>�$DNLD_F�ILTER�SUBDIRCAPCp��8 . 4� �H{ADDRT�YP�H NGT1H����z +�LSq D $ROBOTIG ��PEER�� MwASK�MRU~;OMGDEV���PINFO� � $$$T�I K�RC�M+T A�$( /�QSIZ�!S� TATU�S_%$MAIL�SERV $P�LAN� <$L�IN<$CLU���<$TO�P7$CC�&FR�&Y�JEC|!Z%EN�B � ALAR:!B�TP,�#,�V8 S��$VA5R�)M�ON�&����&APPL�&PAp� �%��'POR��Y#_�!�"ALER�T�&i2URL �}Z3ATTAC���0ERR_THROU3US�9H!�8�� CH- c%�4MA�X?WS_|1���1MOD��1I��  �1o (�1PoWD  � LA��0�ND�1TRYFDELA-C�0G'AERSI��1Q'�ROBICLK_HM8 0Q'� XML+ 3_SGFRMU3T� f!OUU3 G_�-COP1�F33�AQ'qC[2�%�B_AU�� 9 R�!UPD�b&PCOU{!�CF�O 2 
$�V*W�@c%ACC�_HYQSNA�UM�MY1oW2?��RDM*  �$DIS��S=M	 l5��o!�"%Q7�IZP�%H� �VR�0�UP� �_DLVSPAR���QN,#
3 ��_�R!_WI�CT?Z_INDE�3^`gOFF� ~URmi�D�)c�  � t Z!`MO�N��cD��bHOUU#E%A�f�a�f�a��fLOCA� #{$NS0H_HE����@I�/  �d8`ARPH&�_7IPF�W_* O2�F``QFAsD90�VHO_� 5R42�PSWq?�TEL�� P��\�90WORAXQ�E� LV�[R2��ICE��p����$cs  ��)��q��
��
�p�PyS�A�w# kXK	�Iz0AL���' �
���F�����!�p�i��]$� 2Q��r ��������� Q���!�q����$� _?FLTR  �\�W �������!���$Q�2��7r{SH`D 1Q�E P㏙�f��� ş��韬��П1��� =��f���N���r�ӯ �������ޯ�Q�� u�8���\�������� ���ڿ;���_�"�X� �τϹ�|��Ϡ���� ���6�[���Bߣ� f��ߊ��߮���!��� E��i�,��P�b��� ��������/���(��e�T���L�����z _�LUA1�x!�1.��0��p���1|��p�255.0L��r��n���2�����d %7I[3 e��� ����[4���T'9[5U���{���[6���D �/�/)/s��Qȁ�a��a�P������ OQ� ��u.<�/ ?&?�/J?\?n?A?�?�?m�P�?�?�?�?�? O.O@OROOvO�O�O�u.kOl�q��O�L�
ZDT StatusZO�O5_G_Y_�n�}iRCon�nect: ir�c{T//alert^�_�_�_�_mW#_�oo,o>oPobot�2^�P~2g���go�o �o�o�o�o�o	-�?Qcul�$$c�962b37a-�1ac0-eb2�a-f1c7-8�c6eb5138?a8c  (�_�@_���"�p�1!
W��(��"S��JE�`� X��C� ��,$� ��W���ˏ���֏ ��%��I�0�m��f� ����ǟ�������!�4�u�R����� 7DM_�!�����SMTP_CTR�L 	����% ����DF���ۯt�ʯ ��'��Lz�N��!�
j��y�q�u�����Ԙ��#L�USTOM j�2�����  ���$_TCPIPd�j�a�H�%�"�EL������!���H!�T�b<�n�rj_3_tpd7� ��~i�!KCLG��L�i���5�!CR�T�ϔ����"u�!�CONS��M��[�ib_smon����