��  
��A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1RTU4QQ!Rx1R�� � $TIT91� ��� �Td��T0�ThP�T5�V6��V7�V8�V9�W0 �W�WOQ�U�WgQ�U�WU1�W1�W1�W1�W�2�R�SBN_CmF�!@$<!�J� ; ;2�1_CM�NT�$FLAsGS]�CHEK"{$�b_OPTJB� � ELLSETUP  `@�HO8@9 PR�1%x�c#�aREPR�hu0D+�@��b{u[HM9 MN�B;1^6 UTOBJ U��0 49DoEVIC�STI/@��� �@b3�4pBܢd�"VAL�#IS�P_UNI�tp_�DOcv7�yFR_F�@|%u13��A0s�C_WA�t,q�z�OFF_T@N�DEL�Lw0dq�1��Vr?^q�#S?�o`Q"U�t#*�Q3TB��bMO� �OE � [M������REV�B3IL���!XI� v��R  !D��`��$NOc`M�|����ɂ/#ǆ� ԅ��ނ��@Ded p �E RD_E��h��$FSSB6�`K�BD_SE�uAG*� G�2Q"_��2b�� V!�k5p`(��C��00q_ED� �� � t2�$!SL�p-D%$� �#r�B�ʀ_OK1��0] P_C� ʑ0tx��U �`LACI�!��a�Y�� �qCOsMM� # $D
�� ��@���J_\R BIGALLOW�G (Ku2-B�@�VAR���!�AB ����BL�@� �C ,K�q���`S�p��@M_O]˥���CCFS_UT��0 "�A�Cp'���+pXG��b�0 4�� IMCM ��#S@�p�9���i �_��"t����M�1� h$�IMPEE_F�s��s��� t����D_������D��F����_8����0 T@L��L�DI�s@G��� �P��$I�'��%�C�Fed X@GR�U@��Mb�NFL�I�\Ì@UIRE�i42� SWIT�n$`0_N�`S 2C�F�0M� �#u�D��!��v`�����`J�tV��[ E���.p�`�ʗELBOF� �շՀp`0���3����� F��2T��A`�rq1JY1��z _To!�Ҡp��g���G�� �r0WARNM �p#tC�v`�ç` � �COR-UrFL{TR��TRAT9 �T%p� $ACC�Vq��� ��r$OcRI�_&�RT��YS<���HG�0I�E��TW��A�I'��T�M�K��� �202�a1��HSDR�2��2�2J; �S���3��4��5���6��7��8��9�KD׀
 �2 @.� TRQ�$vf��4'�1�<�_U<�G��\�COec  <�� P�b�t�53>B_�L�LEC��!~�MULTI�4�"u�Q;2>�CHILD��;1t���@T� "'�STY92	r��=���)2�������ec# |r056$J ���`���uTOt���E^	EXTt�����2��22"(�0����$`@D	�`&��p%�����(p �"��`%�ak�����s�����&'�E�Au���Mw�9 �% ���TR�� ' �L@U#9 ���At�$JOB����P��}IG��( d p������^'#j��~�L�pOR�7) t$�FL�
RsNG%Q@�TBAΰ  �v&r�*`1t(��0 �x!�0�+P�p�%P"��*��͐U��qh�!�;2J�_R�Ҋ>�C<J�8&<J
 D`5CF9���x"�@?��P_p�7p7+ \@RO"pF̛0��IT�s�0NOM��>Ҹ4s�2�� @�U<PPgў�P8,"|Pn��0�P�9��� RA���l�?C��� �
$TͰtMD%3�0T��pU�`��΀+AHlr>�T1�JE�1\�J���PQ��p\Q��hQCYNT�P>��PDBGD̰�0-���PU6$$Po�|�u�AX����wTAI�sBUF,�8��A�1. ����F��`PI|�-@P�vWMuXM�Y�@�VF�vWSIMQSTO��q$KEE�SPA��  ?B�B>C�B^��P��/�`��MA�RG�u2�FAC<q�>�SLEW*1!@0����
�?�s�CW$c0'���pJB����qDECj�exxs�V%1 Ħ��CHNR�MPs�#$G_@�gD�_�@s���1_FP�5�@TC�fFӓC�Й���qC���+�VK�*��"*�J�Rx���SEGFRf$`IOh!�0STN�gLIN>�csPVZ��1_�A�D2����r� 2��hr�r�A��3` +^?���եq �`��q|`�����t��|aSIZ#�!�� �T�_@%�I��qRS�*s��2y{�Ip{�pTpLF�@�`��gCRC����CCTр��Ipڈ�a���b��MIN��a1순���D<iC �C/���!u`c�OP4�n j�EVj����F��_!uF��N@����|a��=h?KNL�A�C2�AVSCA�@A��r�@��4�  cSF0�$�;�Ir �4�@�05��	D-Oo %g��,,m����ޟ����RC�6� �n���sυ�U��Rޝ0HANC��$L�G��ɑDQ$t�NYDɖ��AR۰N��`aqg��ѫ�X�ME��0^�Y�[PS�RAg�X�CAZ�П���rEOB�FCT��A��`�2t!�Sh`0ADI��O ��y�s"y�n!����Ј��~#C�G3t!��BMPmt@�Y�3�af�AES$�����W_�;�BAS#XYZ'WPR��*�m!�Ɲ	]�R_L
 � 7K ���C�/�(z�J�LB�$�3�x���5�FORC���_AV;�MOM$*�)�SԫBP�H� 1�HB�ɀE�F���P�YLOAD&$EAR��t&3�2�Xrp��!�r��FD�� 8 T`I�Y3���E�&��Ct��MS�PU
$(kpD�&�7��b�9�B�	7EVI�
�!~e�X   $I��B@X��X<&�S]Y5� ��HOP�e�: �pALA�RML�2W�r}rR_�0; hb P�q�`M\qJ@$PL�`A��M����0�E@��	���V��0��qUU�PM3�U��<��TITu�
%��![q�BZ_;��3=� �B pQk��6NO_HEADE^a z��}ѯ��`􂳃����dF�ق�t�Pn��>��Ю@��uCIRT�R�`��ڈL��D�ClB@4�RJ����[Q��н�?�2>���O�R�r��OK��F`UgN_OO�Ҁ$�࠽��T��Ъ�I�V�aCnp�DBPXW�OY���@��$SqKADR��DBT�WTRL��Az�ր`fpbDs���6�DJj4 _�DQ5�AkPL�qwbWA��D^WcD�Ak�A=�|2CUMMY9�6�10�,3v �����B�[QPR��� 
�����C ��Y1$�a$^8�7�L�D�&�� ����0E���/e�PC�1F/U�_�PENEA@Tf��G=/���REC�OR"HH �@��C$L�#D$�PR���+jp��nq�_D$�qPROSS�
���
�r� -�$TRIG� �&P�AUS�#ltETU�RN�"�MR��U2� Ł� EW����?SIGNALA�QR�$LA�0O5�1E{$PD�F$Pİ"�AGc0�A�C~4�3��DO��D��"�!���&GO_AWAY��"MOZq�Z� D{CSG�CSCBg��I Իa#�<�ERIL0Nn�T�`$�������3�2L�@	BGAG~@R�P���44B0D�/ACD�OF�qF�� YF'C�CMA� X�'C�$FRCIN�I_�5#Ӑ@��$SNE�@�F�4L��>� J� ���<Ҡ���R/���P\ OVR10���$Ҡ�?$ESC_�`uDSBIOX��(T\e���VIB�� `s�zLZ��LV��pSS1W������VLP�:�Lk�ZX���ѣ�QPL���USC�P��A���A��MP1�U�C�PP��Rt`�S5QeU� ���Sg�Cg�Sd����dcC��g.���AUTO$�a҃oac�SB����T���C/B���2�f$VO�LT�g��A� ����1D���a��\�@��ORQҀr��$DH_TH�E� PRp� )t&wALPH&t��o�Jw� ! p���.�R�Ӏ{s�5c`r��A��ED��S\ F�!M�q�sV�r�v�ûvL�R�tk�:���BTHR�����T`����zV0ɖ���Q�DE7 ��1K�2P�C�X�C�f� F��#�g��QT,0� ��p���f�d����g����N~��s2>��Y0INHB��ILT� ɡ�T?��3��/� ఩3�P)Q0Q�T)Pe�Z�0Y�AF5�OM� r�o��z���o�)Pڳ�|���o�P��͘o�P�L?�x��o�TMOUXc|��o�� w�+� �1�H��A��g�1Io�����DI~����'�STI�󍣣�O`��� Hҽ�ANǥ��Q�S8��b͑�h!$kЪ���/�_Ig�&yPRAOP�P.C��kӦMCNQe�E�=L�VERSe��bP'PI/�F{�������G�DN��G����o�F�2��ӷo��MԺ�F��_ԴM�D��䧭�ed��3�ea���DO� ��U��2�j�ʹDI��e�۴���번������/�F00�����ON����܅QI�VALȤCR�_SIZJ���A&�REQ�R���2���D�CH)���ʹ���z�D��ō��&�S�_�>X��/WFLG����/U$CV�iM�@VQ��FLX���"�B��-䯤��A�LJP�C��� �bT^�W^� gRxc� cQ�NDMS�mљK�C{P_M�  �S�TW.������h�AL�PY�YQk����V��e�IAG�'�d(7���T�A�P� R��A^��]� `]�d	`]�6[�q_D�� g��c����YP����r��"8Tc� ? �����1��T�ۡ���LH�?��! �0��LDĀ��U0nJFRI�0 �P`��I\15�jIV10U�s1IUP�PZ�0�Q��C�LW���
�PL�C��S��CWC�	/�� �IZ! Fů�T�Q�g��?���g��~�
�P�5RSMI�T��0�  b *�sd2AMWda_T
p5��0?NS_PEA��;�8���ܢSAV������7%I��CAR�؀�P�!<$f�E"CR �����T[#El@I�N\"STD;�[!F�`'�x'QOF7�k%Bf�"RCO҇&RC�� v(���1�R�'=�G%��WMA�Q_naI��A�Q���a$2F�-4I�*7I>R99/Q97��Rk8M�H!C�`Rp � tp�2F��S#DNX�Va�� �5�@�2�AK P $M!��s�S�17��3nc@%j9f��4[�RA�D��0CY_ L L!IG10'1BV�h1@�07H2�NOàx���CDEVIP� M�0$�RBT�FSPc3�C-T�DBY4�A�G3�3�HNDGD�1N ]H�0GRP�HE�!XL<Uj�SDF02�:�4L�` O�Bp���U�FBQ\�FEN�@�uSV��3 �17P d�@DO���PMCS�?P��?P|uRN�HOTSW24:�DpELE�1�U80\�P�RQ T�@I�`[r@  f�o`OL�GCHA8F#��c:�4���3�A�0R � �$MDLb 2Q��EXȃqn6�q� P�i�c�e�cJ]�	�e����#�n�d�g]PTO�a�� tb1U�4SL�AV� S  n�INP���F��By��1_��ENU�1T; $
�PC_eq�2� �RLvw�0�2bpS{HO�� U ���A�a�q�2rr�v�u��vu^rCF\ ?V` ,�xr�OG�W�p�%�q ��Yp�rI��!�M�AX��q0 AY�vW�A (�NTV���rV�E�0�uSKIg�T��`�}�2S���JsX!��C��s��f���_SV��`XCL�UL� �p�ONLdB�߃Y�T��OT�U�HI_V�!��AP7PLY��HI�P�v��_ML�� $VRFY�����=M3IOC_�Z�" 1��l���O�@��LS/"@$DUMMY4x𛐒�_C= L_TPJ�T�8#Cc�1CNF�Օ@_E��j@�1���D#�Q_������PCP�B���R S��k�����u �� W ���� RT_�@`�[uNOC�R X;r��TEL������rzDG��x`Y D���P_BA`L#c��!�ȥ_Ѐ�ҬHУ6Tb�E�� �Znp�R�SAR�GI�!$���`Y�n�SGN�1[ �8�`ЎIGNQ�G�,J����VJ�d�>[�ANNUN��ޕ���_E�'wATCH������Ķ���u\ <�0�@����S$ah�����������1EF I�� �] @�0F��I}T�	$TOT! @�C�����-�M�@NIva^,B�����A�q��DAY�3LOAD�D�&������ �EFV��XI@R_\���I�O���a �AD�J_R_!x``���� 2�"�������`_��PI�cѝD�u�AG����1a �0��\�=� \��䇡��U! ���CTsRLN p b;��TRA��#IDLE_PW��G�XԮQ���V�GV_WЉ`a� �'��Ax`c�� 1$k��P�STAC�#M��Q���R2 A�e����SW��A�����Չ``f�OHα(OPP��#IR9O� �"BRK�Ө#AB��o�㾢��@�  ��F�Չ`b��x�"@�RQDW��MS��6X�'2�?IFECALƳ� 10tND��M���`B��� 5f��CP¢ʱN� Y���FL�A#��OV Y�H�EO��"SUPPOd���gL�p��Q�R�"Xт��Y��Z��W�����P����Bт�XZbq�$Y2@C	O@P�S��2
報��bD!���"g�1I��0�sd `�@CACH�5�VcS���+0LA SUFFI���p7�Yq����6��*�MS�W�e 8vKE�YIMAG�TM@S��&�""@r�2>|�OCVIEN�6�wf ^aBGL[��F��?� 	�����0�g���PST��!�b������������EMA�I�`N��Az@�FAU� 7�h^�Yq��Z�U�3��- E�5�i< $d#�USWи�ITߓ�BUF����DN���H�SUB-$�DC����"��p"SAV x%:"#�_q�X��'�r��P$�UORDO��P_- ^%=��(OT�T��_�P���0LM0$��$g��'AX�3.�bU�X- ���#_GD�
�pYN_��7�jT�D�E��M��U��T��FQ�av��DIBEDT�0ICh�6�k;r�GN!"�&E�$`���QvP���FP l (�pSV� �Tć�[����1��m� �<�n���#C_RYIKQ�#B\� D3p�RE��1DSPd6BP�`hIIMx# ]C�A��1A�U:G��48!CM�IP\�C��~ \DTH^ oSPB2��T\�]CHS�3?CGBSCi�m ��V�d�VP�#T_D*cCONVˁG*cT^ $ZF- FD�A�d?C�0�"1R�SC��DeCM�ER�T�1FBCM�P�S�0ET�S mnFU��DU! b���6ђCDSI��@� �@O���o�G�QR�Q�U=��MS��Z-��P�T�{��Q[�A�1p�� "��Q�4$Z!O�0+�q�$�U��ޔ2�ePM��eCN�$�x�l�l�iGROU�Wd����S� �MN�k u�eu�ep
||�i��cH�p!�ez��0CYC��shw�c��:6�zDE�_D���RO�aP��qf��gv3�O���vO��w�tU���B�u��8��&p�ALA �1q��1z�Г0�PB�ᣠ���ER�T7��Rr �,�0>��%>�G1L~R1q 
MAo�w�Ց�1s�����Ų�R��Pv���C�����U�A��2��0V`t/H *��L�� �	��V°��12�b� 2���2���2���2��*2�7/�8/�9/�D�T1�;�1H�1U�1b�U1o�1|�1��1���1��2��2;�H�2�U�2b�2o�2|�2���2��2��3��3R;�3H�U�3b�3o�U3|�3��3��3���4���2XT�ѡ1u ��\0xf\0�Ug0}��@e��FDR��7vT VE���!�G�RG�RE��F�G�SOVM6C�A��TROV�DTl� 
�MX�IN�8��	���IND(�*�!
Tȑ0E0Z0G-1����PM�3�D��R�IV�Pq�SGEA-R6AIO*�KڲQN�0��1�(��P�0�a>SZ_MCM8 G� �F��UR�Rwx���P!? ���]p?&�C�?&�E
�.�L:!�P���xL��Pq��R�I�;�:#ETUP?2_ y b�9##TD�@
�7%T�`>�p�׎��r�BACQ2Gz T�:"�4)�:�%�PBW�(�IFIf�W M������PTP��FLUI�{ иqd UR��!��B�1P�0 �sEMP�pC2$�b�S�?xn�J8��� �#VRT^��0_x$SHOc�L)��ASSP�!s��@��BG_;�������U���b���o�FORaC�q�!�Qd|�KFU�1�2�2�3q�^ (�} |d�7NAV_a�b�����ְS�q�$VgISI��ۂSC4CSELЮ�� �rV�pOg�$b�ְ�b��$r�I���@��FMR2��~ ���P{r���0 ���������������ڲ_U���LIM�IT_���TC_L�MƤ϶�DGCL�F_Å�DY�LD�>т�5��yϋķ�Mԝ��SJ-	 �T�FS� �T� �Pl�	�3E0$E#X_	 	1!0YP�ba	3B5B�G�'Q��� �d��RS�Wa%ONZP�EBcUG��ߵGR�`�g@U{SBK�aO1n� C�PO ����P��Mt�O,t`SMu�E�"
��F�y`_E � ��0�pm� �T�ERM%�%IaO�RI�1 �%o�S%MpOs� �4&� �S`Z(�f)UP�p ?�� -E�yb��b�)#� �x�G<�*� ELTO7�p�0BPFI*c�1Ѝ�a�@$�$�$UFR��$���!0�U&H OT7BPT�a���#3NST�pPATz�q74PTHJ�a��PE�P�3ap�!AR�Ti �%� i 12�"R�EL{:�1SHFTP�B�!?1m8_��R�P��SX& c $r'�0�@h����]s\1�0I�0�eU�R �pPAY�LO�@nqDYN_�#�O��R?14�Ʌ�@ERV:�
AX�8^�7��p{2ס�eE��R�CN�ɅASYMFgLTRɅ�!WJ�'^�Z�E^�i1�IX��QU�D�pAm5� YF�5aPFP$CFQ�6OR�p�M��i!������>0� Eas�Hs��T� �%2X���POC�!�>��$OP����rc��ֱ��jbRE�PR�#\1��q?3eH�R=5�U�X�1>��e$PWR���u�=@R_�Sb4d�t6�#UD^��VR�"w ���$H�ս!L`ADDRxfHB!GA2eaZaSaTo��R��� Hl�SSC�ף�e壒eU���eb�SE���$ H�SCD��� $N�zP_�p_��2�b�PE�D�<!HTT�P_��H�� (���OBJ�pSb��$^fLE03UPqt� � n�Q�p�%_U�T�arSKP���2�KR�gHIT ����zP��Par��^�0��P�PSS�����JQUERY_F�LA�!_qB_WE�BSOC���HW����!���`�@IONCPUVd�O � vq:�7��d8��d8�b����IHMI_E�D] T �7RHv��?$d�FAV@ ��}��IOLN.�ґ 8l�R���0�$SL!R$I�NPUT_��$t�P��P�� ��wSLAz �������|C��|B������`F_AS����$L��5w�ѿ1��b�!;ࢃ���@HY|�l�E�SQ �wUOP�� `1� ��^f8�\�8�c����PP�3�P��Αc�ےĖ>8aIP_ME��m�7� X1�IPZ`V�_NETV�pd��R|�+��qWDSaP��p���BGV�}`g�MgAm�� lL(�3TA"B<pA�TIԕ�E�� ���0�PS��BU ID �r����P���ad�L��10��v���Ċ���N	� 
��I�RCA̰!� �k �Sy�CY�`EAT�K�}�P�8��3�h�]�RY0�A���AD�AY_w���NTVA7�Ԡ��܂]5����gSCA@��CL�� w�,�Ţz�m����X^2�'�N_�PC�)�Ţ��n����C� \�0rw����`���? 2� b�e����m���ғ�0r��L�AB11�� ��UN�I
���C ITY���e�^e��R����|��?�R_URLF�o�$AL��EN��`�e�t �sTh�T_}U]�ABKY_2���2DIS�����1��J�m���$`ҙE��R����O �A�灋�Jh��F�L+]������Ѭ
��UJR��� �;�F3�7��'��Q����J7��O�B$J8�7`��
���7����83� �AP�HI� Q�P�D�J7J8�2i�L�_KE��  ��KZ�LM� 7� <�XR$�-��C�WATCH_V�A��'@��,vFIE�L�Pcy$ ����� D '1V0@@���C�T���%�)�LG~ ��� $=�?LG_SIZ[t�`2�� 1�(�1�FD<�I0�G��>�/� I� ;�.�S7��� ��(� ��^�� ���A�� _CM32
�
F�A..��T(-��29�S�  S(�S^�_IRi��S k].�RS��N0  MZIP3DU~���LN��r����p2�OԐ��c�KPL�DAU!EA�`Z�nT�7-GHoR��4�B�OO�a�� CK��IT�sk^`�G�REk��SCRX; �sL�DIF�S� n�`RGI"$D�@̆?��T��t4�SAs�3�W�4�?�JG=M'MNCH�s4�FN{�&K?'-�=)�UFK(�0K(FWDvK(HL�)STPK*�VK(��K(rK(RS"�)HPg+<�CT�# �B?��`�9U�a_$@�� %��T�R"G/)�0POV7�*��#�5$W�M)EX;�TUI=%I��B�G���Ar��3#�3; ��$S�ű�	ᰟ�0�NO�6ANA4�{Q²�AI4�Zt�EDCAS���cQC�cQBOWHEOcGS=ӁBnHSzH�IGNG�ŰY�<!��k�ZDDEV�'L�Lu� Y�eФ4���TU$=���P(�A����#Al������P��3��sPOS1IU2IU3IQ��2R@eЦ �S{FP,D��������a�uq0X��VST��R8�Y$��0�P �$E�VC�[ep�`�Vpf`��4dѧ L
� Z���o�0��SxpO��t��`idEp��_ �
pW�q޳��c� �MC�� =���CLDP��s�TRQLI��u��i�dFL\��b���c�1D���g�LD�e�d�eORG{��! r��?RESERV;�Lt�G�LtR��c��� � 	�e�%�d�e&��PT�`��	0q�t}�vRCLMC�t@L^�y]��q��MI��#������$DE?BUGMAS]��������U�T7@��Et���`FRQ���� � "�H_RS_RU�aa�^�Al�#5FREQ�8 t$�00�OV�ER��Y�&��V��PnT!EFI̠%Fa�_���X�yt� q\
Ќ��$U�P�\�?�pűPSHP��	��C@�s�����sU�$�?(� 	���MISC��ծ d��QRQ���	I�TB�̠ 1���1��AXsҀ�|����EXCES"Ҥ\�c�Mj�����t�s�L�b�SC�P O� HY���_���~��������M�K Ա���%�B�_�FLICAdB��QUIRE�#M�Os�O���iPML:c`M�Ų �`z����a��r�aND�����Q�#����DO�INAUT�O�RSM����@�N�r��3�rp�PwSTL�� 4�7LOC�VRI���U;EX��ANG-B-�n
�ODA\��p�1���Ю�MF�e� ���Ybb�0le�� #�gSUPufV�FX���IGG~ � ��pbc��E�bc	6bd ��݂�R4��PD��PS�`4�s3/�W�TI���<p���M~��� �t��MD��IA) ��W@���q��H�����DIA8��Ñ�W����/Q�1��D?)�`�O�Ӧ��� �CUG�VОp-��ՑO�_�=ѹ ���ДS������i�{�P{�� ���P�z�KE2��H-$qB: n֤�ND2�r�����2_TXkdX�TRAWC���r�M8Ԁ4q�`�P.�}X0���P�d�SB)`�U/SWCS;�Tf����V�PULS����N�S��n�
u�JOIN�� u�6`"��r=b��cb���P�r�����cb��o�TA�8�{����� �E&r�SC��PJ��
��R�PL	� �&��LO9>л�m�&� l���Bҍ�܅�Z�RR2g��� 1}�A�q� d$G�I���G�EA��2���p �EPRINE��<;$R��SW0�t��sABCŸD_Jp��z�-���_J3D
>1SP���-�	P>e3dG�8`-���J�s�mr�qO��AI��M�CSKP �j�3�3��J@L��Q�����_cAZ�r�6EL�A<��qOCMP��M�����RTD�a�11���m��P1���0:�Z�SMG� ��v�tJG�`SCLɐ���SPH_�@L����-���RTEaR ����A_D@
�!ڰA�@�SL�$sDIL�23U�kDF��5!LW;(7VEL�aINwb�0^ _BLW@-�f$�� �qV$k'�'|%�s� �ECHR�tTSAY_�����E5`B���B��%�B-���!:5`_S� ��%�"%`��$��9,&Ր�DHɐ��=��8P�$V�����1$��������$�A�Q�R5�>��H �$BEL.�m��_ACCEl!�7<�q�0IRC_ ���?pNT��S$PSɐ�bL����5 �c���63�F@�6�ѩ9�G�3G3�2S�̑_�FQs2P@VA��7��1_MG|�DDsA"��FW�`Q�3�E�3�2��HDE�KPPAByN�7�SPEEfB JQ�O�`�JQ���1>�!$USE_G��P]P#�CTRTY�@��0�q �YNf�A =V� ��=QM9�M��o�m@OX AjTINC'Ԓ��B�D���W����ENCF��-��1x�2���0INPO	�aI�2�U���NTV#>}%NT23_9"���cLOJ ��`��I נ�!f? �#��g`�U"�C� �VMOS�IxA;�Z�VA��L�P?ERCH  >c��� �g���ck�$b�t�k�\T'U-@U@�A�2�eLT�6���Up�$jv:fTRK�сAY���c�Oq�2�^uSs��g��R�McOM)ҍ��MP���C��jsACR���DU��KBS_BC?KLSH_C�2�u 9�_f��ES,� ��R
�|TQ�CLALM�Tpl�p%0<�CHK� |����GLRTYo�����T���Q��Td_UM���C���A�ܧ��@LMTa _L q0O����ˇEō� ؋Ā�5��8v �qYQ��`'��hPC�a�hHp���wE��CMC��\�@�GCN_��N��L���SF�1�iV'R����W�[��2ʕ_�CAT��SH���D �V��q�V~��1~��f��PA���R_P��ys_� �Vv���fs,x�i�JGŰT�v���y�z�TORQU`PgRcoy�@OUW�0jb{�@ݢ_W�uOt��t1��e3��k3��I*�I�Ik3F���P��}@VC�00
Q�tp�1w�u@��v���JRKw�����p�DB�Ms�pMC�? DLe1�bGRV����e3��k3ܱH_p��ڳ"@)�COS6�i6�LN��Y�z�`� e0[ɮ[�-��ʅ�K�b׵ZT�jfܱMYb����B���J���THE{T0*eNK23k3� �_3c�CB%�CB_3C��AS{ I�-�0X�e3X�%�SBe3v�N0�GTS��ACz�R��A���ڔ�$DUf�w����m%��
|%Q�a_;��Q��0�3�Kv�s(R��A��A�J�(�3�3�LP!H6���U�Sz��� �Œ���Ƽ���ƊR�Vc�VX�U0{�V���V��V��V��V*��V��V��Hc�|栂�z�������H��H���H��H��H��OJT�Oc�O	y�O��UO��O��O��O��O��O��F�Eѡ	��ŦV�SPBAL�ANCE_���LmE��H_�SP�!�v�������PFULC�$$���*{1�uUTO_a��i�T1T2e�22NH��2�P���q&P��2�3�qTpO. |�1�INSEG�2�CaREV�C`�QD3IF9u91��,"1�B�OB�,��¶w2Ǡ�PS��LC�HWAR�B�2ABH��u�#C`��\Q�%
��X\qP
�{&:�F2Z� 
|"ڡ�1�U7ROB��CR�b�%�p� �C�1_�d�T � x $WEIGHYPF�P$T��#{�IYQ�`IFQ�@LAG�JR)�SJR�JRBI�L05OD�pF`2S�T�02P�,�0P�0��!� �� 
�Px�2KQ�1  2�Qd^6DEBU3L@z_2��MMY9�5��N2��4�P$D�A�a$�0v�� ��DO_:�0A�!� <� y6�o%�KQ7�BI2A0N��SH_(`KPf2O�9� �� %"��T�P�Q��T��4��0TICK 34 TE1�0%qC�pz@N��TC��R�pKQD"�E�D"�E�0PROMP�YSE6� $I�R��IQo��B�`RMCAIᰄQ[R�E_*0C�C�eq]PR�7COD~3FUQP6ID_�.U��B� �G_SUFF-� �$3@Q�A�BD�O�G��EC0�FGR *3D"lT�CxTD"�UD"��U��lT�4�0�� Hn _FI}19�S7ORDI1 � �2�36��RIQ�0$�ZDT5U�!g0�5��4 *�L_N�A%Az@<b�EDEF_ILh<b�FXd�EP2��FZ4�F�c�E�e�FISྐAp�D�c�CVdё�44��!�Z2�DX�rt~3D��O|� BLOCKE2��fS�O�O�G�alRfPUMkU<blT�clT�elT �bxRnswUgcxT�dxR X6�v�a�SO e��U<b��U�c�S�w�hX?@P@ �dO@�a��0WMx�L�Cs���T�E7��4�( >$1LOMB_f����02VIS��IT�Y2Av�OJ3A_�FRIU�� SI�a��	Rw@҇�@҇)3�32W��W���䰆��_��QEAS 3�R�����p�Bӆ�4Љ5Љ63OR�MULA_I2��E�THR2 �G�,g�� Ч<8�5C?OEFF_O^A�HԔ^A��G
�3S0F�2CA&�?�3$H��3k�g0GR� ?� � $Cp�BXN@TM6wN�Cu�dBKsh�CER�T�,t+d�P�  NL�L�TpS6�_SV t����p��P�� ����P� @�SETU�cMEA�@KPi��0f1�R� � �  ��  �0��'� $�'�q2�Abz@q7qt����Rb��Ap�apn��� �PREC�Q,��d1SK_� 4��� P�!1_USER�"��3 �����VELe���3 �ܵrD!I`��MT?A�CFG���  �|@�Oj"NORaE� $@'��SI�!1��w6M"UX�P��A�DE�� _$KEY_�3��$JOGu��S�V����Ñ!Y�5�SAWj"�aaӍ�T4��GIY:�4 �� 4  �e'2k!XYZ�S���3k ����_ERR���! � ��=AP����1��{�$BUF�f�XX�  �MO�R4�� H� CU �$Ak!j��Aa�����Q$� ���aW�� ���G6�� � $SI���Y�İVOY���O�BJEZ�ADJyU�2\�ELAY`�4�%��D
�OU�P�Ÿj�JQ�R=i�T�9��8��2DIR�=�E����� DY�N��"��TY�"R�O@I0�"�OPWwORK���,�0�SYSBU1�Y�SCOP��?Җ���U��b�PCp���PAð�,���f"Y�OP�PU�!��!M�$�IMAG/�� 1�Z23IMz�M�IN��~J�RGOVRDv���İ'�P)�I� ��P�s��k"LApB�|��'�PMC_E`?ѭ1N1 M��1�211�2�v�SL���� � $OV�SL��c��a�`c�2j"��_v�#�Pw��#�P-B=�2bC�� >`��q?w�_Z�ER7���Z�$�Gd�� ������� �@����%O6PRI\�� 
�P�	���9�PL���  �$FREE�E���9����L����e�Tg ^0ATUS>��TRC_Ta�N�MBR�W@+��c�18,`��� D�1%�fÌ�L���"���QJ ����XEQ3���Ą��� � PUPa��`�aPX�@w"�43�����PG��ڻ�$SUB�?�%�q?�JMP�WAIT�2W%L�O��FeA�RCV!F�A}@R"Z!RV�.R"ACCt R��pB��'IGNR_PL^�DBTB^0P�aFS!BWP�$/�U1@��%IG�@I��T'NLN�&�"R��<r��N�@��PEED|�HADOW^0��/���EK4")!�W`SPD0!� L�<A2�X`k0��y3UCNI*�{w0�R��|LY`� I��P�H_PK����RETRIE�3�)����0�@FI���� ��P�0�4 2}��DBGLV�#?LOGSIZ]��aKKTw!U��0DD�#�� _T���M��C��R�V@?MRPC5���CHECK� X�( ��0!�#��9a�L\#Y�NPA*pT�2����@P1 � h $AR#B !R��S�a��O�P����ATT���"��#F`V@2��aS�3UX���B��PLI�"0!�� $���ITCH�R"�W��AS�ܿ2RRLLB0!��� $BA��DsY�BAM� f�Y��PJ5u�	��R�6�VzQ_KNOWh�C�Rv�Ud�AD�X��v0DðiPAYGLOA,��p#c_O�(,g��,gZ)cL�q���L_�� !@�eb�Q��rd���fF�iC��`j+�cd���I`hR��`g;�|dBd>���JQ��a_Jja:۱��AND:�|�`tjb~a9�*�PL� ?AL_ �^Pv0P���Q��Ce�D(c�Ed��J3p1v�{ T�@PDCK���>����_ALPHAs�sBE��z�AS|� ���!�� �s ��"oD_1)j52SdD�AR����u� ���TIA4�/�5/�6e�MOM�|�;�[�H�[�U��Bn AD;��H��U�PUB��R`���H����U��Q�1p��1 �pف2a� �B�RQ���� e$PI��1�s̱.g$��kHi$�I0�I>�I�L��}�!}�!���}rr�b��/3HIGmS/3o%h4Ɩh4o% � V�Ɩ��՘�!䙥!o%SAMP�o�8��Ɨ9�o%�Ps  ��h��� ��w� �� h0�p�� ������8�ȿ�-pU�H 0��IN Ǭ-p�Ψ�Ťo"Ъ����0�GAMMb��SSԨ ET��dK���D�t��
$4p�IBR�2I�$HI��_f�O������E�в�A��ϰ��LW����Ϲ����r誖0jqC�%CHK����  v~I_�����,r�x,q���z�s����y�1s ��$cx 1����I� RCH_D�!� RN3��#��LEUࡒ���x��}�0MSWFL�$�ہSCR(100;�,@v�37B[֝��`�;���o�h0~�PI3}A�METHOBX���%��AX �qX20��2ERI��J8�3d�R�0�e	�"�pFU�9�}�⌣��&�L��9�;�O�OP}���Qጡ��APP�3F��@U�v�a岣RT��0�O ph0.ŧ��턱 1�#��k ��L����RA�@MG$����SV��P΢CURA��GRyO50��S_SA�QX��3��NO�pC� ��t3����4oFoR������x��R���� �DOg1A��bAw�qڪ� ���Aϗ�A��1-���ic'�QM�� 7� �YL"��a
����S�b4�7B�@I��0��ď�a_��9CѣM_Wb��!A���=�M� ��`�0q|$J�R1I��"�PM$��� ��A{ ��WC�$��L1QVaC�tA��tA�tAUt� ͰN��P��dS��-pX�0O��s,qZ��Py ��+ ���M��x�u� ��������2������5uL�q_XR� |tq �3�[��&H��&U�3� 4��'�&N�sQ}��0���q"
��0W`q$P��A�PMON_Q}U=� � 8�@�QCOU���@QT�H]�HO|80HY�SPES�R80UE�#0)��@OVT�  ��0P!��T�RUNW_TO�OPO��N�� P`�5C��|A�INDE��R�OGRA� HP� 2>A�NE_NO�4�5�IT��0e0INFO�1� `Q�:�1ڎ�1OI�2� =(��SLEQ�� A諕 @�6	e0S_EwDIT�1� �PR�Kށ����E��sNUpGjHAUTO�mECOPYށ���L��[�M��N�@�KKƯPRUT� �BNuF�0UlR$G�2|�D=RGADJ�1�� htpX_� I����#V�#VW!XP@!X�#VϓP��Np�_CYCoSN�S_h3�q 	�L�GOXã�NYQ_/FREQÂW֠:�N�QSIZB��L^`�r�P!QV�֠��CR1E����Y�IF>��3�NAA�%�T_G>��STATUt ��w7MAIL?��q=a<�34LAST=a�qކTELEM�Q� ��qNABot�EASI|a1l�� XЀkb��<�f�ҳ���I �0�īR��;1� ��b�ABS1SpE�0ӐV_a�fBAS]r�e���āU񐳐H�$,qwRM�R�c�� ��:s�𐠲Xat����R��| 	�b 2� ���� �v(r�w]r ���(r8�w� �DOU�3��^p��$$CX`S0��� ���c�fc� �pY�SI9����XK�IRTU�����A� _WRK 2� @� �0  �5��w���t��� ��	ɀ��ݏc�A�!�ˏ�����,��8�ȁ>�s�����Q�B�SSA� 1"��? <a�ҟ �����,�>�P�b� t���������ί�� ��(�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢ� ����������� �2� D�V�h�zߌߞ߰�������ߝ�CC�@XL�MT0�����  d��IN����]P�`EXE'�S��6�^0-r ��@�Q�D�V��Svp@�S��%select?_macro�߫�����IOCNV��c	� ��P��U�p(㲗��0V 1]^�P $N���0H�B�E�A�?���j  h�z������������� ��
.@Rdv ������� *<N`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6 HZl~���� ���� �2�D�V� h�z�������ԏ� ��
��.�@�R�d�v� ��������П������*�<�N���LAR�MRECOV ����6�!�LMD/G 1�<������_IF �1��d  RVO�-003 Dea�dman swi�tch r��as�ed 	�TCP)� d out t�ion for BWD��7�?��S��e�w�������, �
 ��ҿM�>I�PL_FANUC�_SMPLG> � LINE 0 ��T2  ABO�RTED��JO�INT 100 �%׿:�!�$�R�P_CLO�@���k�E�SBN-0�60 Inval�id attri�bute syn�tax data����������NGT�OL  j� 	? A   1�C����PPINFO �� ��v߈�8�߬��  ���� �ߕ������)��%�_�I��m���O��������	��-�?� Q�c�u�����������PPLICATI�ON ?������L�R Handli�ngTool� �
V9.40P�/17B���
8g834�F0F3170	�K'7DF5 ����None��F{RA�� 6c~��_ACTIVi��]�  ��*�  ~�UTOMODi����(��CHGAoPONL +oOUPL��1	ة� hl~���CUREQ 1
�ث  T���	����$��� ��//'/9/�/]/ޖ��� �$H�k�*HTTHKY�/
���$\~/�/>?? r/,?J?P?b?t?�?�? �?�?�?�?:OOO(O FOLO^OpO�O�O�O�O �O�O6_ __$_B_H_ Z_l_~_�_�_�_�_�_ 2o�_o o>oDoVoho zo�o�o�o�o�o.�o 
:@Rdv� ����*���� 6�<�N�`�r������� ��̏&�����2�8� J�\�n���������ȟ "�����.�4�F�X� j�|�������į�� ���*�0�B�T�f�x�����������俬T�O���DO_CLEAN8�o��NM   � ���������ߠDSPDRYRv�&�HI��@��q� �ߕߧ߹����������%�7�I��MAX@��V���Gg�XV��fcf�PLUG�GVW�cPRC*(�B����`�R����O��1�C�SEGF/K��*�ϩπq�����������$�LAPN�a��#1 CUgy�������*TOTAL����KUSENU
N�[ <�@鲬�RGDISPMM�C-�!1C5�y�@I@C�[OL�n�9��W_STRING� 1'
�kM S�

��_ITEM1�  n���//*/ </N/`/r/�/�/�/�/��/�/�/??&?8?�I/O SIG�NAL�
�������Ӱ�����޼�ƭ��خ��ޮ�����5��9�����ײ�޿ = 100������������۸���3 ��1�2t3�5��3ʰ��ް�� t�MH ��װ��A����??=??OQOcOuO�O �O�O�O�O�R�� R���O,_>_P_b_t_ �_�_�_�_�_�_�_o�o(o:oLo^opo�OWOR-���a_�o�o �o�o*<N` r�������8��&�PO�e	L��k5�o������� ��ɏۏ����#�5� G�Y�k�}�������şG�DEVO��c�ݟ �)�;�M�_�q����� ����˯ݯ���%��7�I�[�m�PALT]���on���ο� ���(�:�L�^�p� �ϔϦϸ������� ���GRIl��8Ѭ� �`�r߄ߖߨߺ��� ������&�8�J�\�@n����&�R] ��P߶���(�:�L� ^�p���������������� $6H��PREG��� ��Z� ����&8 J\n��������N=�$ARG�_�`D ?	����/!�  	$N6W	[C(]C'�N7�d)" SBN_CO�NFIG�0/+�1�2�!|!CII_SAVE  N4��!�#" TCELL�SETUP �/*%  OME_�ION=N<%MO�V_H� �/?RE�P��M?*UTOB7ACK� /)�!�FRA:\�n X?n� '�`�0n�8� ��;�  2�0/07/31 �12:49:12ne(nO OMODO�<��mO�O�O�O�O�O�On��O_._@_ R_d_v__�_�_�_�_ �_�_o�_*o<oNo`o ro�oo�o�o�o�o�o����  �1_�p3_\ATBCK?CTL.TM;�S�ew��b;INI◰�5�&j3MESSAG� �q�!7 �#|�!�qODE_D� �&�%�xO��j3�PAUS`� !��/+ , 	��e /%d�r�,		\������������� ڏ��� �J�4�n�X��z���7�A�TSK � G��?�m0UP3DT�p�wd���XWZD_ENB8�t�*�STA�u/!��!!XIS� UN�T 2ǖ�!� �� 	 ��l��J7C�� ��� ]��� �n
|����T��!"�������,��Я�|�G�P� �b u�+� %M> A8R ��N'ȯ)��M��+^�MET��2�j��� P{�B9�5@�-A�B�4@��A/��yB"�v7�>��8=�&�=��Q�<�I=?��*��7_�SCRDCFG 1/%;�1 ��%�"E��+�=�O�a�s��?n
Q�)������� ���߄�Aߨ�e�w� �ߛ߭߿�&�`�'p1�GRc��%���6pN5A0.+	p4�ַ_ED�p1�� 
 �%-<pEDT-��*:|��6��Y�#��f�q2o�n
e"cO6h������2�);�� l�*��q1:���������"�
�3��M�*q� ��q����`��
�4��=���= ��,�
�5u� �	���	/Pb��
�6A/��/����j/�//./�/R/
�7 ?}/Z?�/��6?�?�/�/�??
�8�?��&O��]��OmO�?�?\O��?
�9�OO�O9O` ���O9_�O�O(_�O
�CR�H?�_�_~=�_�oJ_\_�_�_��K�N�O_DEL
��GE_UNUSE���IGALLOW� 1.�   �(*SYST�EM*4�	$S?ERV_GRE{�`nA�REG�e$�c4��`NUM�js�m�PMUi`4��LAYu�4��PMPAL�p?uCOYC10Jn]~Gp<K~�sULSU=�m�_rA��cL��tB�OXORI�eCU�R_�p�mPMC�NV9v�p10|s~%�T4DLI%����i	*PROG�RA�dPG_cMIK~u���ALU����~���B���n�$FLUI_RE�SUcw��o�!�MR�n�`lo,�e� w���������џ��� ��+�=�O�a�s��� ������ͯ߯����'�9�K�]�o���\bL�AL_OUT ��k���WD_A�BORdp�n���I�TR_RTN  �T��i�NONgSTOB�� ���CCFS_UTI�L .���CC�_AUXAXISw 3N� h����Ϧϸ�����CE_�RIA_I�`��Кa@�FCF�G N�Y�M��
�_LIM�b2�U� �P� 	���B\��TP
����Y�ZU�Y������Թ��`Yq��Q��$��v��X
_��"�9�PA�̀GP 1r�#��k�}���`�C�`C�@C7��J���]��p�������� C�����প���������̪������������������;���pCkT�������������������������������� D�� DK�K��K�K� �V?��3�HE8`ONFI�-��m�G_P�1r� Uerŷ� ��������#5m��KPAUS�q1r�� sr7}r� k����� �9IoU����?�Aii�4��M�NFO 1vH�$� �]�x9/T^��h>FQϿ]/�A/�� �D&t�����D)�³��?²E�´x/�)@�O� �*ز!�LLECT_�!0H��ذ#�#ENU�Ÿ�b�Ҳ!NDE�#�#H�Y�12�34567890�I7R�a$�G?Y6��H��S)�?�?�\�?�? �?�[�?�?BOOO1O �OUOgOyO�O�O�O�O _�O�O	_b_-_?_Q_ �_u_�_�_�_�_�_�_�:oo#6B�$�+ ��-'2IO &29��k#Ƽo�o�ol�o�gTR?�2'nm�(�؈2o ~x�(�m*z-��&_MORS�3)r͌a��u]� �y�������rT:�q*r�,}�?f�f�f���Kp���4�%P,2,�/.�e／ Ώ�������8u�k)@o,�k#� � ja�(P�DB.0.ʼ)dc?pmidbg]���L��ʓ:�n��p��|��Ȗ  �n��A��X�!��l����f�mgz�ӯ�� �f¯�� �>-`ud1:@�i��+ꂑDEF -���c)T�cy�b?uf.txtt��u���=�/nm��>�����a�MC&�r20��|cdC�$��s212ͤ!�q�k&�CzkЎ1^�A���hAӡ�A��߈B5O����C�4 y�H+C3/��C%;]C���D}�C����D�F-Ev��@F?�UE�f�E�v�E�/F��n�?���l�<�23nlD�)�h1��!��2�ӧ�5���
&pxc������ D4q��λ�G��  E%q��F�� E�p����F-F�P E���fF3H ?��GM����_�>�33��i�G��nc�G�@�5�����G�Ai�k$=L_��<#�{u�`�V��c:��RSMOFST +����EP_T1�4�nmA g���MO�DE 5���`���3q�w!;�-��O�I�?���<�{MܾTEST��)2����R�"6�/y��uƦ� Al�k(�� �b���C�0B͖��CE�������:d�{s +���*!����^��T_��PROG %G�%ӿL[��`�NUSER�`K�EY_TBL  �G�!$"�	
��� !"#�$%&'()*+�,-./R7:;<=>?@ABC���GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������&��������������������������������������������������������������  L�CKjp�aj ST�AT�\�X1_A�L-�p1}_AU_TO_DO6o�~#FDR 38��2hk)U;`/r/�/�$O/�/H�-�k� �/5����)�/�/�/<? >O?5�\�J�N/�?�? �?�/�?!Oe�T���8O bOh3fOPO�O�OnO�O �O�O
]�?/_A_S_�? d_�_4O�_�_�O�_�_ �_�_�_o(o^opo_ �o�o�of_�o�o�_ *o,Xf<z ����o��#��o 4�Y�z�t������ ��Ώ�����.�@�� g�y���6�����l�� ܟ�����(�6��J� `�����V�ϯ�󯞟 �)�ԟJ�D�b�d�V� ����t���ȿ��Ͼ� 7�I�[��lϑ�<��� ��ʿ�Ͼ������� 0�f�x�&ϟ߱���n� ���ߤ���2�4�&� `�n�D�������� ��+���<�a��� |��������������  6H��o��>� ��t���� 0>Rh��^ ����/1/�R/ L/jl/^/�/�/|/�/ �/??�??Q?c?/ t?�?D/�?�?�/�?�?  OO�?"O8OnO�O.? �O�O�Ov?�O_�?"_ _:O<_._h_v_L_�_ �_�_�_�Oo!o3o�O Doio_�o�o�_�o�o �o�o�o�o>P�_ w��Fo��|o� �
��8�F��Z� p�����fߏ��� �9��Z�T�r�t�f� ������؟� �Ώ G�Y�k��|���L�¯ ��ڟܯί���*� @�v���6�����ӿ~� �	ϴ�*�$�B�D�6� p�~�TϒϨ����Ϟ� �)�;��L�q�ϒ� �ߪϬߞ����߼��� �F�X�����N� ������������ @�N�$�b�x�����n� ������A��b \z�|n���� �(��Oas ��T����� //�2/H/~/�/> �/�/�/��/?�2? ,?J/L?>?x?�?\?�? �?�?�?�/O1OCO�/ TOyO$?�O�O�?�O�O �O�O�O__N_`_O �_�_�_VO�_�_�Oo �__ooHoVo,ojo �o�o�ov_�o�_ $I�_jd�o�v ������0��o W�i�{�&����\ҏ ̏��ޏ�&���:� P�����F���џ㟎� ���ď:�4�R�T�F� ����d������ ��� '�9�K���\���,��� �����������̿
�  �V�h���ϡϳ�^� ���ϔ�
��"�$�� P�^�4�r߈߾���~� ��	����,�Q���r� l�ߌ�~������� ��&�8���_�q���.� ����d�����������  .BX��N� ������!��B <Z\N��l� ��/�//A/S/� d/�/4�/�/��/�/ �/�/�/?(?^?p?/ �?�?�?f/�?�?�/O O*?,OOXOfO<OzO �O�O�O�?�O_#_�? 4_Y_Oz_t_�O�_�_ �_�_�_�_�_.o@o�O goyo�o6_�o�ol_�o �o�_�o�o(6J `��Vo����o �)��oJ�D�bd�V� ����t���ȏ���� 7�I�[��l���<��� ��ʏ̟�����ܟ� 0�f�x�&�����ïn� ԯ������2�4�&� `�n�D�����ο࿎� ��+�֯<�a���� |Ϛ��ώ����Ϭ���  �6�H���o߁ߓ�>� ����t��������� 0�>��R�h���^� ��������1���R� L�j�l�^�����|��� ����?Qc� t�D�������  �"8n�. ���v�/�"/ /:</./h/v/L/�/ �/�/�/�?!?3?� D?i?/�?�?�/�?�? �?�?�?�?O>OPO�/ wO�O�OF?�O�O|?�O �O
O_�O8_F__Z_ p_�_�_fO�_�_o�O o9o�OZoTor_tofo �o�o�o�o�o �_ GYko|�Lo� ��o�����*��@�v�\��$CR_�FDR_CFG �9Z�~�q
UD1:�w:�tJƄ  Ҁ�|���HIST 3:�Z�  ��  w?�r@�UA�B�C�p�UD�E�I�g�p�o�w�h���INDT_EN���t������T1_DO c �u��z�T2��~��VAR 2;����� h�� � A&���&��r��'L�'L�΍C��rZ��STO�P����TRL_D�ELET6�Ɣ �n�_SCREEN� Z���k�cscy�U_�MM�ENU 1<��_  <�|%� ���tۯ�:��s�=� v�M�_�������⿹� ˿�*���`�7�I� ��m�ϥ��ϵ���� ����J�!�3�Yߒ�i� {��ߟ߱�������� F��/�|�S�e��� ����������0��� f�=�O�u��������� ������)b9 K�o����� ��L#5�Y k���� /�y��?_MANUA3�e�n��ZCD��=㙼��/%  "��r�Ԇ
*n'
*?|(���pd<'GRP �2>��B� h ���"h ��$DBCO��RI�G�����"G_ERRLOG ?ʫ²q�/1?C?U? ~�!NUMLIMē��!��
�!PXW�ORK 1@ʫ� ?�?�?�?�?�?m�D�BTB_y� A=���!;Bl ��DB_AWAY�#��qGCP ��=s�ׇ2UB_ALs0..�"_�"Yb��������S@ 0 1B�+ , 
�?�O
$�O�_H_M���_L@}�%UONTIM�������GV�I
�}P�GMOTNE�N.�.&}[RECO�RD 2Hʫ y�_�sG�O��Q �_
+`B	oo-o?o�X Gono�_�oo�o�o�o qo�oo4�oXj |�)�!�E� ��0��T��x�� ������ҏA���e�� ��>�P�b�t�㏘�� ��+��������:� ��3�͟��������'� ܯǯկ�����J� \�˯��k�y���%�7� ���m�"�ϣ�X�ǿ ٿ�Ϡ�7ϯ���E��� i�{�0�B�����x��� ���������ߑ�QB�TOLERENC�^DBȧBl@L���� CSS_CCS_CB 2I�,DP
$�O
.c���� ?�������(�:�L��p���
+�`����� ������!3EW i{������ �/ASew �������/ /+/=/O/a/s/�/�/C ���/�/���+V:�LLE�JI�UQ|<C9 C���C�{0.0��F? A��+�p+ഄC�P��q1�- 	 A��k0�0B�ߍ9?�  �6��?�?�(DPc��qP��B��րHC[�3OEOWO��{O�(kO�O[O�OO���K��L�d������?�8;V�ȥ[D�O���OH_#2��@��7_�_�_�_���vPA.��_c8.�A  �_o�WqQm1�1m1!m�QB�QBoLb)e�YoP�o�o�oQZP��`�`�0�D20Ca�� @��
�!X8N�k   5_��>7�����Yk}�"w�a$1W2�!"{$5 �ךO��O��8�0J�\���MaCH+�>1��?3B�Dz��D ~���%O��ď�ݏ��K	���2%���"�CR�A�P�W 1_�/�t��=R�t�r� R���ʟ����Пޟ�9��#�q`H������ ���a����*3Ʃ��� ���!��E�W�6�{� Z�l���ÿ�o�b�"���q2��Az&�4���B7YB#��@�m@$Y*���ʿB�T�f�x����"Hy`^���� ���ϊϴ�!��E�W� i��0ߝߐ�����r� �߮��-�?�Q��u� �����߆����� �)�;���_�>�P���`t��s����x�  h���0'9f] o������� �,��OY�} �������(/ /1/K/U/�/���/�/  z/���/�/? ?5?(?Y?L?^?�?�? �?�?�?�?�?�? O1O 8UOt/^O�O�O�O�O �O�O�O�O__$_Q_ H_Z_�_FO�_�_�_�_ �_�_oo o2oDoqo�hozo�o�o�o�oԷ	o  �a��`�����`�/- R=va�C�' �<�q
S�����h�:�2����#��K�����i�A�   ����m�@�C  Տ�͂С���Ѡ=�賖 ���Ͽ�+Ă�C��  M�3�t��~Ӄ>�{�����S��@@��������B�S�>����C�������͂��<��o?�PH�)S�B����������Bܿ�ͅ1�"+��9�� m�b��i�20K��5��!��@�	�@$X��9����B]A��
�y�@q.^B]���т��¡` � ?��ͥͿ�u�{?����e�ܱ�Ծ��$DCSS_CL�LB2 2K�����p�~'�NSTCY 2L����  h�믊�������ҿ �����,�B�P�b� tϊϘϪϼ��Ϸs)��DEVICE 2%Mm���(�� >�P�}�t߆߳ߪ߼� ��������C�:�g�y�������)�HNDGD Nm���Cz�k)�LS 2Om�G�9�K�]��o�����������PA?RAM P8�����H��RBT 2}Rm� 8�p	<	������Q�T������R��1ʹ@� �CW  �B\`6怈B	�� ���� �@R����b��I������. ���	>,�YkJk����c��; M� T����0///f/��A�S�D �C��ׂ!т1�@#��@I&��@R�\@g�;�?��j��B�&�fB�DC�C3$C2��oC3Ф����A���B8��yBB�A��.���mB���C��RC3�C4
_C3��a�(�35P<8�@"E/W/ �??/m??�?�?�?O �?�?8OO!O3OEOWO iO�O�O�O�O�O�O�O �O__j_A_S_�_�_ l��_�_�_�_o	oBo To?oxo�[?�_�_q_ �o�o�o�o�o4 /ASe���� ������f�=� O���s������_o� �,��)�b�M���q� ���o��ŏ򟭏۟� :��#�p�G�Y���}� �����ůׯ$���� Z�1�C�U���y���ؿ ����� ϛ�D�/�h� Sό�wω��ϭ����� ��.���)�;�M� _߬߃ߕ��߹����� ����`�7�I��m� ����������� J�\��π�k������� ��������"��+�=� jAS�w��� ���T+= Oas����/ ��//'/9/�/ �/�/�/�/�/?�/(? ?L?^?9g/y/�?}? �?�?�?�?O�?�?O ZO1OCO�OgOyO�O�O �O�O_�O�OD__-_ z_Q_c_u_�_=?�_�_ 
ooo@o+odoOo�o c?u?�_�o�_�o�o �oN%7I[m ������� �!�3���W�i����� ������yo"��F�1��j�|�g�����ğ�h��$DCSS_SL�AVE S������~ښ_4D  ���AR_MENU T� ��R�d� v��������bA�֯��֞'�SHOW �2U� �  ��Ձ/�9�@�^�p������������ܿ� �  (�"�L�I�[�m�ϑ� ��ʿ��������6� 3�E�W�i�{ߍߴϱ� �������� ��/�A� S�e�w�ߛ����� ��
���+�=�O�a� ��������������� '9Kr�[� ��������� #5\�k}�� �����//1/ XU/g/���w/�/ �/�/�/	??B/??Q? x/�/�/2?�?�?�?�? �?O,?)O;OMOt?nO �?�O�O�O�O�O�OO _%_7_^OX_�O_�_ �_�_�_�_ _�_o!o H_Bol_io{o�o�o�o �o�_�o�o2o,Vo Sew����o� ���@=�O�a� s��������͏ߏ�  �*�'�9�K�]�o���ਏ"���ɟ��CFG7 V������FRA�:\	�L�%04_d.CSV�	��m}֟ ���A O�CHW�z��g�񏋯���  �u������į֯�u����JP����u��������RC_O�UT W�����+�۟_C_F�SI ?Q� �u����� ��޿ٿ���&�!�3� E�n�i�{ύ϶ϱ��� ��������F�A�S� eߎ߉ߛ߭������� ����+�=�f�a�s� ������������ �>�9�K�]������� ����������# 5^Yk}��� ����61C U~y����� �/	//-/V/Q/c/ u/�/�/�/�/�/�/�/ ?.?)?;?M?v?q?�? �?�?�?�?�?OOO %ONOIO[OmO�O�O�O �O�O�O�O�O&_!_3_ E_n_i_{_�_�_�_�_ �_�_�_ooFoAoSo eo�o�o�o�o�o�o�o �o+=fas �������� �>�9�K�]������� ��Ώɏۏ���#� 5�^�Y�k�}������� ş�����6�1�C� U�~�y�����Ư��ӯ ��	��-�V�Q�c� u������������ �.�)�;�M�v�qσ� �ϾϹ�������� %�N�I�[�mߖߑߣ� ����������&�!�3� E�n�i�{������ ��������F�A�S� e��������������� ��+=fas ������� >9K]��� �����//#/ 5/^/Y/k/}/�/�/�/ �/�/�/�/?6?1?C? U?~?y?�?�?�?�?�? �?O	OO-OVOQOcO uO�O�O�O�O�O�O�C��$DCS_C_�FSO ?����Q P �O�O<_e_ `_r_�_�_�_�_�_�_ �_oo=o8oJo\o�o �o�o�o�o�o�o�o "4]Xj|� �������5� 0�B�T�}�x�����ŏ ��ҏ����,�U� P�b�t���������� ����-�(�:�L�u� p���������ʯܯ�  ��$�M�H�Z�l��� ������ݿؿ���%π �2�D�m�h�z�_C/_RPI^._�� ����Ϩ�_���W�X��{�^SL��@L� ���� �����H�C� U�g��������� ���� ��-�?�h�c� u��������������� @;M_�� ������ %7`[m�� �����/8/3/ E/W/�/{/�/�/�/�/ �/�/???/?X?S? e?w?�?�?��9��߬? �?OO+O=OfOaOsO �O�O�O�O�O�O�O_ _>_9_K_]_�_�_�_ �_�_�_�_�_oo#o 5o^oYoko}o�o�o�o �o�o�o�o61C U~y����� ��	��-�V�Q�c� u������������ �.�)�;�M�v�q���𕟾���&�NOCO�DE X=���'�PRE_?CHK Z=�А�A А�< �Ր=�E�W�=� 	 <9������3 y�ïկ�������� A�S�-�w���c����� ��������+�=�� a�s�i�[ϩϻ�U��� ������'���]�o� Iߓߥ�߱��ߵ��� �#���G�Y�3�e�� �ϗ�����q������ ��C�U�/�y���e��� ��������	��-? KuOa��� �����);_ qK������ �/%/�I/[/5/G/ �/�/}/�/�/�/�/? �/E?W?�/{?�?g? �?�?�?�?�?O�?/O AOOMOwOQOcO�O�O �O�O�O�O_+_!?3? a_s___�_�_�_�_ �_�_o'oo3o]o7o Io�o�oo�o�o�o�o �o�oGY3}� I_w������ 1�C��/�y���e��� �������я�-�?� �c�u�O�������� �󟍟�)��5�_� 9�K�������˯ݯ�� �����I�[�5�� ��k���ǿ��ϟ��� ���E��1�{ύ�g� ���ϝ���������/� A��e�w�Q߃߭߇� ���������+��� a�s�M�������� �����'��K�]�7� ����m���������� ��5G=�/}� )������� 1CgyS�� �����/-// 9/c/Yk�/�/E/�/ �/�/�/?)??M?_? 9?k?�?o?�?�?�?�? OO�?OIO#O5OO �OkO�O�O�/�O�O_ �O3_E__i_{_U_g_ �_�_�_�_�_�_o/o 	ooeowoQo�o�o�o �o�o�O�o+�oO a;m�q��� ����!�K�%�7� ����m���ɏ��Տ�� �o5�G��S�}�W� i���ş�����՟� 1���g�y�S����� ����寿�ѯ�-�� Q�c��K�������Ͽ Ώ�����M�_� 9σϕ�oϹ��ϥϷ� ����7�I�#�m�� u�gߵ���a������� 	�3���i�{�U�� �����������/� 	�S�e�?�q����ߣ� ����}�����O a;��q��� ��9K%W �[m����� ���5/G/!/k/}/W/ �/�/�/�/�/�/�/? 1??U?g?A?S?�?�? �?�?�?�?	OO/O QOcO�?�O�OsO�O�O �O�O__�O;_M_'_ Y_�_]_o_�_�_�_�_ o�_o7o-O?Omoo o�o�o�o�o�o�o�o !3?iCU� �������� 	�S�e�?�����Uo�� я㏽����=�O� )�;�����q���͟�� ��ݟ�9�K�%�o� ��[������������ ��#�5��A�k�E�W� ������׿�ÿ��� ���U�g�Aϋϝ�w� ����ɯۯ	�ߵ�'� Q�+�=߇ߙ�s߽��� ���������;�M�'� q��]������������$DCS_SGN [���-��^�>	�29-NOV-�25 10:31� ��6�0- 7-�E�  12:49� `�`� [�}S�n�P�f4�n�j�`��k�2�ե��U�Þ�;"�0>~�  �HO�W \��� `��VE�RSION �%�V4.5.�2��EFLOGI�C 1]���  	������+	���:PROG_E_NB  ��"�c�[ULSE  �@s_AC�CLIM���ud�WRSTgJNT�-���EMOdb�w� INIT ^
����OPT_S�L ?	���
 	R575��VE74J6K7K50o1o +	�|(TO  4���V� DEX҆d-�`�#PA�TH A%�A�\�S/e/��HCP�_CLNTID y?��" ,����/��IAG_G�RP 2c������b�	 �@�  �"ff�?aG��%��� BG�  ?��1� 0�C?1>@c��j2!��7@�z�@^��@
�!���mp2m15 �89012345�67�0���� � ?��?��=q?��
?���R?�Q�?ѯ�?ʼ0��0�?(�?�z���0�`�@�  AG�A�p�0�10A� 0� 0G�B4�� ��4`�
�1@����@��\@~��R@xQ�@q���@j�H@c��
@\��@U�@Mp����?�?�D��#@��7IH���@C\@>L@9���@4x0/\)@)��@#\@{@�jO|O�O�O�O8G�?���?��0��� G@?}p�?u?n{?[@;?\�0Q��O_�_,_>_PX�
=?���0�tP_U� 0z��H?p�0h��?^�R�_�_�_�_��_PX�5�\P�� �� 0� `�0?�tP� � #`o o2oDoVo8G ����oAS�o' q�y��[m� �+�	�O�a��m��ÀqbRB�@jRcQ�`
=?��ʆ�\Pׄ
=�5!��4V����
=�b��a&���U?� @C��``3�=q�=b���=�E1>�J��>�n�>��H�
=<�o ~��s������ �`�C޷`<(�Ub� �4�"��@ß���A@`�?5������ 8�J��Ȼ�V������ද��گ쯖�>J����bN�
=�'�G�6���@{`^��pP��0k�@f�fZ>!T@��33�푒�(��
=C��� ��I�CH��)C.dB؃�
= B׿ݱɼ' �  �
��a'�B3Ğ�,��N�B��`�X���wωϰ���3~���l�_?�(�k�R������!�`�~�lD&t�����D/�`�>�s���o�ߢ˻6�<҂������ ²X����AD
� ��߯ߚ��߾��������n��*Iҥ	��W��!CT_CON�FIG d�'|�d�egA��!STBF_TTS�
s	�����e�:���MAU� h~��MSW_CFv��e�+  ��OCoVIEW��f	�1���/[�m���� ������I����� &8��\n��� �E���"4 F�j|���� S��//0/B/� f/x/�/�/�/�/�/a/ �/??,?>?P?�/t?��?�?�?�?�?^�RC�gΥ��!j?NO ;O*O_ONO�OrO�O���SBL_FAUL�T h�:��AG�PMSK���Gj�TDIAG iz��������UD1: 67890123451R��%Q��EPD�m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�oLV�!V�i�
\_�od�TORECP
_Z
*T CW5{[_Xj|� �������� 0�B�T�f�x��o�o�o����UMP_OP�TIO%��NځT�R���I��PM�E���Y_TEM�P  È�3�B+�O��*�9�U�NI���O���YN_BRK j4�~�EDITOR����(���_�`ENT� 1k�9  �,&IP�ANU�C_SMPLGRP_CLOSEȏ�&FS_MOV_5DEG �'OPE%��������EAS_W�RK2FpG��A�NIMA�_DR�Oq�W��30�K��� �-BCKE�DT- _PIC�ɯ��HOME ��*�&PROG_1 �������|J��MAIN q�>��&DE�C����GETDATA4˿ݿ��1 ���&&�1 �B���AAA �R���&�y϶��TE�� 4?���@�1 ����&�O4�1䜐MGDI_STAb�>�O���✐NC_INF�O 1l	������@����ߢ�n�V�;1m	� �~������
�d��=�O� a�s��������� ����'�9�K�]�o� ��������������� 	*�8J\n �������� "4FXj|� �
�����/! +/=/O/a/s/�/�/�/ �/�/�/�/??'?9? K?]?o?�?�?�?��? �?�?�?/#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�?�_�_�_�_O o-o?oQocouo�o�o �o�o�o�o�o) ;M_q���_�_ ����o%�7�I� [�m��������Ǐُ ����!�3�E�W�i� {�����ß՟��� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9� K�]�oρϓϥϷ��� �������#�5�G�Y� k�}ߏߩ��������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u����� �����������) ;M_q���� ���%7I [m������� �/!/3/E/W/i/ {/�/�/�/�/�/�/�/ ??/?A?S?e?w?� ��?�?�?�?�OO +O=OOOaOsO�O�O�O �O�O�O�O__'_9_ K_]_o_�_�?�_�_�_ �_�?�_o#o5oGoYo ko}o�o�o�o�o�o�o �o1CUgy �_�����_�	� �-�?�Q�c�u����� ����Ϗ����)� ;�M�_�q������� ˟�����%�7�I� [�m��������ǯٯ ����!�3�E�W�i� ��������ÿտ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�sߍ��ߩ� ���������'�9� K�]�o������� �������#�5�G�Y� k��ߏ����������� ��1CUgy �������	 -?Qc}�o� �������//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?u��?�?�?�?� �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_�??�_ �_�_�_�?�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]w_�����_ ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�o]� ������������	� �-�?�Q�c�u����� ����ϯ����)� ;�M�g�y�������]� ӟݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�_�q� {ߍߟ߱�˿������ ��/�A�S�e�w�� ������������ +�=�O�i�s������� ��������'9 K]o����� ���#5Ga� k}������� �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???YK?u?�?�? ���?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_Q? c?m__�_�_�?�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /�_[_ew� ��_������ +�=�O�a�s������� ��͏ߏ���'�9� S]�o��������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�K�9�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)��C� �$ENETMODE 1n����  S�S�N�p߂��R�OATCFG {o��������C���DA_TA 1p_���]���*��*�� �!�3�E�T�dT�u���M�y������� ��������E�W�i� {��������=����� /A����w� �����]o +=Oas�� ����//�� K/]/o/�/�/�/�-R��RPOST_LO��r��C%
���/?�?/?Q�RROR_[PR� %_�%4/�q?@8TABLE  _����?�?�?��+RSEV_NU�M n�  ��i�@�!_AU�TO_ENB  q��g�@4_NOA� s_ہ�B�  *�`@�`@�`@�`@@+_@yO�O<�O9DFLTR%O7F�HISCE!g�2K_�ALM 1t_�� �C$`LM�+ �O9_K_]_o_�_�_�O�_�2?@  _��^A���ZR�TCP_�VER !_�!�`?�_$EXT� _7REQ�F�0I*c�SIZ3o%dSTK�PiNE�'bTOoL  E!Dz�B��A %d_BW�D�P�`�F�a�ҢcDI�a u���'��<E!�kSTEP�o�o|R��`OP_DOro�P�FDR_GRP� 1v_��Ad 	��_p��aps�Y��q'�M"����l��T� ����vas���}�tA
�A��IZA$@�����{��{/���?�e�P���t����}?�԰W@/Ơ@9�?��ܷ�
 F@ �q<ԁE!@	���R�����B�-�f�Q�A@<�p��@S33��P�@����O�؟�ap�x �ŜapG�  (��Fg�fC�8R�4�ȝ?�΀Q�Ǟ6��X�x��875�t��5���5�`+�ȟH �������%V��ArEATURE� w���`���LR Han�dlingToo�l �E"En�glish Di�ctionary���Multi L�anguage ?(CHIN)�&��KANA/�4D ;St�ard����Analog I�/O^�g�gle �Shiftz�ut�o Softwa�re Updat�e��matic ?Backup�ͱ�ground E�dit���Cam�erau�Fy�Co�mmon cal�ib UI��n���Monito�r(�tr�Rel�iab����DHC�P��Data ?Acquis7�`�?iagnosɱr�~z�isplay�?Licens^�d��ocument �VieweC�b�u�al Check Safety#�~��hanced#�4���s��Fr�����xt. DIO �3�fi��D�end.�ErrB�L��`�J8�s_�rp�O� �`��FCTN Me�nu�v^ò�TPw In��fac����GigE������p Mask Ecxc�'���HT���Proxy Sv���#�igh-Spe�Skiҳ#��~S�mmunicȰ7onsZ�ur�С��u�v���conne�ct 2��ncr��stru	�����e����J��0�KA�REL Cmd.� ���Run-Ti�@�Env���el� +̰sʰS/W���������v�Boo�k(System�)�MACROs�,Q�/Offse���0�HSв�s�5�MR<�8®�M����R��l��MechSt�op/�t����0�iqґ� x�r�ʰ���od��witch�.���.��TOpctmf��0�fi��2��g��0�-T����PCM funt���	a��tiz�z�o��Regii�Yru��ri��F��4s�Num Se�l��O>� Adj�ue�Jw���ta�tu0�����RDM Robot��scove��e�a�@�Freq �Anlyu�Rem���S�nU���Se�rvoS�A ��SN�PX b1�SN���Cli��_.��LGibr�/� ԑ K&oN�t��ss#ag�0��P �����a��P/I���%MI�LIB?�"P F�irm���.P��A�cc��TPTXo��$eln��?�!x��-orqu��imulaA���6uH Pa*��.�\�:b&/�ev.�%���ri��t?USR� EVNTO-@n?except� an��(E9�{�VC�rp�g���V���B<?h�E�+�KSr SCn5��OSGE�O�EUI~a�Web Pl� ^=!��ET7�������ZDT Applxn��QEOAT�!,Ѵ��iPj�ax)�_ Grid����].�_iR�B.U�f����O��RX-10�iA�_m�ll SmoothU���c��scii/�vLosad��tjUpl�`Η�toS��0ri�tyAvoidM�,�sW�t�0g`	�y�c���;@�c�C9S/�. c�� xJo=tL�r� x�u��� xc��a3bo���RL�0>�2Y��or��O�0��S�Fit��{tl�nt���wHMIo Dev�� (S!m� d��in�#?�
<���sswo\����ROS Eth (��a�!��$�[L%�ga �b�L%dhUpv�E!�%[�t �Нi�Rs��{�64MB� DRAM��F�RO#����l<f F!lH����6m �aZ�opq���e``v��#sh����Ɨc�Õ���p�6؜ty��sa�)�r'��j"b~ .z�pq/sJs��d� �vx��� 2:�ap�pornv�h�<"V�q�T1*�cFC/��E�Fs=Ȏ�Hel�U!��T[yp��FCE h�фvR@St�{����l�uA $ꃨPG �j����Rj��No� m �c߷ dOL;�Sup���0�OPC-UJk"�T�遼�5��j��cr.p�lu� �����quir��� Om���%�T0.
���es�tL%IMPLE ���VJ'S;�eq�tCex��dhz�I(p��[B�?CPP���E8����bTeaH �9�ߚDrtu���v�Yp���4���UIFg��ponsRfstd�pnKe SWI�MEST f� F	01ᚥ� bC�:�L� y�p��������� 	� ��?�6�H�u�l� ~������������� ;2Dqhz� �����
7 .@mdv��� ����/3/*/</ i/`/r/�/�/�/�/�/ �/�/?/?&?8?e?\? n?�?�?�?�?�?�?�? �?+O"O4OaOXOjO�O �O�O�O�O�O�O�O'_ _0_]_T_f_�_�_�_ �_�_�_�_�_#oo,o YoPobo�o�o�o�o�o �o�o�o(UL ^������� ���$�Q�H�Z��� ~��������؏�� � �M�D�V���z��� ����ݟԟ��
�� I�@�R��v������� ٯЯ����E�<� N�{�r�������տ̿ ޿���A�8�J�w� nπϒϤ�������� ���=�4�F�s�j�|� �ߠ����������� 9�0�B�o�f�x��� �����������5�,� >�k�b�t��������� ������1(:g ^p������ � -$6cZl ~������� )/ /2/_/V/h/z/�/ �/�/�/�/�/�/%?? .?[?R?d?v?�?�?�? �?�?�?�?!OO*OWO NO`OrO�O�O�O�O�O �O�O__&_S_J_\_ n_�_�_�_�_�_�_�_ oo"oOoFoXojo|o �o�o�o�o�o�o KBTfx�� �������G� >�P�b�t�������׏ Ώ�����C�:�L� ^�p�������ӟʟܟ 	� ��?�6�H�Z�l� ������ϯƯد��� �;�2�D�V�h����� ��˿¿Կ���
�7� .�@�R�dϑψϚ��� ���������3�*�<� N�`ߍ߄ߖ��ߺ��� �����/�&�8�J�\� ������������ ��+�"�4�F�X���|� ��������������' 0BT�x�� �����#, >P}t���� ���//(/:/L/�y/p/�/�/�/�* � H551��#�!2�(39�(0^�%R782�'56�J614�%ATU]P'6545'86�%�VCAM�%CUI�F'728c6NREv652V6R63�&�RSCH�%LICކ6DOCV�6CS�U6866J60^26EIOC�746�R69V6ESET�?7U7J7U7R68��&MASK�%PR�XYo87�&OCOBH3?86@&83^F�J6%8 :�GLCH^FFOPLG?70vF�MHCRGFS�GM�AT�6MCS>80�"G5526MDSW�+WiGOPiGMPR�jF�0�H06PCM�n75qW@26�@�G5�1J751�X0J6P�RSG69^FFR�Db6FREQ6M�CN�&97SNByA�7�GSHLBf�M1g�0X26HT=C>6TMIL86�TPA�6TPTXFcfELf�@�787�0�&J95z6TU�TjFUEVFUE�CFFUFRb6VCuC�hO�FVIPnfwCSC�fCSG�6��0I�%WEB>6HTT>6R6�8�h;0�FvCG]wIGEwI�PGS�vRCnfD�GiGH7�X6�'Ru7	GR�XR51�8�6vH2vH5V6�0J�X�X6z7L=i�'J�87"G87�G83�J6R55vF@26Rk64�g5��R6�G�R84��79�H4vz6S5]GJ76^F�D0626F �RT�SfCRDFCR�XjFCLIZXI7C�MS�6S�>6STY:ng6)WCTO>6�0��77�7�0z6ORS��F7@6FCB�6F�CF�WCH>6FC�RFFCI�vFCR�GJ�pOWG*�M�X7NOM�6OLWKP��6OP��SENDvGFLU�FCPR�W�L	wS��C�8ETaS^�T��0zgCP�6�TE%�S60�&F�VR�6IN�WIH�agIPNnfGene�$�(1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹� ��������%�7�I� [�m��������� �����!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�w��� ������џ����� +�=�O�a�s����������ͩ  OH551ϧ�2��39��0�R78�2�5�J614��ATUP?�54�5?�6�VCAM��CUIF?�28n��NRE�52~��R63�RSCH��LIC��DOC�V��CSU�86��J60N�EIOuC��4.�R69~��ESET_�}�J7�}�R68�MAS�K�PRXY��7.�OCO�3_�.�4��>�3��J6=����LCH��OPL�G_�0��MHCR���S}�MAT��MkCS^�0��55N��MDSW����OP���MPR��۰.�0.�PCM��5M���N���.�51n�51���0n�PRS~�6�9��FRD��FR�EQ�MCN�9��SNBAϻ�SHLB�MM�۰���2�HTC^�TMsIL��TPAN�oTPTX��EL�ċ�.�8-�+��J9�5��TUT��UE�V~�UEC��UF]R��VCC^O��wVIP��CSC���CSG���I�W�EB^�HTT^�Ra6ͼ��[��
CG�{IG�IPGS�RC��DG��H7Zm�6�R7m�R��WR51^�6��2��I5~��J�ܞ�6���L]��J87��8�7.�83n�R55���k�N�R645v�+R6��R84n+k79�4��S5��wJ76��D06N��F<RTS.�CR�D~�CRX��CL9I.�m�CMSN�{0�^�STY��6��C#TO^��N�7-�˰���ORS�ګ��F�CBN�FCF��C�H^�FCR~�FC-I>FC��J�uG�M��NOMN�cOL����OP]KoSEND��LU~�WCPR��LmS�<C�ETS�K|<;����CP��TE=;S�60�FVRN�I�N��IH��IPN��Gene�Ψ�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� ������������ '9K]o��� �����#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů�  נST�DҤLANG ����0�B�T�f� x���������ҿ��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V��h�z�������RB=T�OPTN���� ��	-?Qcu��������DPN�);M _q������ �//%/7/I/[/m/ /�/�/�/�/�/�/�/~?ted � ʨ9?K?]?o?�?�?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_�_�_�_�_ �_	oo-o?oQocouo �o�o�o�o�o�o�o );M_q�� �������%� 7�I�[�m�������� Ǐُ����!�3�E� W�i�{�������ß՟ �����/�A�S�e� w���������ѯ��� ��+�=�O�a�s��� ������Ϳ߿��� '�9�K�]�oρϓϥ� �����������#�5� G�Y�k�}ߏߡ߳��� ��������1�C�U� g�y���������� ��	��-�?�Q�c�u� �������������� );M_q�� �����% 7I[m��� ����/!/3/E/  �N/l/~/�/�/ܴ/�-99�%�$�FEAT_ADD ?	����!�0  	 �(??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q������� ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ�������� �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o�������������$DEMO� w�)   �(4�*�<�i�`� r��������������� /&8e\n� �������+ "4aXj��� �����'//0/ ]/T/f/�/�/�/�/�/ �/�/�/#??,?Y?P? b?�?�?�?�?�?�?�? �?OO(OUOLO^O�O �O�O�O�O�O�O�O_ _$_Q_H_Z_�_~_�_ �_�_�_�_�_oo o MoDoVo�ozo�o�o�o �o�o�o
I@ Rv����� ����E�<�N�{� r���������ԏޏ� ��A�8�J�w�n��� ������Пڟ���� =�4�F�s�j�|����� ��̯֯����9�0� B�o�f�x�������ȿ ҿ�����5�,�>�k� b�tϡϘϪ������� ���1�(�:�g�^�p� �ߔߦ��������� � -�$�6�c�Z�l��� �����������)� � 2�_�V�h��������� ��������%.[ Rd������ ��!*WN` �������� //&/S/J/\/�/�/ �/�/�/�/�/�/?? "?O?F?X?�?|?�?�? �?�?�?�?OOOKO BOTO�OxO�O�O�O�O �O�O___G_>_P_ }_t_�_�_�_�_�_�_ oooCo:oLoyopo �o�o�o�o�o�o	  ?6Hul~� �������;� 2�D�q�h�z�����ˏ ԏ���
�7�.�@� m�d�v�����ǟ��П �����3�*�<�i�`� r�����ï��̯��� �/�&�8�e�\�n��� ������ȿ�����+� "�4�a�X�jτώϻ� ����������'��0� ]�T�f߀ߊ߷߮��� ������#��,�Y�P� b�|��������� ����(�U�L�^�x� �������������� $QHZt~� �����  MDVpz��� ���/
//I/@/ R/l/v/�/�/�/�/�/ �/???E?<?N?h? r?�?�?�?�?�?�?O OOAO8OJOdOnO�O �O�O�O�O�O_�O_ =_4_F_`_j_�_�_�_ �_�_�_o�_o9o0o Bo\ofo�o�o�o�o�o �o�o�o5,>X b������� ��1�(�:�T�^��� ��������ʏ��� � -�$�6�P�Z���~��� ����Ɵ����)� � 2�L�V���z������� ¯����%��.�H� R��v���������� ���!��*�D�N�{� rτϱϨϺ������� ��&�@�J�w�n߀� �ߤ߶��������� "�<�F�s�j�|��� �����������8� B�o�f�x��������� ����4>k bt������ 0:g^p ������	/ / /,/6/c/Z/l/�/�/ �/�/�/�/?�/?(? 2?_?V?h?�?�?�?�? �?�?O�?
O$O.O[O ROdO�O�O�O�O�O�O �O�O_ _*_W_N_`_ �_�_�_�_�_�_�_�_ oo&oSoJo\o�o�o��o�o�o�o�o�o}  x.@R dv������ ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t�����������|��  � �2�D�V�h�z����� ����������
. @Rdv���� ���*<N `r������ �//&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� ��6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L ^p������ � ��$�6�H�Z�l� ~�������Ə؏��� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я�����*�<� N�`�r���������̿ ޿���&�8�J�\� nπϒϤ϶������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ������������,� >�P�b�t��������� ������(:L ^p������ � $6HZl ~������� / /2/D/V/h/z/�/ �/�/�/�/�/�/
?? .?@?R?d?v?�?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O �O�O__&_8_J_\_ n_�_�_�_�_�_�_�_ �_o"o4oFoXojo|o �o�o�o�o�o�o�o�y�$FEAT_�DEMOIN  �#t�Np�$p�6tINDEXC{�Rq�6pILECO�MP x����qQr1uzp�SETUP2 �y�u�r� � N �qws_AP2BCK 1z�y?  �)x�"�{%� �$p�p� K�!u�w����*��� я`������+���O� ޏs������8�͟ߟ n����'���4�]�� �������F�ۯj��� ���5�įY�k����� ���B����x�Ϝ� 1�C�ҿg����ϝ�,� ��P����φ�ߪ�?� ��L�u�ߙ�(߽��� ^��߂��)��M��� q����6���Z��� ���%���I�[���� �����D���h��� ��3��W��d� �@��v�/ A�e���*��N�r�/�y�pP�� 2�p*.cVR /j/�*m/��/��/�/�T PC��/�/�FR6:D�/>�/>?�+Tbp b?t?5_?�<Ep/?�?�*.FW/�?�	3�?"L�?FO�;STMQO{O20gO"�M5O�O�;H�O�O��G�O�O�OO_�:GIFY_�_�Eo_,_>_�_�:JPG�_o�E�_0�_�_Wo�*JSao�o��cxo5o%
J�avaScript�o�_CS�o�F��o�o %Cas�cading S�tyle She�ets:�
AR�GNAME.DTi��@\};�a�t�j�pDISP*���t����q4�B��CLL�B.ZI_��@:�\��\��Ɖ�aC?ollaboƏr�
PANEL1�O� ��s	�C��qiPe�ndant Pa'nelJ��	9�:�"�5���R�d����2?�(�3��ԟ�{���2ß������X�j����3G�0�3��ܯ���3˯������`�r���4O�8�3� &�����φ�4ӿ�������h�z��vtTP�EINS.XML��=�:\)��ϥqC�ustom To�olbarj��yPASSWORD���FRS7���n��Passwor�d Config �ߥ7���0�m����  ����V���z��!� ��E���i���
���.� ��R���������A S��w��<� `���+�O� H��8��n /�'/9/�]/��/ /"/�/F/�/j/�/? �/5?�/Y?k?�/�?? �?�?T?�?x?O�?�? CO�?gO�?`O�O,O�O PO�O�O�O_�O?_Q_ �Ou__�_(_:_�_^_ �_�_�_)o�_Mo�_qo �oo�o6o�o�olo �o%�o�o[�o x�D�h��� 3��W�i������� @�R��v�����A� Џe�􏉟��*���N� ��������=�̟ޟ s����&���ͯ\�� ���'���K�گo��� ���4�ɿX�j������$FILE_D�GBCK 1z������� < �)
�SUMMARY.sDG	���MD:=��}���Diag� Summary�~��CONSLO�Gs�V�h���ߐ���sole lo�	TPACC�N��\�%D߁ߌ��TP Accou�ntin#ߋ�F�R6:IPKDM�P.ZIP�߹�
����ŝ�Exception
��i��MEMCHECK�w���lύ��Me�mory Dat�a���:n )x�RIPE��f�x�����%�� Packet L"ߞ�L�$�K���S�TAT��� ���� %)�Sta�tus��F�	FTAP����|�������mment TB�DF� >I)ETHERNE_����L�]���Et�hern2��fi�gura)DCSVRF������  verify all"��(4�DIFF��#�9diff�ZL�� CHG01���`)/��Q/\2��2///�/�N/`/��3�/�/�/1? ��/X?�&VTR�NDIAG.LS�]?? ?�?��u1 �Ope�4� ��n�ostic��'�)VDEVy2DAT�?�?�?�?���Vis�1Dev�ice�?�;IMG@y2��O&O�O"�QD�Imag]O�;U�P@ESO�OFORS:\_B]���Updates OListB_���@�FLEXEVEN���O�O�_���Q ?UIF Ev55���-vZ)
P�SRBWLD.C	M�_��-R	oD_��PS_ROBOW�EL;�:GIG���o�_�o��Gi�gE�H�_�N�@��)�aHADO�W�o�o�oO��S�hadow Ch�ange����.d�trRCMERR�G,>����pC�FG Error�W@tailv M�A�S�CMSGLIB���Y��b����bPic ��7�)E�ZD�o���B�׏��ZD�`a�dy�� rNO�TI���ȏ]���Notific����,�AG)�CRSENSPK�O����\���� �CR_ؑOR_PEAK柍�.�@�� d�翈������M�� q�����<�˯`�� ���%���̿���� ϣ�%�J�ٿn����� ��3���W���{ύ�"� ��F�X��|�ߠ�/� ����e��߉��0�� T���x����=��� ������,���=�b� ��������K���o� ����:��^p+ �#�G��} �6H�l�� 1�U��� /� D/�U/z/	/�/-/�/ �/c/�/�/?�/�/R? �/v?�?C?�?;?�?_? �?O�?*O�?NO`O�? �OO�O7OIO�OmO_ _�O8_�O\_�Om_�_ !_�_E_�_�_{_o�_ 4o�_�_jo�_�o�o[o �oSo�owo�o�oB �ofx�+�O a���,��P�� t������9�Ώ]�� ���(���L�ۏ폂� �����s�ܟk� ��� �6�şZ��~�������C�دg�y�����$FILE_FR�SPRT  ���������'�MDONL�Y 1z;��� 
 ���~�˯�� ﯯ�ؿ������ �2� ��V��zό�ϰ�?� ����u�
ߙ�.߽�;� d��ψ�߬߾�M��� q����<���`�r� ��%��I������ ���8�J���n���� ��3���W�������"���F��S|%�VI�SBCKY�C�h��*.VD��; �FR:\� ION?\DATA\�^�; Visio�n VD file�ASiwa �*��`��/ +/�O/�s///�/ 8/�/�/�/?�/'?�/ 8?]?�/�??�?�?F? �?j?�?�?�?5O�?YO kO&O�OO�OBO�O�O xO_�O1_C_�Og_�O��__,_�_!�LUI�_CONFIG �{;���[ $ �S^��V#o�5oGoYoko}o�i`|x�_�o�o�o�o�o| �o0BTfx� �������,� >�P�b�t�������� Ώ��򏉏�(�:�L� ^�p��������ʟܟ ��$�6�H�Z�l� �������Ưدꯁ� � �2�D�V�h����� ����¿Կk��
�� .�@�R��vψϚϬ� ����g�����*�<� N���r߄ߖߨߺ��� c�����&�8�J��� n�������_��� ���"�4�F���j�|� ��������[����� 0��Afx�� �E���, �Pbt���A ���//(/�L/ ^/p/�/�/�/=/�/�/ �/ ??$?�/H?Z?l? ~?�?�?9?�?�?�?�? O O�?DOVOhOzO�O #O�O�O�O�O�O
_�O ._@_R_d_v_�__�_ �_�_�_�_o�_*o<o No`oro�oo�o�o�o �o�o�o&8J\ n���������tRobot� Speed 100%�:�L�^�p�|���r  x������$FLUI_�DATA |����Ł��q��RESUL�T 3}Ņ�� �T�/w�izard/gu�ided/ste�ps/Expert��%�7�I�[�m���������ǟٟ���Continue with G�ance�"�4�F� X�j�|�������į֯6� ��-��Ņ>�0 ��p��ǃƁ'����ps �r���������̿޿ ���&�8����_� qσϕϧϹ������� ��%�7ߏuт�q'���+�=�+M�cll�b�ToolSe�t��g/Dist�Work@����� ��%�7�I�[�m���.0������� ������%�7�I�[�m�����w{ݐqo�t��?�&M�rip����Num/NewFram�+=O as��������0x��
. @Rdv�������p��c�/���E�M���imeUS/DST�y/�/ �/�/�/�/�/�/	??�-?�Enabl a?s?�?�?�?�?�?@�?�?OO'O9O����/sO5/G/Y&24d/�O�O�O�O_#_ 5_G_Y_k_}_<?N?�_ �_�_�_�_oo1oCo Uogoyo�oJO\OnO�O�B���
�ditor �o/ASew������� To�uch Pane�l s (rec_ommen�)� $�6�H�Z�l�~�����0��Ə؏� ��o�o���o�oracces`�p���������ʟ�ܟ� ��$�?�C�onnect t?o Netw��g� y���������ӯ���	��-�싘O����#���!E�pInt�roduction6�˿ݿ���%� 7�I�[�m���u��� ����������
��.� @�R�d�v߈����]�`�߁���Us�_ #�5�G�Y�k�}���0�������q1��� �%�7�I�[�m���� ���������a
��ѐ��������)����A��ve���{�� �������
0xFE/^p ������� //$/2*�c.L/� 2D/Macr}o�s/New�" _��/�/�/??(?:?�L?^?p?�?�0x0�?�?�?�?�?�?O O)O;OMO_OqO�OB&0��]/�O�/�,�/�+�"Open�#_5_ G_Y_k_}_�_�_�_�_ �?���_oo1oCoUo goyo�o�o�o�o�o������O�O��-�O�OoClos�w�� ��������_2+�Q�c�u����� ����Ϗ����)�@�o�iR���=���SetMethod.���ӟ���	���-�?�Q�c�u�8��c�[������W�n��?�ړ������ ̯ޯ���&�8�J�\�n��� ="iqr��Oa�s���$����t�raightOffset���,�>� P�b�tφϘϪϼ����=�X�g����g������,�>� P�b�t߆ߘߪ߼����l�����ѿ�%�S�M�X��o�� �������������#�>.0<�'�Q� c�u����������������)A��h  ��+�=�O�Y*� ���/AS ew6������ �//+/=/O/a/s/�2DV�/z��tZ~/?)?;?M?_?q?��?�?�?�?�?�1?17.762��? OO1OCOUOgOyO�O��O�O�O�/�/�$B�#�%�/�/׺)�/���RotationIWW�Oo_�_�_�_�_��_�_�_�_o�?180�Ko]ooo�o�o �o�o�o�o�o�o#�OXC3�_%_7_I_onP&��� ���/�A�S�e�$o �������я���� �+�=�O�a�s�2�/`�/hz��nRz� �)�;�M�_�q�����8����x�-99o� ��(�:�L�^�p����������ʿ����´ȩ����,"ݟ�tp�3Zdir/Tp3zοd�vψϚϬ� �����������?<� N�`�r߄ߖߨߺ��� ������ӿ��O���� +1��Mea�surement�/Straigh ?����������+� =�O�a� �2ߗ����� ������'9K ]o.�@�R�d�v���/We��Nums//New�sv '9K]o����v�0x��� / /$/6/H/Z/l/~/�/�/�/�/-`��)��#�.��Tool�Use�/l?~? �?�?�?�?�?�?�?O)j1OAOSOeOwO �O�O�O�O�O�O�O_$_-a
�/���/Y_x?-?�PartR? �_�_�_�_�_o#o5oGoYoko*B2oo�o�o �o�o�o�o%7 I[m,_��K_�r�(�_�s/G�� �r� �2�D�V�h�`z��������� �����0�B�T�f� x�����������{}�ȣ�#�)��yPa�yload1Cm �b�t���������ί�������p��[�c�Ȃ��c-���L�^�p� ��������ʿܿ� ��}�ٟ�/5��� 3��Y϶�����������"�4�F�X�j��10׏�ߤ߶����� �����"�4�F�X�j�՟W�A ��[���=�2O���,�>�P��b�t���������'��ێ�5��� $ 6HZl~���@υ�C����}P&�����Advanced�\n���������/{�0x��:/L/^/p/�/�/ �/�/�/�/�/ ??u�A��1?u�%%���Mass/Center�1?�?�? �?�?�?	OO-O?OQO cOҏ�O�O�O�O�O�O �O__)_;_M___v��0?�_f?��?ss ��j_oo+o=oOoao so�o�o�ohOzO�o�o '9K]o� ���v_�_�_�_�[),�_��G.c�2�XX�^�p��������� ʏ܏� ��o�o6�H� Z�l�~�������Ɵ؟ ���������'�9�sY���į֯ �����0�B�T�� %���������ҿ��� ��,�>�P�b�!�3�`E�W�i�{���sZf� ��*�<�N�`�r߄� �ߨ�g�y������� &�8�J�\�n����@��uχϙϫ�.����p�P�\L�[�m�� ���������������� ��3EWi{�� ���������`�� ��$�6�rt�� �����	//-/ ?/Q/"�/�/�/�/ �/�/�/??)?;?M? _?0BTfx�rt��OO'O9OKO ]OoO�O�O�Od/v/�O �O�O_#_5_G_Y_k_ }_�_�_�_r?�?�?�?����<TCPVer�ify/2cMethod�_Vohozo�o��o�o�o�o�o�o�L�Direct Entry8J\ n���������H�_'��_�_j'o+ofyJ����� ȏڏ����"�4�F� X��O|�������ğ֟ �����0�B�T��_�A��_��[�m��fy ���
��.�@�R�d� v�������k�п��� ��*�<�N�`�rτ� �Ϩ�g������ϯ���ӯfy�?L�^�p߂� �ߦ߸������� ￰�117.762 ǿ/�A�S�e�w��� ��������������B�%������/mW��������������1CU�80ÿ����� ��!3EW�D�C39�G�Y�k�}�PZ�//+/=/O/ a/s/�/�/�/���/�/ �/??'?9?K?]?o? �?�?�?d���Ϛ���yR�?IO[OmO O�O�O�O�O�O�O�O�-9m&_8_J_\_ n_�_�_�_�_�_�_�_�_�?�9´�?�?L�*O#OfyMeano�o�o�o�o�o�o 0B_*gtS �������� �"�4�F�oou�3o�EoJ)eowo�`ax V����)�;�M�_� q�����Tf˟ݟ� ��%�7�I�[�m�������b�������K"���ˁIntroductio�o?�Q� c�u���������Ͽ� �%�2�$�6�H�Z� l�~ϐϢϴ��������ϵ ��ѯ���B�ˀ ߇ߙ߽߫� ��������)�;�M� �q��������� ����%�7�I��6��,�>� M#a�fil�e2/cycle�powƆmode T�����1CU�gy���#�z��b�g�X�^�[�g���� 0BTfx����&e�!� Џ�����La�ui�dedȄSafety�5/G/Y/k/}/ �/�/�/�/�/�/T�? ?1?C?U?g?y?�?�?@�?�?�?�?�?g�g���O�����/don���O�O�O�O�O�O �O_ _2_D_?h_z_ �_�_�_�_�_�_�_
o o.o@o�?O#OmoGO/ȄReg,��o�o �o"4FXj|����Europ O�����#�5�@G�Y�k�}�����abAzc�o}o�oML�o� Timez}@EU��5�G�Y�k�}��������şן韨wE�ET Ea rn �sa�o+�=�O�a� s���������ͯ߯�
���c`�ߏя㏡o��24�������� ��Ϳ߿���'�9� P_]�oρϓϥϷ��� �������#�5�G�^o��*�<�RO`�24/currentL� ������)�;�M�_��q���s29-�NOV-25 17:29 ������ ����*�<�N�`�r�����_����yߋ��� �߿�Year ��2DVhz�������v2025�*<N` r�������� 
����  ����-/��!��Month��/�/�/�/ �/�/�/??)?;?�u11C?j?|?�?�? �?�?�?�?�?OO0OBO/' /�O�U/��DayFO�O�O �O_!_3_E_W_i_{_�_L829�_�_�_�_ �_oo*o<oNo`oro�o�oUOgHsO�o���O��Hou -? Qcu������L97��$�6�H� Z�l�~�������Ə؏�ꏩogH�o)���"|�og(inute� ��������̟ޟ�� �&�8��_\�n����� ����ȯگ����"��4����o-�;�Q �Q���NetDon r�ѿ�����+�=� O�a�sυ��nA�ϻ� ��������'�9�K� ]�o߁ߓ�W�W��� �ߍ�O"��	��-�?� Q�c�u������� �����)�;�M�_� q�������������I����߽�����X j|������ �0��Tfx �������/ /,/����!3E �/�/�/�/�/??(? :?L?^?p?�?A�?�? �?�?�? OO$O6OHO ZOlO~O�OO/a/s/�/ �/�O_ _2_D_V_h_ z_�_�_�_�_�_�?�_ 
oo.o@oRodovo�o �o�o�o�o�o�O�O�O��O��W�Summary�ov���� �����*��_N� `�r���������̏ޏ ����&�8���	�-?��RobotOp<�ʟܟ� �� $�6�H�Z�l�~�=��� ��Ưد���� �2�@D�V�h�z���O�O��a�������&��cl�lbWtToolS�etting�Off��(�:�L�^�pπ�ϔϦϸ����ϛ�1����)�;�M�_� q߃ߕߧ߹����ߣ��
�iͷK���%��n��{���� ����������/���23�Y�k�}������� ��������1�ߢ��q��.E�/��SpeedLimit/Max� 6��� 2D�Vhz��	1000.�0���� ��/!/3/E/W/i/�{/�+IsDz � gy����Val�/,?>?P?b?t? �?�?�?�?�?��O O(O:OLO^OpO�O�O �O�O�O�O�/�/�/�/����//Introductioi� p_�_�_�_�_�_�_�_  oo$o��HoZolo~o �o�o�o�o�o�o�o� 2M���M'_���A_� lectWork4�������/�A�S�e�w�6iLightwe��} �qpiece�� ��Ϗ����)�;�pM�_�q���  ErA�Sew�4��/Load�No�tHW_l��W�W ����.�@�R�d�v����������Я;d.3 �?���"�4�F�X�j� |�������Ŀֿ�OÙ�>�����ɟ7�8�����CenterMassڿ�Ϙ� �ϼ���������(� ��?Q�c�u߇ߙ߫� ����������)�� �C���3Z5=�O�a�omml�.����� ����1�C�U�g�y��<cEOAT w?/o par��� ��������
.@Rdv;xA﫟� w��/����+= Oas����� 8��//'/9/K/]/ o/�/�/�/�/�/4�8X����2�� g�n?�?�?�?�?�?�? �?�?O"O�FOXOjO |O�O�O�O�O�O�O�O�__�/�/?c_%?�/9?K?���_�_�_�_ 
oo.o@oRodovo�� �_�o�o�o�o�o *<N`r�C_��y_�+�_��� "�4�F�X�j�|�����8��ď�h10;O�� ��,�>�P�b�t����������Ο9_�yA  Y_�}_��~a?k�}� ������ůׯ���� �6OC�U�g�y����� ����ӿ���	��ڟ�V_`�"�,5�G��_ ����������*�<��N�`�r߉b�cith�o�߷��������� �#�5�G�Y�k�<�P���r��6��/� �ContactS�topInvalidArea/�PlusZz�$�6� H�Z�l�~��������� ݏ���� 2DV hz����-ϓ������7�����Min�v��� ����//��</ N/`/r/�/�/�/�/�/ �/�/??������51C�XY	�XY"?�?�?�?O O%O7OIO[OmO,/�O �O�O�O�O�O�O_!_ 3_E_W_i_(?:?L?^?�p?��)�?��NotHW_l�o!o 3oEoWoio{o�o�o�o �o�AR��o�o& 8J\n������P�_����_���_U����\�n��� ������ȏڏ���� �o4�F�X�j�|����� ��ğ֟��������9���� -��1S�peedLimi o��ïկ����� /�A�S�e�$������� ��ѿ�����+�=� O�a�s�2�D���h��Sy����Modet� ��)�;�M�_�q߃��ߧ߹�|GDo �not Use �(Recommended)�� �� $�6�H�Z�l�~���T������"���� �ϳ��\��9�K�]�o� ���������������� |�5GYk}� ������yH�����7�#�� ������// */</N/`/�/�/�/ �/�/�/�/??&?8? J?\?-?Qcu �?�?�?O"O4OFOXO jO|O�O�O�Oq/�O�O �O__0_B_T_f_x_ �_�_�_�_?�?�?�? �?,o>oPoboto�o�o �o�o�o�o�o�O( :L^p���� ��� ���_�_�_ oo~�������Ə؏ ���� �2�D�V� g�������ԟ��� 
��.�@�R�d�#��� G�Y�k�Я����� *�<�N�`�r������� ��˯޿���&�8� J�\�nπϒϤ϶�u� �ϙ�����"�4�F�X� j�|ߎߠ߲������� ���˿0�B�T�f�x� ������������� ��)���M������� ����������( :L^���� ��� $6H Z�{=��a�u� ��/ /2/D/V/h/ z/�/�/�/o�/�/�/ 
??.?@?R?d?v?�? �?�?k���?���/wizard�/cllb/st�eps/Summary�?HOZOlO~O �O�O�O�O�O�O�O�/  _2_D_V_h_z_�_�_��_�_�_�_�_
o�2��7�?�?�?�(O/�Configur�ationCompleteo�o�o �o�o�o(:L ^_������ � ��$�6�H�Z��6A#o5o�Yo�3qo�/SignalN�umberAss�ـment/SPIރd�	��-�?�Q��c�u�������ju1 ��ٟ����!�3�E��W�i�{��������1
@�9��a���2ŏ׏�D�U�g�y��� ������ӿ������ -�?�Q�c�uχϙϫ� ���������į֯�����
ߐߢߴ� ��������� �2�D� V�mz�������� ����
��.�@�R��:߉�{�U������ ��&8J\n ���c����� "4FXj|���?�?������� /./@/R/d/v/�/�/ �/�/�/�/�/�?*? <?N?`?r?�?�?�?�? �?�?�?O���GO 	/nO�O�O�O�O�O�O �O�O_"_4_F_?W_ |_�_�_�_�_�_�_�_ oo0oBoToOuo7O �o[O�o�o�o�o ,>Pbt��� �o�����(�:� L�^�p�������eoǏ �o돭o�$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ����� �ۏ=����v����� ����п�����*� <�N��rτϖϨϺ� ��������&�8�J� 	�k�-��ߡ�e����� �����"�4�F�X�j� |���_��������� ��0�B�T�f�x��� ��[ߥ�������� ,>Pbt��� ������(: L^p����� ��������/E/ l/~/�/�/�/�/�/�/ �/? ?2?D?h?z? �?�?�?�?�?�?�?
O O.O@O�/#/5/�O Y/�O�O�O�O__*_ <_N_`_r_�_�_U?�_ �_�_�_oo&o8oJo \ono�o�o�ocOuO�O �o�O"4FXj |�������_ ��0�B�T�f�x��� ������ҏ����o�o �o;��ob�t������� ��Ο�����(�:� �K�p���������ʯ ܯ� ��$�6�H�� i�+���O���ƿؿ� ��� �2�D�V�h�z� �Ϟϯ���������
� �.�@�R�d�v߈ߚ� Y���}��ߡ���*� <�N�`�r����� ��������&�8�J� \�n������������� ������1����j |������� 0B�fx� ������// ,/>/��_/!�/�/Y �/�/�/�/??(?:? L?^?p?�?�?S�?�? �?�? OO$O6OHOZO lO~O�OO/�/s/�O�O �/_ _2_D_V_h_z_ �_�_�_�_�_�_�?
o o.o@oRodovo�o�o �o�o�o�o�O�O�O 9�O`r���� �����&�8��_ \�n���������ȏڏ ����"�4��o )��M��ğ֟��� ��0�B�T�f�x��� I�����ү����� ,�>�P�b�t�����W� i�{�ݿ����(�:� L�^�pςϔϦϸ��� �ϛ� ��$�6�H�Z� l�~ߐߢߴ������� ����Ϳ/��V�h�z� ������������
� �.���?�d�v����� ����������* <��]�C�� ���&8J \n������ ��/"/4/F/X/j/�|/�/M�/q�/�+��$FMR2_GR�P 1~�%�� �C4�  B�� 	 � !?3<0F@� I?@�+0G� � q1Fg�fC��8R}5a=?�  x�?�,06�X��2��875t��5���5`+�a=�A�  �?�;BHx�4_0E@S33!EB�,4COTM0@A jO`>TO�O�O�O�O�O �O_�O2__/_h_S_��_�#�"_CFG ;T32�_�_�_|�_�YNO :/
F0.a 3`�\�RM_CHKTYP  �!� 00�� �!ROMI`_MsINO`�#��{`u�:@X� SSB�S���% 6�o�%�c�o�o�U�TP_DEF_O/W  �$3�g�IRCOMN` ��$GENOVRD�_DOpf�-}TYH�0rd dJud3to_ENB 3p�RAVC�#��g�` �A5�o�y_��a<��1J ��qOU 0�<�6a18r15< x`�?��/�}���͏�#C��3�!���o"�^�!>����Br0��49p��o�pSM�T�#��y0�`���$HOSTC�R19�9�`���0� MC�$
��ȟ�&  27.�0�1�  e ��E�W�i�{��*3������Я������	a�nonymous@	�7�I�[�m�� ǟ0���������,� 	��-�?�QϘ�uχ� �ϫ�οh������ )�;߂��Ϧ������� �������Z�7� I�[�m��������� �������V�h�zߌ� ��{��ߟ��������� .�/ASv��� m�����*�<� N�+bO��s�� ������//8 ��]/o/�/�/�/� �"$/?X5?G? Y?k?}?��?�?�?�? �??B/T/1OCOUOgO yO�/�/�/�O�?�O,? 	__-_?_O�Ou_�_ �_�_�O�_O�_oo )o;o�O�O�O�O�_�o �O�o�o�oZ_7 I[m�o�_�_������|���EN�T 1�P� P�!�V�  'p D���p���h�ɏ��� ����ԏ"�G�
�k�.� ��R���v�ן����� П1���U��y�<�N� ��r�ӯ�������ޯ �Q�@�u�8���\��� ��ɿ����ڿ;��� _�"σ�Fϧ�j�|��������%���QU�ICC02��!�192.168.O1.10K�@�1��^� ���D�2�߮����!�!ROUTER"���!r�I���?PCJOGr�M�_!* t�0{�~=�CAMPRT��ƞ�!r�����RT�;�����`� !S�oftware �Operator? Panel=�o�����NAME �!3�!ROBO����S_CFG �1�3� ��Auto-s�tartedidFTPtoI�o� t�o�����- (:]K�� ����Kn"4F #/Z|:/k/}/�/�/ h�/�/�/�/?0/�/ C?U?g?y?�?�?Rodo vo�o?	OP/-O?OQO cOuO<?�O�O�O�O�O O�O_)_;_M___q_ �?�?�?�_�O�_$Oo o%o7o�O[omoo�o �o�_Ho�o�o�o! 3z_�_�_�_�o��_ ������o/�A� S�e�w�������я ����N`rO��� s��������͟���� ��'�9�\�]�🁯 ������ɯ�"�4�F� H��|�Y�k�}����� h�ſ׿����0��� C�U�g�yϋϝ���� ����	�P�-�?�Q� c�u�<ϙ߽߫����� �߆��)�;�M�_������_ERR ����o��PDUSI�Z  �^�����>��WRD �?���  �guest ������%�7�I����SCD_GROUoP 3� �
�IFT��$P�A��OMP��� ��_SH��ED��� $C��COM���TTP_AUT�H 1��� <�!iPenda�nU�`'!K?AREL:*`i{KC���� �VISION SETy���'?:�^p���������/C�TRL ����I(�
�'F�FF9E3/���FRS:DEFA�ULTn,FA�NUC Web ?Server��\! L"/����,�/�/?�?,?>?}�WR_C�ONFIG �.~���cn/��IDL_CPU_kPC� �B����0 BH�5MIN��<��5GNR_I�O������0HM�I_EDIT ��~�
 ($I�PL_�"_SMP�LGR3 LOSE�Icon 2B��^OOPEN2Bt7H�51 FOXO2�2mOO$ bkt�lead-ins�t_basicp�ick_star ^I/�O�O__;_&_�__J_�_�_Z!($*uninit� t[�_�_�_o�_/oo ,or_wo�oto�o�o�o�o�o�o�?$IN�PT_SIM_D�O�6�:NSTA�L_SCRN�6 ��UzTPMODN�TOLkwT{�!RT�YJx�1Yv3 EN�Bkw��3OLN/K 1���������1�C�U�g��rM/ASTE�0�yH"��qSLAVE ݒ��H D�uSRAMCACHE��|��5O_CFGǏ��s߃UO�ۂC�MT�@� �2���Y�CLƏ��� _AS�G 1�s7��
 i�������ԟ� ��
��.�@�R�d�v�\q�_�NUM�����
ۂIPďևRTRY_CN(���gqG_UP�����q��� ۂ���</  0I$3��0@gr�?��� ���DmplGrp/�Sar�e_Config.stm�� ������ѿ�ր�� �#�5�G�Y��}Ϗ� �ϳ�����f����� 1�C�U����ϋߝ߯� ������t�	��-�?� Q�c��߇������ ��p���)�;�M�_� q� ������������� ~�%7I[m�� ������� !3EWi{
� �������// A/S/e/w/�//�/�/ �/�/�/?�/+?=?O? a?s?�??&?�?�?�? �?OO�?9OKO]OoO �O�O"O�O�O�O�O�O _�O�OG_Y_k_}_�_ �_0_�_�_�_�_oo �_CoUogoyo�o�o,o >o�o�o�o	-�o Qcu���:� ����)���_� q���������H�ݏ� ��%�7�Ə[�m�� ������D�V����� !�3�E�ԟi�{������ïR�K�_MEMBERS 2�"�w2� $"����^������RCA_AC�C 2���   [}�z�}ZT�6�)ps�  &T��T�g�x�r�|�n����� I�BUF0�01 2�V�= �x�u0  uW0x�����곩y����#��.�9�F�Q��\�i�tā�ČėĤİ�Ļ������j�����z��U����(��3��U@��L��W��d���o��z�ć�ċ`  `wX곫we"�q"�|� �� A�x�xR�"�)�x1�x9��xP�I�xQ�xsJ관괋�q�xy�+x�괺���ǹ2Կ��������� �������� !��)��1��9�� A��I��Q��Y�� a��i��q��y�� ��������� ������걸��� ���������������� ���������������� н�	н�н���  ��(�-�1�-�9��� A�B�H���Q���Y��� 2�h���B�x���R�� �ґ��ҙ��ҡ���z� ���ҹ����������ǹ3���������� T����'�)� 7�9�G�I�W� Y�g�i�w�y� ���§��� ��T����������� ������������� �	����'�.)� 7�.9�G���#P�_� ��;h�w���y҇��� c�ӟ���ү�������������CFGw 2�V� 4�� ,T�T�<�!!]�HISѲ�V�� �g� 20�25-11-29�T� T�;  Gs#�/�/�/R�!XT� - h�$��v xr$z�{/�/?^=[|�pY(8e) ?^?p?�?�?�?�?�?��?�?T���� R��x�Y"1-07-06A?.O@OROdOR�^�s#�":�$ �$x�$�O�O�OT�/R�X�H5O
_x_._@_  T�#X��/p_�_�_�_�J▁H2�O�_�_�
oo.o@oRoP���x�O�oR�QgAY"0-08-31�_`�o�o�o�o
gAso�0BTf�boP�g2��o���E^���; -v fa#oP�&�8��Ӯ7&��C/U/g*bQd�y ��G���ɏ�*!d ��� 邚���� �� � ��"�4�"?4?�|� ������ğ֟���� �;�Oh�U�g�y����yH6  [� 8���`���� c �@邔�߯��O�OL��9�K�]�KZ8  ^]P}�h�������ѿ �_�_��+�=�O�a� s�ao���ϗo�o������'�x9  _0�[�m��m�����������	 U-�@ c�p��ɯ :�L�^�L�9$��h�z�g*�qy �������� �*��-��� �ⶠ�� � �����G�Y�G�Y� �ߡ����������� 1���2���z���yH��)��@6� ����lYk} k��]P����� ����,/>/P/b/t/ �/�/�ϩ�/����)/ ?(?:?L?x�/{?�? �?�?�߱��?�?OO �sra�6B�p6B�j?�_OqO�Oq�A_I_�CFG 2���� H
Cycl�e Timeq�Busyw�Idl�B�Dmi�n{QUp|�F�ARead�GDow�H�O���Q�CCount>�A	Num �B�C��{s]pKQY�P�ROG�B�������(/sof�tpart/ge�nlink?cu�rrent=me�nupage,1�53,�!s^�Uo��W631,�P l�e_Config.stm�Oo�MJU�y�SDT_ISO_LC  ���~���OJ23_DS�P_ENB  �^j��`INC �^kul`A   �?�  =����<#�
ka�i:�o �a�o�o��o�$xgOB�PC�c��E�f>qG_GRO�UP 1�^k>��< �tP�a(�	�,?��_� �!���(��L�^��p����6yG_IN_AUTOKt��i`POSRE�FXvKANJI_�MASK膯h��R�ELMON ���|_�yG�`�r���������N��S��W�Ճ�ʕ�քKCwL_L��NUM�`���$KEYLOGOGING�����*���e�PLANGUA_GE ��f���ENGLIgSH t�|�LG�A���ZR�'��  ��H � �� '�7  �W 
���� /o�=f ;��
�(?UT1:\��� ��'�9�P�]� o���������ɿ���(O���HQ�N_D?ISP ��o X���z�LOCTOLu��Dz�Pga�a���GBOOK ���-��Q��-��Ԫ������/��A�Qݑ�Sc�?�	���ԩ�q9j�߼�Q���_BUFF 2=�^k ��%�����>b��G �Collaborativ �%�7�� v����������� ��E�<�N�{�r���~��DCS ��Y �b�a`ܟ���E�'9��IO 2��� �@n�@�P�r������ �$6JZl ~��������/"/MER_ITM[nd��{/�/�/�/ �/�/�/�/??/?A? S?e?w?�?�?�?�?�?8�?��P"SEV��F�]L&TYP[nj/�KO]OoO�=�RST����SCRN_F�L 2�[�P� ���O�O__+_=_O_F�OTP3�[o:B�NGNAM�d��f��6�UPS_ACRx�@ꏾTDIGI�X�IU_LOAD�CpG %|Z%�HOME\_^_MA?XUALRM��Q���e
Bb�Q_�P�U�P ��a�B`CA���͜o�������ddpP 2��� �=�	:O�o+ OaD�p�� �����'�9�� ]�H���d�v�����ۏ Ə����5� �Y�<� N���z�����ן�̟ ���1��&�g�R��� v��������Я	�� ��?�*�c�N�����|� �����Ŀֿ��;� &�_�q�TϕπϹϜ� ���������7�I�,��m�Xߑ�:hDBGDEF ��e��o���_LDXDIS�A�P{[KMEMO�_AP�PE ?|[
 ��z�� -�?�Q�c�u���B`�FRQ_CFG k��g��A z��@���|�<��d%��������b��k{��*Q�=/S� **:\�|� O�a���|և������� ������2~ߍe[�2 L�p��,( 0�C��( 9^E�i������ //�6/8jI�SC 1�|YB� ���~/���ߔ/��/�/�/B/T"_MST�R �M5SC/D 1�
��/c? �/�?r?�?�?�?�?�? O�?)OOMO8OqO\O �O�O�O�O�O�O�O_ �O7_"_4_m_X_�_|_ �_�_�_�_�_o�_3o oWoBo{ofo�o�o�o �o�o�o�oA, Qwb����� ����=�(�a�L� ��p�������ߏʏ���'��K�6�o�?M�K���#=�ၟ$�MLTARM��u����� ������METP�U��b���+9N�DSP_ADCO�L����CMNT6.� !�FNJ�N�>�FSTLIo�`�0 �#>®����گ�!�POSCFz��Y�PRPMM����ST,�1�#;; 4��#�
^�j� ^�n�|�Z�|�~���ҿ ��ƿ����>� �2� t�V�hϪόϞ������!�SING_CH�K  r�$MODA���\+����~�DEV 	���	MC:N�HS�IZE��b���T�ASK %��%�$1234567�89 �����TR�IG 1�#; l�����		�J�F��YP�ѣ0���EM_INF 1��6�`)AT&FV0E0O����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ����H�F���:�n���Av���Y��������� �������� �w*�������� ��+O �8J\���/ :'/��]//�/h/ �/�/j�/���� 5?�Y?�/j?�?B/�? n?�?�?�?O�/�/CO �/??�O�OP?�O�? �O�O�?_�O?_&_c_ u_(O�_LO^OpO�O�_ �Oo)o`_Mo _qo,o��o�o�o�oG�NIT�OR��G ?b� �  	EXESC1f�r2x3xE4x5x��v7x8x9f�r�Ryt rytryt+ryt7ryt CrytOryt[rytgrytTsrys2�x2�x2�xU2�x2�x2�x2�xU2�x2�x2�x3�x�3�x3r�R_G�RP_SV 1��� (j�����b��w���o�ƥ�_Djb��ԃIO/N_DB$й(�b�_  �ސ�ސ)�A���`@����  
lF�m�A��`N   4�Z�&��=�-ud1tՊ����� ��PG_JOG ����ƫ
ˠ2���:�o��=���?�ˠ����*�ܞD�V�ˡm���n�00�'�ˠ+�@������ѯ�  �ѧ��L_NAME �!�� ��!�Default �Personal�ity (fro�m FD)Y��R�MK_ENONL�Y�G�R2�� 1��L�XLy� �O�l dm� ������ѿ����� +�=�O�a�sυϗϩ� ��������ߥ��$� 6�H�Z�l�~ߐߢߴ����� "���� #�5�G�Y�k�}��� ������������1� C�U�g�y��������� ������	-?Q cu������ �);M_q �������//��<��;/M/_/q/ �/�/�/�/�/�/�/?���E�a�� */ݟ*?_?��PN?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�Oh? z?�O�O�O__)_;_ M___q_�_�_�_�_�_ �_�O�Oo%o7oIo[o moo�o�o�o�o�o�o��o!o�ots����bt{x�d��8�� �{���w��G{���pN�A�7� .� Y�O�a�s�������׏�-�Ӑ��
���	�`C�=�O�a� �3�A�D�������[� A��̙(��q�q��"����tS|�_�  �tp�p�E�C{  ��&�G�"�k�V�{������ů�x�qH�j�p�����p+�� �� ��� @oD�  )�?�/���?Ā1�ā@I��)���˯  ;��	lA�	 ��X  �����y� �, � ��������K�oȩ���]�K��K]�/K	�.��_�Zx�����@
���J��Կ��T;f��I��Y�,�A�{S�ٽ�>  �3���Ck��j�#3��?2}H����bā��|S-��Ͽ�B���ᗸX�畨� D	�����g  �  �!ֵ�?���	'� � �]�I� � � �ٕ�:������È=�����-�@�߯�ھ���G��-���yN}�+�  'A���B�I��@�p��Q�V�Cj�Cn�C��� y�~�J1��|���܀ �{ Nſ A 0ݹB}���|��弝���āDz��$���H�3��X�~�i���������А #4P���ąz���r�б�p��?��ff������� �&8j�8ĀN\
C>L����=�ݺ(Ā�P�������q��� xi�;e�m���KZ;�=g�;�4�<<�0���/���y�ɐ?fff?��?y&;�@=0M?��YH�|�6 B�ݹ1��/��u� ��	/�-//Q/�</u/�/r/�/J�zF}��/�/�/?�,? ��/_?�/�?n?�?�? �?�?�?O�?%OOIO 4OmOXO�˜O��X�? �OB?_�O_A_S_e_ z_�_&_�_�_�_�_�_o����3dՙG��Cojoo�o����ؘo�o�o�oH��"{�k�}��dD
p,��L�d��`�aUqI���!n,ȴA2=q�@��T@|j@$�?�V�^��z�Ð���=#�
>\)�?��
=�G��}�{=r ��,��C+��B�p���p}B6���C7n����?6`��(���5}G�p��Gj��F�}��G�>.E�V�D�K�����I2`�F�W��E��'E����D��;�����I+aE����G��cE�vmD�����9 ��ď���ӏ���0� �@�f�Q���u����� ҟ������,��P� ;�t�_�������ί�� �ݯ��:�%�^�I� [��������ܿǿ � ��6�!�Z�E�~�i� �ύ��ϱ������� � �D�/�h�S�xߞ߉� �߭�����
���.�� +�d�O��s�����л�����p(�q343�]����9���x!�7��U3~�mU�g�I�5Q����I�Ǔ������Q��������=+(aO�EP�P��A�O���������#\ Gl�}���� ��"//��O�OL/�/p(��/�/�/�/ �/�/�/??C?1?g?�U?w?�?�P2/�? � B�;`p�1CHpz;`�P@BoOO@+O=OOOaOrM�C�?��O�O�O�O�O�S?���C�  @�S$�P�P�aS�4�U
 �ON_`_r_�_ �_�_�_�_�_�_oop&o8o�z(Q ��}���'x#�$MR�_CABLE 2��} ��tT� �f���o�	�o wI�`q�c�ow}� 7]1g��y ������3�Y� �-�c�����u����� 珽�Ϗ��/�U���k�1{B��o����˟������������*A�** qcOM� �~i��^�6 *[�|��+%% 2345?678901~���! {�����{@�{@�15{@{A
���m�not segnt J�ӣW��TESTFE�CSALGR  eg{J�1dC�QڡY
S�� � {D�Xbp�n������� 9�UD1:\ma�intenanc?es.xml����  +Z�D?EFAULTvLqb�GRP 2�b� � �{@}6*[�V{F  �%!1�st clean�ing of c�ont. v�i�lation 56��ڏ�	P����}5+*�}J���������X�%i�mec�hp�cal ch�eck�  �BS��@]�d�}5�π�ߣߵ����(�y�roller;�M�_�����U�g�y�����(�Basic �quarterl!y���$��,D��`#�5�G�Y� �M2���{@"8��N�N���}5�����b��t�C��O��s���������&(�Overhau��6|�' x{@18}5�ew���{@$V����wI T)/;/M/_/q/��/ ��/�/�/??%? 7?�/[?�/�/�/�?�? �?�?�?:?�?!Op?O �?iO{O�O�O�O O�O �O6O_ZO/_A_S_e_ w_�O�_�O�O�_ _�_ oo+o=o�_ao�_�_ �o�_�o�o�o�oRo 'vo�o]�o��� ���<N#�r G�Y�k�}������� ��8���1�C�U� ��y�ȏڏ쏢�ӟ� ��	��j�?������� ��������ϯ���� T���x�M�_�q����� 䯹�˿��>��%� 7�I�[Ϫ��ο࿵� ��������!�p�E� �Ϧ�{��ϟ߱����� ��6��Z�l�A��e� w�������� �2� �V�+�=�O�a�s��� ����������� '9��]������� �����N#r ��k}��� j�8�\1/C/U/ g/y/��/�/��/"/ �/	??-???�/c?�/ �/�?�/�?�?�?�?O T?)Ox?�?_O�?�O�O�O�O�O@JnB	 X`�O__(_lIB IO W_UOWE__�_�_e_w_ �_�_o�_�_7oIo[o o+o�o�o�oso�o�o �o�o�oEWi'�9������|� �wA?�  @nA 5_0�B�T��nF�������lH�*ŏ** F�@ �q�vp�����!���E�W�i�{��� zOFFߏ��ϟ�󟵟 �)�;�M�������� �����������Y� k�}��m����S��� ǿٿ�1�C���3�E� W�i�+ύϟϱ������WDnA�$MR_HIST 2��u}�� 
 \B�$ 2345678901�#��Ͽ��9Ozߌ�C�u� O�����߯���.�@� R�	��i���c��� �������*���N�`� ���;�����q����� ��8��\n%��nD��SKCFM�AP  �u��q���n@���ONREL � nD�����E�XCFENB�
8��FNC�JOGOVLIM��d�^�KEY��aj_PA�N�|x�RUN�Qa	�SFSPDTYP5 ��SIGN�T1�MOTS�_�CE_GRP 1��u���@r� _/nCL/�/�s/�/k/ �/�/�/?�/?D?�/ h??a?�?U?�?�?�? �?�?O.OORO	O\O �OoO�OcO�O�O�O_��K�QZ_EDI�T���TCOM_CFG 1͹ae_w_�_ 
FQ�SI �6+����_�_��_o����O@oXT_A�RC_�@T�_MN_MODE���=Z_SPL�co#UAP_CP�L�o$NOCHE�CK ?� � �o/ ASew����������NO_?WAIT_L�;W6& NTNQϹ�Ez�Y�_ERR0!2й	����'���Ə؏��_�/�~`�O��ю�|}�Z/oW��<���?���v�\�� I���P�ARAM��ҹ���G�������(� = V�E�W�_� 9�����o���ɯۯ��0������C�U���y��cUM_RSPACE�i��Q������$ODRDS�P�c� OFFS?ET_CAR1P�o��DIS���S_�A~`ARK�<YO�PEN_FILE����Q<VαPTION_IOr�s��M_PRG %���%$*�Ͼ�O�WmO;��6'��Ar����:!5�� '� ��	�j�	�G	 ��	��&���ϰRG_DS�BL  �� �r�v��RIENTkTO� �C�� ��A �U�`IM�_D{����ϰV~ӰLCT �c��8RҼ��d����_�PEX�`��RA-T�g d ����UP ���b��; �{��s����/$PAL]��c���_POS_CH<��&���Ő2/#�L��XL���l�j�D�V�h�z� ��������������
 .@Rdv����22�����#5GYk}� ������// %/7/I/[/m//�/�/ �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_k���_�_ oo+o=oOoaoso�o��o�o��E�a :Ҭ��o�����o	:�P�o3EWi{� �������� /�A�"w������� ��я�����+�=� O�a�s���T�f���͟ ߟ���'�9�K�]��o���������ɯۮ���;����j�dg�8�J�/�m�{���e�������进� 8�׷���	��9�?π]�����ϲ�:�ֵ	`�����	���:�o��'�9�K�|]�f�A�  t٨и_�_��"��x������  ����#���C{  ο ��ʿ���#�I�4�m�`��_��Z��OU���/��/��H'���� ۷ ���� �@D�  ��?������?���៑C4�����s�  ;��	l��	 ��X  �/�4�%� �, � �E�J���Hʪ�U򏓤�H���Hw�z/H�P���x������B�  ������������>  ?�3���C������c��������B���������R��f�ek���������T Dڵ�����g  �  ���]����	'� �� 	I� ��  ��Ռ�=����-?��@U[�����[������N%�� � '���C C C�� �*��/�a�`�$�z��{ Nq� A 0��B%Ѕ%$ё%d�l�%��DzV��//�/�/�?*?���A2���I2А #4PI"Z5��z��^��|���l ?��ff���?�?/? ���?�;��8���?JC>LO~ ���(��6EP?HZ9<�3�7��C1 x��;e��m�B�KZ;�=�g;�4�<<a�m��O�?�����|%Bq�?fff?l�?&�@��@=0�E?��U�Y$� �A�����=_��\_�G !��?�_|_�_�_�_�_ �_�_!o3ooWoio@o �oxo�o(_J_L_�o �o/S>wbt �������� �H����o���o�� z��������O&�8� ҏk�V���z���ş��"�"�ߔ}��C���x��:�%�?��D��K���o����� %�~�D��د�^��^�]��@I��͞,ȴA2=q�@��T@|j@$�?�VT���z�Ð���=#�
>\)?��
=�GH����{=@��,��C+��B�p��[�B6���C7n����?���(���5G�p��Gj��F�}��G�>.E�V�D�K������I2`�F�W��E��'E����D��;������I+aE����G��cE�vmD�����:�� 7�p�[ϔ�ϸϣ��� �������6�!�Z�E� ~�iߢߍߟ������� �� ��D�/�T�z�e� ����������
��� �@�+�d�O���s��� ����������* N9r]o��� ����$J5 nY�}���� �/�4//X/C/|/�g/�/�/m�(m�343�]�/mA���%�%x�/�/U3~�m??�"�5Q-???�"Ǔ�Y?k?Q�����=�9�?�?�?�?(O�<n�P�BP?N^�[�hO�/tO�O�O�O�I�����O�O_ �O_>_)_b_M_�_q_ �_�_�_�_�FP�R��_.oh�1o;oqo_o �o�o�o�o�o�o�o�#Is02�_t � B�琾��qCH��z�s0@�@�����t�c�H�Z�l�~���s3?����=@ @s35ts0s08���[ts5
 ������0� B�T�f�x���������pҟ�c�ԁ ��);��'x#�$PA�RAM_MENU� ?�5��  DEFPULSE��	WAITTM�OUTH�RCV�[� SHEL�L_WRK.$CUR_STYLF�;��OPT�q���PTB����C��R?_DECSNS�0E �\���!�J�E�W�i� ��������ڿտ����"��SSREL_�ID  �5YA��1�USE_PRO/G %,�%σ�2�CCR_�C�YA4����_HOST �!,�!���ϐ�T P@���û�����0�>��_TIME]�C�����GDEBU�GA�,�2�GINP?_FLMSKY߈�sTR�߈�PGA��e x�7���CH��^��TYPE)�5���M�v�q��� ����������%� N�I�[�m��������� ��������&!3E ni{���������WORD ?�	,�
 	RyS���CPNS�E���:JOɡ�B�TE�DCOL��E����L_� ��0�s0ȫ�dm�T�RACECTL �1ׅ56� }=@ *=@�7@��DT Q�؅5 �D �� i� U' 	+$
+$+$Q+$�0-"+$+$TC�-"+$+$+$e+$+!/C�/ WA-"��-"Ѐ-"��-"Ȁ-"Ā-"+$*/</ N/`/r/�/�/�/�/�/ �/ ??$?6?H?Z?l? ~?�?�?�?�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�o&8J\n���#!�%k� }�������ŏ׏��� ��1�C�U�g�y��� ������ӟ���	�� -�?�Q�c�u������� ��ϯ����)�;� M�_�q���������˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���!�3�E�W�i�{� �ߟ߱���������� �/�A�S�e�w��� g������������!� 3�E�W�i�{������� ��������/A Sew����� ��+=Oa s������� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�? �?�?�?�?�?OO1O COUOgOyO�O�O�O�O �O���O	__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o %7I[m� �������!� 3�E�W�i�{������� ÏՏ�����/�A� S�e�w���������џ �����+�=�O�a� s���������ͯ߯������$PGT�RACELEN � �  �����3�_�UP ���e�b�j�N�c��3�_CFG ڦb�L��
c�����������E����  ���w�DEFSPD ۂ���E��3�H_�CONFIG ��b�J� �j�d)��B� ��,�PôƱH����3�INz�TRL �ނ���8õ]�P�E�����b���(���3�LID�{����	��LLB� 1�� 5�I�B8�B4Ӵ� I�!��LŶ� << �?�K�j�K�b߄߲� �ߺ����� ����@8�f�L�n���4� �������M���<�/��A�r���GRP 1������@A!����4I��A� �Cu�C�OCjVFx����-�Ʊ����(�(����q�C���#´B$BE l�L6H�l��?&�B34����`�j4M J�n��,�����%//  DzJ#S/��:/{/*/�/ �/�/�/�/�/�/?? A?,?>?w?b?�?�?�?��:)�1
V7.10beta1���+�@�*�@��) @�+A� )�?��
?fff>����1�B33Aж�0�
CB(��A���AK���9AD�	AVOhOzO�O�O��p2���8�@@>K���@A���?�ff�?�@�������Mb��� ����?��?�,_>_@(_b_L_�_�1)�l���u)A�Zb��_��_�o���1EE�A�S BfڰB�:o,eBHbc��T���MdI�Q��T��Q��Tx�dxo�o o�o�o�o l���2��-?s)W�M_	t���KNO?W_M  �������SV ��?�Y�i/�� ��_�D�/�A�z������M����� �B	~��6� I�^���Z���O
�b�T�@ڱ�1ڰ$�� �2����MR�����T�_^+�����~��OADBANFW�D���ST��1 �1�b��p4�EOAT w/o part��B�����=LQ�0�B��� f�x��������ү� )���,�>�P�b���@������ܿR��2����4ڿ  �</���3�+�=�Oς�4l�~ϐϢ��5 ���������6�$�6�H��7e�w߉ߛ߂�8���������M�AҐ����O�VLD  ��ޏz��PARNUM  ����#��n�SCH]� k��
�������UP�D���^��_C�MP_��`����p'�ޕv�ER_CHK����ޑǂ�������RSq�՟�q_�MOҟ��_��
�__RES_G���
ROʽ_d��� ����7*@[N`3�@P �5k����7�� ��/7�/</A/ 7d�\/{/�/7�Л/ �/�/7
��/�/�/7�V 1��fې���@`h���THR_INRq�bፂޕ�dm6MASSz? �Z�7MNy?�3MO�N_QUEUE ����ޖ �@ *
�N{�U��N�6�8��3ENDAIEcXE*OE@�BE)@|O�3OPTIOG�(�0PROGRAoM %�:%�0�8?���2TASK_�I_�qNOCFG ���?���OPDAkTA���[`a��2ƅu_�_�_�_�_ h_�_�_oo)o�_Mo�_oqo�o6_INFO
���S]��4?o�o�o  $6HZl~ ��������� �2�D��g�d�S\ �nQ��DIT ��_����TWE�RFLKH`3�CRG�ADJ �A	���? ��1���1
P�a���?���z��cQ<@	����f% �r�وn�!�MQ2�/��b	H��0lA7_2<�>������t$��*�/� **�:�� ������6�1����;��� a�C2[�)���9�K�y� o����������ۯ� g��#�Q�G�Y�ӿ}� ������ſ?����)� �1ϫ�U�gϕϋϝ� ��������	߃�-� ?�m�c�u��ߙ߫��� ����[���E�;�M� ��q�����3��� ����%���I�[��� ������������� w!3aWi�� ����O�9 /A�ew���X6	"_F/ۀ4/m/X$ 㙏/�[/�/W/�/�/����*SYST�EM�V9.40�107 27/2�3/2021 gA%݀
7��#��PREF_TLA( $GRID@�ES  $B�ARcB]2STYL�E]1��?0OTO�ENTJ0 � $P_NAM�s0!�0{2]1z1X�Y(�J1 � �$LIST_POsRT]2�3ENB�8�SRV�0)�4�6DIRECT_1�2��42�93�94�95*�96�97�98�1x1sF_HRK0  Q0_VALUEv�S0�OUPv�$AX�ISzAWC�4� !$ENABr0� �1G�3�%$CUR��wERcAN�C�Bn0AR�0�YPoA$TOTAL_TI�Ar@�C�PWRpBIC1�DR�EGEN�JRpBE3XE\A�A$]C�A�^1REe0�EMON�TR_R)Q�2�A_�Sx@WWP:SV_L�IM�0tV@�1EG�RE�CG0?PHzBO�VERU0�TV_H�d0DAYSV�QS�_Y�A$MAX�SIZ9SSUMM�AR�P2 $�CONFIG_S�ET�CUP�2{AL�A�0RUQ=QC_�o6$CMPR�4� cDEV�@�P/bI��@Z c�S]1XBE�NHANCE�A | 
�E*a�@TTN�QINT�0QM(�|^1��_MASKj3PD_OVRD�3�GE2IX�0JPAX�yPZ5OVCyQ�TB�UqRWCF5 4 �S?e71[o6�PS�LG�P�A \ �$PS_�V=pMO�P^1�AS�0ra3aU<q�fTv�SDbtAUx1-p80P�A (0Q�Ar�JvOPCrFI�L_McS�qVELL:S�0TQLP�3N�0�.PCPSUL�P _ 	$V�{C��P_�po@�M'�V�1&�V14�2C�2�4�3C�34�4C�44��A�0 ��@��ܿ0��MINщVI#B1+0��2�*1T����3��3��4��4���@�L��@@���@̇Ʌ݅ɅPLUS_TORQnAp؅����+pSAVba�	d $MC_FOLDER`	$SLđÑse��@M�pIsc��LO}A�`  $��2cΐKEEP_H�NADDّ!�R�#�CCOMi0`;�{1ڒ=p<�OP ��b�ؑ_0<�xg<�REMS�;��A�2x�ԏ���U�4e;�HP�WD  �S�BM�a�0COLLCABLt�@>p�AE�a��@ITSa��r�$NO�FCAL(c�CDONrb�qÒܚa�0
 ,Q0FL�ANGoA$SY�NҐI�M�0Cb�~�@UP_DLY�1=C�DELA{��A�k2YPAD�Q$TABTP_R���QSKIP:�g Ĵ0�PORk������P_�Pʰι �@J��b�}Q���Q�� @��@��+@��8@���E@��R@��9�a�R=A�3 X�P�B��gMBa�NFLIyC�3��REQU�0<�cqwNO_H��r��,`�_SWITC�H�2RA_PAR�AMG�q ��_0mhUSE_WJ�[r
��SscNGRL�T{�O�q$WA�RNWpYp(c�STb�@J1���rAP#`�WEIGH�3J43CH�01�OR�11���bOO�@;RATI�O/�J�@D�0�bS�A��&e�ӓ�OBO4�D^0x0J2���1��bEXD_RT=QTD_IT�C���@0����a�V`RD�C�A=� � Ȏ`�`��R݀��THx?Q����RGEAPR#IO��8�W�G `�Y�?PER���SP9C���UM_�бs2TH2N�a���ѿ 1 (�E�D{1�2  D� liX�LVL2+_P���Sgq�Q~P�L10_CA�q�����a  h:q�0��j�0(S�@�qJ�H��М�Ձ� b񩓁�@�Bb�p�D��`�� P��DESIG"���1
�1�����10��_DS�q�10��FPOS11�1 l�B�ZrH��C��SATq����pU��EIND�`�1= �=0���HOME�g 	2 /ASew0�3������4);PM_q5�������L06/#/5/G/Y/k/��7�/�/�/P�/�/�/�'8?�?/?A?S?e?��S|ߠ1  �Q P��e�����ЎB T��D�FC�IO�q=II�0bO�_OPIEaC�B���� WEӁ �@H�����D �C��B$DSB�?pGNA���v�Cx���PBS232#E'  �9��5H�3`gICE��SPE����Q��IT�Q qOPyB��RFLOW�P�TR1��Q��U�SCqUPi�a�UXT�a|�Q�`ERFACTڀ�U%P��RS;CHca! t�Ր�_	P`^�$FR?EEFROM�PPs�Aq�(�A`ۑUPD��)��PT�0&eE�Xذ�X�S!��FA��p2b��@PdPca"�� 塏5�A�L�q�9P�EX`PIHQb�P1PY8e�B_�r0��4aQSfWR�a�?��9DP�wfP��6FR�IEND:�p$�UF��t�`TOO�L�fMYHՐ�bL�ENGTH_VT�E�dI�q�c��$� �`�hUFINV�_ y�ARGI��q6�ITI��gXؕ��g=vG2=gG1�Ga^P��WrhwPRE_�b���D���a�� ���S�cEQӀC��b��q�v����lS~Q# @.@P�Q꒬zWhpjU�jU��B�|�P�T$X �-M�PCTQcH��YhPP�/U)d�SG��WI`�m�҂�D��a@K�q���ʰ������=$�v 2#�qa� wi1�hr`2uk2
�3uk3�j։-��i��I��60`�0`!�$)V��bV>uV!��qQ	�q�rP%7�kV ��ߡ_��vCR�����b_�Z���Ee���c����5$AG���PR����p�S!�PR�q�R&A& �����+�ˀ$�В�ˀ%�π�P�p^Pβ
@�S^�A' ؠ�R�Ѹ7A\�/@UNN�@A)X%Q�pA�`L�ar�^��THIC��G����@�^PFEREN|Z���IF_CHkc´�Iug���6��G1@���0$���p<�7_JFE�PRL�_���RVW�A~Q( � $X�;Q  .^�VALE� ��j��:�)�Bn�  2(� �S,�0*
/  �$�_���a�����γT�Ь�γgDSP嶫�LILSpE
��A��šȳ���AX��UVK�P_M#IR�!āpMD�B�AP2� �E/`b�AԎ��SYS8�R��P�Gw�BRK�r�VNuC��I�1  ��0vc��в��AD;Aγ�;�BSOCٶ3@N���DUMMY16m6�bSV\�DEfA�SFSPD_OViR��^���LD�&�ORצ0N��ֱF�֫�OV�S!FTڥ�W��Fp�Q�%Ås���alCCHD�LY�RECOV(��pT�W��M���� �������
�_��\�g @��,pVEz@.�1OFS,pC���cWD8���4����2[Ŗ��TR��	A��E�_FDO[�MB_�CMKAF�B BL ��@�hⰑ+�VlQ�R��PY�ƳP�Gi�|�A�Mz�\��P������_�M��NRMŰ9B��T�$(���Q�3T$HcBK�Qg��IOueq�YA��PPA��?�$�O�7���YB��DVC_DB/s��h� �B����2ј�1������3����ATIO"1�]Q,��Uzc�8FCAB
�tb�s=� ���0���QT�_RPg�?SUBCPU���Si��@R��P�S�p���B�$HW�_C<P�����A�kq���$UNIT��� � ATTR�Ij���CYCL��NECA��L�F�LTR_2_FI`��H��F�QLP˼����_SCT�sF�_�F_�8�
FqS�A��CHA�a� y��CRxRSD��зB��գ��Y@_T���PRO��@�9PE%M�0_�Ц�Tfw�� f���DI�`i�RAILAC4��4M��LO���c��7�b��������+PR��S�qn�W!�Ct��@	��FUN9C���RIN�ps�0o` w$8QRA� �b� �#
@	��#W3AR5���BL�q�'��$A�+��(�(DA`���!8�#�%LD�P Ѕ�33汪!�33�TI�S5ɱ��$��PRIA�QRAF
D P0�~3�Є5�8����MOI� C�DF_�`�ӸQ;PL�M��FA��HRD]YPdORG80H��ao`0�5MULS�E�`j�S���J��J6�K�F�FAN?_ALMLV5SRA�WRNYEHARD@���V`�p�P� 2QA�QƱ��_��g�AU�mPRkORTO_SBRv�E��J� v�|!�CMPINF�����D)1�CREG�vfNV�P!c��DA��`R�FL��$AM0��RG�ࠠ`HVgUCM�N��Y�#NONI�NE�PYB8jRs&� �I��ι�+ ���a$.Aa$Z$q��������,$ �o�EaG�γ��QARఄ����23#e� |�A�XE�ROB�RKED�W�a��_]m���SY��8a��fS��gWRI��f� SCTR䵼@��*�E����d8�A�B��`���f9'#��OT�OQ����ARY��r!!�����FI���,�$LINK(�1��'qc�_�c�����3O��`OqXY�ZwBYz�jsOFF���&rNrBxpB�l"�t���p �sFI� �ww����l"��_J���(�3sP���@�d�j3p���#TB�qB5�C� kƓDU���32�7"TURT@XZ3n�q�B1X�`���FLm��Р`��pu�i39�^
� 1+��K
�	Mg�\�54%S�S%�ORQ��##� ��␂�1��0�<�j�8�#QQ�OVEX���M,0��Sr��Sr��R q��@o�p�� o�B� q ,�0��Y�9����� 0�j�Y�v����S������ER��!	8"E���|�D#9�A瑠���u�%�w11AX�ӆ�1� �(r�� ���A��ƀ��쀞� ����3 ���`���`��1fp���0���0���0 ���0˩�0۩�0��0 ���0��0�8�,�� ��2~�DEBU}�$x!�C���JrA!B'�8�R�V�| 
©��/�m ;�e�;�Ɓ;��;��� ;�3!;��a;��a�4:���2ϒ�sLAB�r8�y ��GRO� �}L��B_� ��d 1ӽp�@����ձA �ANDڀ8 .���Su1��A]� ��Q�``q�1��� RpNTd@�ӣ�VEL�͔���!���r�0ҭsNA��phbC�T�`s3#�,��b{�SERsVE���P- $�pܤ ��!)�PO�J�� _�T9P!��1�P. w $M�TRQ���
L�hbV�/Z�22�.k�b0 _ 0� lT�AERR��ra�I���͔��TOQ͔ʐL<`���b����G+�%<q|� � L�RE0 1� ,'�o��/ёR�A� 20 d�0�f��P�b� 2�P$f���0����OC1x�3 � ��COUNT��a ��PFZN�_CFGU�4 4� %V�T|�z��ೌ���� 4 ���S5 �,�M�+B�`�pɓo��FAq0ؕ6XX`-	��H�Ga,�� XaPzB��PHELAP��6� 5�pB_B;AS|�RSR$V` ERcS<L1� 1�窙 2�
3�
4�
5*�
6�
7�
8���RO�� �-pQpNL��Q@�AB8�
 � A�CK�IN^�T_�UUU�@	@�AL_P�UX�~Be2OU:�P�� %Xy��@�`y�T�PFWD_KAR���-Q��RE7��0P8#p1� QUE$Yf� Y�I���~@�AIU@��yOp���VOqSE�M�q?&E��0AS�TY[SO* P�D�Ig�@��!x��1_�TM9SMANRQܘ&OpENDN�$�KEYSWITCaH��z!$HEI��BEATM�PE�(`LE��� ��(UҾF.$�S$DO/_HOM�0OzAOEF9�PR�q��ja�`UUC
0O�1���OOV_M��pE�pGOCM;�'E�D�vxHK�Q7 DLq$&W��U��"M`��K�<�FORC*SW�ARձ�RzOM>` 8 @���s*�@U�cP`1FgP�D3F4��c�O��L�29�%XUN�LO���ZDED>�A  �S+0��G: <NP�1y���MSUPGN��AC�ALC_PLAN��C1�pAY�a�|zB��; � �@9�PA�$�MQ{Aϵ���`���%Md0���r��F�Td��RSC��M �P�ѱ� �<Q���p�jOTYWZZWZEU AR㐡PTaՈR�P�V~�2NPX_AS��w< 0� ADD����$SIZeA�$VA���MUL�TIP<�S@A��1= � $ ��P>2�p6bS��ayC��"fFRIFa��^�S�IB4`NF�$ODBU�`��#efcai7�CM�!$�ձ������Ƃk� >!�> � �P���TE��
��$SG%L�aT5r��&���cx���`�`STMT���sPSEG8" qByWY��dSHOWunb�BAN�@TP�p@���,��7�l�mV+�_G��? ��$PC��_�+���F�B�1P�xSP A�f�u�VD�p���@� ���A00���q@�w@�w)@��w3@�w5�y6�y7*�y8�y9�yA�y�@��w @�w���v�@�wF�x+����y1�y�`����1$�11�1>�1�K�1X�1e�1r�1*�1��1��1��:�Tx��y2�y2
�2�U2$�21�2>�2K�U2X�2e�2r�2�U2��2��2��3�yU3�y3�y3
�3��3$�31��H�K�3�X�3e�3r�3�3���3��3��4�y4��y4�y4
�4�4�$�41�4>�4K�4�X�4e�4r�4�4���4��4��5�y5��y5�y5
�5�5�$�51�5>�5K�5�X�5e�5r�5�5���5��5��6�y6��y6�y6
�6�6�4�6A�6>�6K�6�h�6e�6r�6�6���6��6��7�y7��y7�y7
�7�7�4�7A�7>�7K�7�h�7e�7r�7�7ꌉ7��7������pP_UPD�qAs Z��C 
J��V\b�qB x �$TOR��`  �7SO�� l ��Q_w�RE�r��'��`��S��C1����_�U;`�� J�YS�LO�C �  �Udb��Qd�W$05�0<�RVALU��q����R�F
�ID_YL�#z�HIu�I�2?$FILE_���Ƶ$?3�0�SA�V�qD h����E_BLCK���q>��D_CPU���P ���Pu������� ��R E � �PW�`.I`XLAqSR��]ngRUN�@G�\��g� ��\�gH`�s� g�AT2��_LI�2F  ]'G_O:"��P_EDI2�PTo2SPD�G��PIDq`I`
�D�CSy Gi�H � 
$JPCwT�s� SPCOC^�$MDLQ$�u0~TCP�UF�� SCOB�� ��<�r�pI�0"M\��Oz~r?TABUI_<�pyJ�B< HD".RI$2#A�S�`�LLB_AVAI�2�q2#�qK $n� SEL� NEs.� RG_� N�`�A�x@2#SC�0LS �o!B@TB�I01!_M�@�pM 1\��PFo1L_���&)M�b-@G�pUy2]t]6:rPS_XbP�`� �P,5Ew"�TB;C2�EN ��`�@l�@�B$�FT@pqag4"PZ�TDC�e�� �0�P;c�5{7THDX`�1�4��7R�{$�PERVEn3��4{3�4�aF2_AC��0 OX -$A�@n3D{3@� rPI`aPLOW�'F1A��2HG*P���`3C\`ERTIA�5T��pI��@�KDE|�EXaLACEM��CCcC��V2�P�F8�E�G�ATCV�L�A�GTRQ�LUZ�r �C�q:U�C�qJQ��DQZ�Ja��p�E�Q
�EA2� 9p*!@l�C�0JK�VVK|q �Q�1�Q�a�PJpq�Q��SJJ�SJJ�SAAL�S�P�S�P�V�a2�R5�3)PN1\)`�K�@uD�!_qq`R�vG1CF�"P `��GROU`��aZB�q�N^0CpS�`REQ�UIR�2>�EBU�3�1�� 2aO�a�0�fG1SGL5�Q�  APPR�PCw ��
$� NN�hCLO-yS�5Xy�E0 BC� AR �d0M�0�@P��2Wt_MG��apC��p��kx�0lwBR�KjyNOLDjvS?HORTMO��z$�}[uJ�!3CP�T�@ �S�@�S�@c�@c�@#1�r7�u8�1�0>M4S� �b(B�n1G��1U�PATHQ�j�`�j�-Hf�GpZ�`R��NT� A%ذw�b`qIN BUCht@[A��C?PUMɈ	YJ@# iPЁ~��1�늣0��P�PAYwLOA�wJ2Lf�'R_A� *�LY 6��2�&�B�kuR_F2�LSHR�4o�LO�7���p�̓~�̓AC�R���������2H�S�uB$HkrޒFWLEX�c@qJK6T P�b\?n?�?�?�Z@�� EU : OF�@p���"O�1�@+O=OOLF1��ե駀^OpO�O�O�O�O�E �O�O�O�O
__._@_ R_��TW��T��� s_�_�_���ZTa��X��gQ�U\�D��U�� ���_�_�_�P�Ue�U�eo1oCoUi}!BJhdV �W0uo�o�o�Z�g�AT��a^PE�Lp��"�ҳhJ�`Uv�`JE�pCTRw"��N���֤gHAN/D_VB���_��M4W� Q@kv�46M�SW���G0EvX� $$MT� Xy���q��q�쳰���r��A��#�[v����d}Au|C��zA�{A��{��v{ �zD�{Dʤ{P��Go m�STЉwu�yu�N�xDY � �`kv����4�@f� ��f���%��WDį����uP�u�u�
����%�.� z�L5Y w�\�O� *�s)q�ASYM��P`��`��XR`������_SH\b��؄�}�H� ����*�J1��p�C�cYb��_VI�+��)s�V_UCNI�3���n�J�U ��������& ��^P���pß՟f%�����D2E�pCH~h Z �l�dO�TO��PPD��V�3�$�5��R��P��q��Xq� �$�!� _�u����0�%�!����P�ROG_NA�}$Tj$LAST�q�R�CAN���3� XYZ_SP���$X7�� �l6S� 05q1sEN�p14CUR�(�5��`HR_T�b[A�1y3N��pS��O�4���0�\ ����I�A�$�� A`��C����r���0 ] � Y�MEX���)Bc"�T�0PTFe�q�QAU`Yd�(VHqA�eITGZa $�DUMMY1��o$PS_ �RF �  q��F�FL�Aj`YPR��BYC?$GLB_T���5p�EQ@�@pLIFh�^�E��f�@OW�+@O�UVOLY�L� 0Q_2Ɂ�D2.���@�pP�6R�00S�@T�C�$BAUD,��SST6�B��@�ARITYpSD_[WA�TAIUYC��r�OUv��Q�YT�LANS�@�[��SyZ\C'�BUF_�R�L����X�0�YCHK]_0CESɡ��+JOG@E�AQ!4hRUBYT:�KiH� Kd�rn�nf`�Q��!�čfH��>���1_ �X
���aSTY����SBRU M21�_� �T$SV_cERR�e�cCL�@��bAq�O�"�0GL��EWh` 4 �$[A$�Q$�Q$W3sy��!U�#0Rɂ�@sUua� b�"4$GI��}$q q`tLphb L$p\nv}$FEvv�NEARR�?2$�F�yO�TG1��/�J�0R�� cc�?$JOINT����f�qMSEThd�  kwE�ur���S��_�t��he�k  ��UX�?���LOCK_FO���`��0BGLV�GmLg�TE:0XM�N&�EMP�pz����BR�$UP�r{ #2a��Ls��b|�\�4W���`�aCEo�s�Ҁ $KAR��M>�3TPDRAp�qVEC�� ��pI�U��c��HEY�T�OOLɣ%�VȤR�E�IS3H�E�6L/��!CH�� d�1�ONWE�D3Wc;�I��"6P@$RAIL__BOXE{!��gROB0��?��a?HOWWARp!��<�@m�ROLM�BǕ�d�j�ؒ��6P�;�O�_F��!��HTML5x1K3��P��]p_�hf�~� � �W�hg�r���q��8Vv�Phh t�Э��`NA�Ҵ�R���POJ[�1IS0��NP��;���_����2��!ORDEDW�� Q��p�XT��%1)�2R0M�O@ i D �@OB���W� ��C�@���SYS�ADR�Ѱ0Q@|� �� j ,b�NV$A^�!5\�|=5�APVWVA,A?k � 0r��5PR�"$E�DI1��VSHWeR������IS�p�Q`ND;@wcس�cHEAD+` �;���KE�Q�@CP\i0�JMP�L�5C�TRACE�4�l��Q�I��S��C%�NE.����OTICK/��M�1��!2�HN�am� @��O��7C7�P8�6���@STY�"k�LO�A�"2�ens�
0 6%$���"4=��SW�!$@�{ @A�Ea�EP� Έ6SQU�RLO<�B�TERCU@Z��TS�o  up�`�׭ s������1OV@ICU IZ�D"1�E�A%a�B���A�P9P�R��_DO?2[��X�PS�1�3AXI��Q����3E� Tx���P�REQ_��,�ET-�*P33����F���A��e�D9BX�0 �q�TSRdpl mз����s��
���B��VJ1��h���A���q��@��A8���I���� ��D+��P?�$��C��,�C=�p%7I^SSC�@� q h�DS������@SP� A	T*�J2�ь�[BoADDR)c$�P�� IF3��_2C�H+�/`O���m ��TU�`I�� rF�rCU�PN���V<�I�2sM�t�.�C�
��
VrVj����0't \�`��������@0�C^��Q��
����b��TXSCREE�u�0_P���INAs|pL"4p�.�.Pv TA� �`�B,��a�����+��ҕ��RRB`�q+����D;�UE7�w# ���!a�@Sq,�'RSM����U۠W��6!�0S_Fs#&�� !&)A'��.�CL��ހ 2vGUE���x�2�bf&1M_TN_FLj��1x�`��@�BBL_o�9W�@�0y ����"5O@q�"LE^�#x����$RIGH�T�RD�dTCKGRĂ@5Tܠ
71WIDTHBSͰB���A�+b��UI��EY���z d$p
�Ɛ���6P��BACK����B~5q4@FO�ɡ�7LAB��?(�4@I-�P�$URL���0 V1:@H�� { 8 $��0T_�l�2;@R �PR�GSu��AU2�P�f �`|��w�PU�� /CR`�ґLUM8/C�N ERV����I�`NE^4} � b�GE�2�qY�L��LP�EW�ET���)�G��H��HY�*�I5�K6�K7�KMP��@RҚӸ��pDU1xY�=`A |V1�USRt~ <ĺ`�0Urr�rrFO\� rrPRIj�my���рPTRIP���m�UNDO6�ipЙP�չ���p���+�` ��2\KP$aG ��T되��m�ROSr��VR 1��S+��!�"4s ;~b�����U�A�!��o.o<#�B���SOSFF��� � Dc�O�`�����d�d��GU&�P�a\��c����gk1SUB�� }��E_EXE6��V���SWO�� e�c`�W�WA���KPq�0J V_�DB-sEp RaR	T`�䅖��q��;#sORo�uuRAUD "vtT�yD�[q_��7��� |��D�OW�N��s$SRC���0�D���u��M�PFI����-�ESP�є�d=�^CޱZG�K���u���� `�e`rs��2�COMP�$���P_�p`x�o�k�v�7rCT3�q)�qK���DCS�ŐPL��4 C3OM\PZ�Q�{�@xҏ��}�HcCq�a���o�VT�Qg`
�bY�Zޱr`K�F�� �ѷSB$�>�r���_�M*�e��gDIC_�AY�.��PEE0T�1��#VRq���1������0C�� <����� W���~ Gg5�vsF��ܴ�� ��SH�ADOW�Q
�_�UNSCA���OyW���DGDE_LEGACi�����C��C\c�� A��%������R��w�0�w�@Cr@w�D�RIV��8��C��!��h�� ܂ MY_UBY+T���c ��1�d)��0�̱�_ ���&�L��BMv�!$Z�DEYI�cEX� ��o�MU&�1X=�l� US*��{P_RbC�pPc���D�G_�PACINj��RG�q����zc`��9c��K#o�RE�2�ba\�\���� �S � a�G��P/H����]�R`� �f0�(@�L1�b	n���RmE=�SW��_A���� k���OAQ-1A(o�s¨�E��U��ϒg T0]�HK���%@��EП�o����EAN��prprżEP]�MRCV�!�; �z@ORG�Б�¤2	Ҍc���REF�'$����a�k@[� I�PP�Z��Z�)�|�ֱ�_�p�ʲ�����SP��ˣڅ�Q]��$� ��?�Q\Q�Х�OU�؛� g����2�� 0Mq�jP�-���F� N UL_ �f.�CO�i��\�Y�NT)��䩂��A��8Q��e�L)���0����A��8Q�VI�Av� �pHD<w v0$JOP�"��$Z_UP|���Z_LOW5���d��1�"���$EPY��S�Y%��@�G\FG �q���o 5-PA81{ -CACHf�LONѷ���]���C1T���C��I_F�����T������$HO�rps��Á���O � 3�L2���q}A���VP�� 0�_SIZf��Zd��5�؇7q3MP�
FA�I��GV���AD�	o�MRE����GP R��py�AS�YNBUF�RT�D-9�3OLEO_2D_tcUW9c$����UK���Q���ECCU�VEM�հ�����VIRC �M5�9_~�jX�P�P�AGIR_�GXYZE -#_�W/� (L�$k1�Tb�L��IM�L�C0��G�RABBa<�{�L�ER��CN�{�F_1D(���.V50�()���%B���䒬���2LAS902ћ�_;GE��� ����q�O�%T���b�/��9R�I4����B�G_LEV�1��PaK����Q�GI� 	N�0t�Z��0�����k��P��S� ��N$�4 �L
q����σ�cAO�*SbD�QDE�Y��q�8��8B�W��v���p�b�WP��:ڄ0T8S��Q�D�tQ�   �rPT�ĂUfq� $&qIT�RyP�1���b�VSFd���  ��Po���_�UR��S�M�U��R�xAD�J]@���ZD�F�3 DHV�AL?�� �t U�PERI�"�$MSG_QM�$���P7r��gp���RzG�Q^�cG �X�VR�T��"�PT_����2��ZABCBbu�RڃC�
XA��AACTVSg� � � $�U<3 
SCTIV�1G�IO���SB��ITlU���DV�
���Y0���q `P	Sݑ�r ��rGސaGLST��G��lM�\f_S������A��CH�r� L mq�c�U���j�D���� GNAET`��G��_FUN?�G �Po�ZIP�t�TR�Q�$LˢA��RMPCFbu��Bp�R��qڡLNK0�
�	q ct� �$@��tCMCM��Cx�Cb�Zq0��P�Q $JxsrtDv~r�r�w����u��rw�ԍr�wU9X!uUXEq��v !�u�u�u�q�q�y�q�wpFTF��~s8��2�
�Z�e� ��K�d �0R�Y�^�Dg  � 8��R� U�$H�EIGH��zH?(�a�gVB�qPR�䥏 � �D/ѱP$�Be�����SHIYF�HRV��FPC����PC�srhqx䀈@���3p�#9�kD,I�b`CE�PV!�P�)�PHER�� �� ,a���������y@GNp�)� � �������X@X@�Q ���IORITY �P��ʒ����$`SP�@�����ԕ��;���8�ˑגODU��x�����W�5��G�GL�H�1�H�IBHQO���TO�E�1D�  _(!AF��E ��ӯާ!tcp|ޯ�!ud��~.�!icm��V�5�XY�� ��� �ԑ)�� *������X@� ��Ϳ��������� �S�:�w�^ϛϭϔϐ�ϸ����*4�p�����%+�=�O�a� o>��/c�	�=/�� **:��哈9߮�����ض�A}��,  �ΐ�����*��`���Z��m�������ENHANCOE (���A>��d�����  �D1�����ѓ�����QkR�X@�|��RTREP�<w�g�SKST�`�SLGu 渫���ԑUn?othing��� �� ��CUgY����TEMP �D�xz�4 _a_�seiban�	 Š����2 VAzew��� ���//@/R/=/ v/a/�/�/�/�/�/�/ �/??<?'?`?K?�? o?�?�?�?�?�?O�? &OOJO5OGO�OkO�O �O�O�O�O�O_"__ F_1_j_U_�_y_�_�_x�_�_��VERS׀�A�` di�sable��]S�AVE 	D�	�2670H70%0�X�_po!��ro�o/��o 	�h*�|�$�o�e�o�e;M_qz*|�o��9�/gƁ 1
��]`�p'��5���\'���URGh�Bu���h�WFA�������/�W̠b�K�f�WR�UP_DELAY� ����_HOT %3�,�����s�R_NORM�ALňL�Տ*���S�EMI	�/�n�֑Q/SKIP�s3��sx�_���_ן����� 3�"�0��P�b�t�:� ������ί�򯸯� �:�L�^�$�n����� ��ʿܿ�� ���6� H�Z� �~�lϢϴ��� �������� �2�D�3���$RACFG c����|��bѿ_PARAM��3��� @��@�`��|�2C���|���Cg�G�Bb�BTIF����bпCVTMOU��v���b�DCR�s}�� �ʑ�=t�B8*�B(^P@����@-�S;��޾�����}վ-?��T3�
�̟����;e�m���KZ;�=g;�?4�<<���J�8���� �:� L�^�p���������������� }�RDIO_TYPE  7���u��
EDPRO[T_f���C�|�BHg�E��X���2h ���B��Я�
����� �+�\[��� �ߴ����"/ /F/T'rw/��>/�/ �/�/�/�/�/�/�/? B?d/i?�/�?$?�?�? �?�?�?O�?,ON?SO r?$O�O O�O�O�O�O �O_�O(_JOO_nO0_ 
_p_�_�_�_�_�_�_ o4_9oKo
oloo�o ~o�o�o�o�o�o0o 5TohV�z� ����@1���~XINT 2ȉz��q�G;� o������祐j�f�0 Ǐً����	�� �S�A�w�]������� џ����۟�+��O� =�s���k�����ͯ�� ���'��K�9�o� ��g�����ɿ��ٿ����#��G�T�EFP�OS1 1'	  x���t ���ϩ����ȈϚ��� 5� �Y���}�ߡ�<� ����r��ߖ���C� U����<�����\� ���	����?���c� ���"�����X�j��� ��)��M��q n�B�f�� %��mX�, �P�t�/�3/ �W/�{/�/(/:/t/ �/�/�/�/?�/A?�/ >?w??�?6?�?Z?�? �?�?�?�?=O(OaO�? �O O�ODO�O�OzO_ �O'_�OK_]_�O
_D_ �_�_�_d_�_�_o�_ oGo�_koo�o*o�o �o`oro�o�o1�o U�oyv�J� n���-���� u�`���4���X��|� ޏ���;�֏_����� ��0�B�|�ݟȟ��� %���I��F���k�2 1w�!�3�m� �֯��3�ίW�� T���(���L�տp��� �������S�>�w�� ��6Ͽ�Zϼ��ϐ�� ��=���a���� �Z� �ߦ���z���'��� $�]��߁���@��� d�v����#��G��� k����*�����`��� ����1������* �v�J�n�� �-�Q�u� 4FX���/� ;/�_/�\/�/0/�/ T/�/x/?�/�/�/�/ [?F???�?>?�?b? �?�?�?!O�?EO�?iO OO(ObO�O�O�O�O _�O/_�O,_e_ _�_ $_�_H_�_l_~_�_�_ +ooOo�_soo�o2o �o�oho�o�o�o9 �o�o�o2�~�R �v���5��Y���}��������3 1��N�`����� <�B�`���������� U�ޟy����&���ӟ ����k���?�ȯc� 쯇��"���F��j� ���)�;�M����ӿ ϧ�0�˿T��Qϊ� %Ϯ�I���m��ϑϣ� ����P�;�t�ߘ�3� ��W߹��ߍ���:� ��^�����W��� ��w� ���$���!�Z� ��~����=���a�s� ���� D��h �'��]��
 �.���'�s �G�k���*/ �N/�r//�/1/C/ U/�/�/�/?�/8?�/ \?�/Y?�?-?�?Q?�? u?�?�?�?�?�?XOCO |OO�O;O�O_O�O�O �O_�OB_�Of___ %___�_�_�__o�_ ,o�_)obo�_�o!o�o�Eo�o��Ƅ4 1 я{o�o�oE0ioo �(�L���� �/��S�� ��L� ����яl�������� �O��s����2��� V�h�z���� �9�ԟ ]������~���R�ۯ v�����#���Я�� }�h���<�ſ`�鿄� �Ϻ�C�޿g�ϋ� &�8�Jτ�����	ߤ� -���Q���N߇�"߫� F���j��ߎߠ߲��� M�8�q���0��T� ��������7���[� ����T�������t� ����!��W��{ �:�^p�� A�e �$ ��Z�~/�+/ ���$/�/p/�/D/ �/h/�/�/�/'?�/K? �/o?
?�?.?@?R?�? �?�?O�?5O�?YO�? VO�O*O�ONO�OrO�O<�o�d5 1�o�O �O�Or_]_�_�O�_U_ �_y_�_o�_8o�_\o �_�oo-o?oyo�o�o �o�o"�oF�oC| �;�_��� ��B�-�f����%� ��I��������,� ǏP�����I����� Οi�򟍟����L� �p����/���S�e� w������6�ѯZ��� ~��{���O�ؿs��� �� ϻ�Ϳ߿�z�e� ��9���]��ρ���� ��@���d��ψ�#�5� G߁�������*��� N���K����C��� g��������J�5� n�	���-���Q����� ����4��X�� Q���q�� �T�x� 7�[m�// >/�b/��/!/�/�/ W/�/{/?�/(?_ T6 1+_�/�/!? �?�?�?�/�?�?O�? OAO�?eO O�O$O�O HOZOlO�O_�O+_�O O_�Os__p_�_D_�_ h_�_�_o�_�_�_o ooZo�o.o�oRo�ovo �o�o5�oY�o} *<v���� ��C��@�y���� 8���\�叀�����ޏ ?�*�c�����"���F� ���|����)�ğM� ����F�����˯f� ﯊�����I��m� ���,���P�b�t��� ���3�οW��{�� xϱ�L���p��ϔ�� �������w�bߛ�6� ��Z���~�����=� ��a��߅� �2�D�~� �������'���K��� H������@���d��� ��������G2k �*�N�����1�U;?M47 1X?N�� ��/�8/�5/n/ 	/�/-/�/Q/�/u/�/ �/�/4??X?�/|?? �?;?�?�?q?�?�?O �?BO�?�?O;O�O�O �O[O�OO_�O_>_ �Ob_�O�_!_�_E_W_ i_�_o�_(o�_Lo�_ poomo�oAo�oeo�o �o�o�o�olW �+�O�s�� �2��V��z��'� 9�s�ԏ��������� @�ۏ=�v����5��� Y��}�����۟<�'� `��������C���ޯ y����&���J���� 	�C�����ȿc�쿇� ϫ��F��j�ώ� )ϲ�M�_�qϫ���� 0���T���x��u߮� I���m��ߑ����� ���t�_��3��W� ��{������:���^�����hz8 1 �/�A�{�����#� A��e b�6� Z�~���  aL� �D�h �/�'/�K/�o/ 
//./h/�/�/�/�/ ?�/5?�/2?k??�? *?�?N?�?r?�?�?�? 1OOUO�?yOO�O8O �O�OnO�O�O_�O?_ �O�O�O8_�_�_�_X_ �_|_o�_o;o�__o �_�oo�oBoTofo�o �o%�oI�om j�>�b��� ����i�T���(� ��L�Տp�ҏ���/� ʏS��w��$�6�p� џ���������=�؟ :�s����2���V�߯ z�����د9�$�]��� �����@���ۿv��� ��#Ͼ�G�����@� �ό���`��τ�ߨ� 
�C���g�ߋ�&߯������MASK 1���������?XNO  �� �~�MOTE  "����X�_CFG �_��Tԓ��P?L_RANG[�W�������OWER ������SM�_DRYPRG %���%\����TART ����UME_PRO�����v���_EXE�C_ENB  <���GSPDO��v����TDB�����RM����ING�VERSION �#�e���I_�AIRPUR�� �W�0�l��MT_���T��]����O�BOT_ISOLEC ��h ����/NAME�-���OB_CATEG ���1�$�8@�ORD_NUM �?��eH700  T��{����PC_T�IMEOUT�� �x��S232x�1� #��� L�TEACH PENDAN�tד�$�[�Y����� ���� ce ConsT��/-&"'/U���ֳ e-W//~K�No Us�/p�/�/�NPO)�\������oCH_LR�!���	F1?!U�D1:l??R��VGAIL\�T ����PACE1 {2"#�
? ���,zӑ��U i�)L< ��0?��;PO�?0O�O�O~O �O�G�?�?OO�O>O `OV_w_6_�_�_�]#� #��]�O�O__�_B_ d_Zo{o:o�o�o�o�o �O�_oo,o�oPoro h�o�����o�o (�Lnd��� D�������Џ� �� $�6�H�Z�|�r�@��� ��ɟ������ �2� �V�x�n���N���ů ��گ��
��.��R� d�j���J��������� ����*�<��`��� xϙ�HϺ��϶���� �&�8���\ώ�t��πTߪ��ߢ���;�12�<� �?�*�<� ��`ߒߕ���u���������3�'�9�K� ]�������������"#�46�H�Z� l�~�0������ .CD5Wi {��Q���>@�./O/&/d/e6x ����r/�/?�_/�/O?p?G?�?�/7 �/�/�/�/�/�??7? :O�?OpO�OhO�O�?8�?�?�?�?O�O&O XO[_�O;_�_�_�_�_��OG &�K� �_�
(` o  �EHoZolo~o �o�o�o�CX�m_�_�o�_2�dHp-o?o m������o �o�n�z!�3�P�CU �������ˏݏ�� �	��=�O�p�c�u� ����ǟٟ�������)�;�]�o� `�_ @Ш������������� �����*�l�~���R� ��ƿؿ�������2� ����JόϞϼ�r� �������������R���"�
֯���_M?ODE  �IR^��S '�K��L�J�/_ү��M�r��	m��+�CWOR�K_AD����{n-�R  �K��@������_INOTVAL��T��C~��OPTION�� �N V_D�ATA_GRP �2)(��AD��P ��o���~������� ������,<> P�t����� �(L:p^ �������/  /6/$/Z/H/j/�/~/ �/�/�/�/�/�/??  ?V?D?z?h?�?�?�? �?�?�?�?O
O@O.O dOROtOvO�O�O�O�O �O_�O*__:_`_N_��_���$SAF_DO_PULS�����/�c�Q�PCAN�_TIM�ў�0���QR */��0���/&`&b,ら�A�cK��Q��  ��6oHoZolo~o�oo��o�o�o�o�o�o��b27t�Q�QdCx:qJq���Sy��������fy�z \��t��_; ��  T�����#�5�B�T D��B�k�}������� ŏ׏�����1�C��U�g�y����&�xz���ڟ쟱� � @�;�oȨ�
�K�p���
�?t��Dik�a>7�  � ��b�� e�Q��F��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�N���r� �ߖߨߺ�������� Q�%u.�@�R�d�v����������0 �r\�S�h���!�3� E�W�i�{��������� ������/AS ew������ �+=Oas �������\� /'/9/K/]/o/�/�/ �/�/"��/�/�/?#? 5?G?Y?k?�����b �?�?�?�?�?OO)O ;OMO_OqOI�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofoxoM�衟Q��o�o�o �o�o,>Pb t�������z��o�$�.����2��	12�345678s��h!B!��W 
F��`�� ������ʏ܏� �� $�*��oM�_�q����� ����˟ݟ���%� 7�I�[�m�~�<����� ůׯ�����1�C� U�g�y����������� ����	��-�?�Q�c� uχϙϫϽ������� ��ֿ;�M�_�q߃� �ߧ߹��������� %�7�I�[�m�,ߑ�� �����������!�3� E�W�i�{��������� ������/AS ew������ ���=Oas �������/ /'/9/K/]/o/.�/ �/�/�/�/�/�/?#? 5?G?Y?k?}?�?�?�?�?����?�?�5�/�O1OCO_�Cz � A��j   ���h2�}� >OF
�G�/  	��2�?�O��O�O�O\�oL� �OR_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o7_�o�o �o&8J\n ���������"�4�B�A�A�B�<_� U��A  �o���sC�u@l��A�At  �v@��ŏ�@(ۃ `Rl����iMu@0\��$SCR_GR�P 1,0+�04� � ���B |E	 `��h�y�r��^�~E����������ڟRM��@גD�#\���כ0\CRX�-10iA 01�23456789�0�@N� \��@fN�0 k��A
X�j��	���K ��h��W���W�0S^�"בv�����	�����*�<�N�^��G�H����l�W� ������ſ׿���o�A��Ϯ�?�XG0�w��\Ch_@,[}xx�  �䄑B� � BƊψ¡Ą�Av@��  @�@�ń�s@����� ?����H��߳ʄ�F@ F�`+�3�*� W�B�{�fߋ߱ߜ��� ���ߤ�������$��!�3�E�B�S��ߙ� ������������ ;�&�_�J�����/^�ß����|G�@��"@I���e@M7 B�bX������?�TA�����$��� 0Q��A ���/��DPb1 (�@�(����{��� /)L�����='£�7�ECLV�L  Q   ���Ǣ� Q@P!L_DEFAULTX$�L!��@~l#HOTSTRx-���"MIPOWEKRFW ZE�%�$oWFDOy& �%�6�ERVENT �1-_!_!�# L�!DUM_EI�P/8�j!AF_INEx =?TO!FT?l>3?r�?!���? �?��?!RPC_M'AIN�?�8��?(ON�3VIS�?�9�O�tO!OPCUA�uO�JcO�O!�TP�@PU�O&9d��O_!
PMON?_PROXY_)6Ae�OX_�B&_"=fG_��_!RDM_S�RV�_&9g�_�_!#R��o'8h�_<oK!
�0Mo_#<i+o��o!RLSYN�C�o�i8wo�o!�ROS?�l�4��o !
CE�@MOTCOM!)6k�l!	5rCONSdm(7l[�!5r�WASRC�_)6m��!5rUSB��'8n�P�!S#TM� j�%:o?�����?���S����#ICE_KL ?%�+� (%SVC�PRG1�1��2�1�6� �3Y�^� �4����� �5���� �6џ֟ �7���� �y�$A�<�9I�N��o v� �#��� �K�Ư � s�� ���� �ß>�  ��f� ���� �;� �� �c�޿H����H� ��.�H�ܯV�H��~� H�,���H�T���H�|� ��H����H�̿F�H� ��n�p��� � �� �����@��&��J� 5�n�Y��}����� �������4��X�C� j���y����������� ��0T?xc ������� >)bM��� ����/�(//�:/^/I/�/�_DE�V �)��UT1:�'4����$GRP 21��%� �bx 	�� 
 ,�  �/?�"�/.??R?9? K?�?o?�?�?�?�?�? O�?*O<O#O`OGO�O �O�/�OqO�O�O�O_ �O8_J_1_n_U_�_y_ �_�_�_�_�_o"o	o Fo�O;o|o3o�o�o�o �o�o�o�o0T ;x�q���� ��_o,�>�%�b�I� ��m��������Ǐ� ���:�!�^�p�W��� {���ʟ!���$� �H�/�l�~�e����� Ư������� ��D� V�=�z�џo���g�Կ ����
��.��R�d� Kψ�oϬϾϥ����� �����<ߓ�`�r�Y� ��}ߺߡ߳������ ��8�J�1�n�U��� ���������U�"��� F�X�?�|�c������� ����������0T ;x�q���� ��,>%bI ��������/�:/!/3/p/�#d Խ&	^/�/�/�/`�/�/�/?";%�"?<G?�#���`11 `5p?~7h?�?�?�?�? �?�94?O\9�?FO4O jOXOzO|O�O�OO�O *O�O__B_0_f_T_ v_�O�O�__�_�_�_ oo>o,obo�_�o�_ Ro�oNo�o�o�o :|oa�o*��� �����T9�x �l�Z���~�����ď �,��P�ڏD�2�h� V���z����ן韠� ��
�@�.�d�R��� ʟ���x��Я��� �<�*�`�����ƯP� ����޿̿���8� z�_Ϟ�(ϒπ϶Ϥ� ������@�f�7�v�� j�Xߎ�|߲ߠ���� ��<���0���@�f�T� ��x��������� ��,��<�b�P����� ����v�������( 8^�����N� ��� �$fK ]6~��� ��>#/b�V/D/ f/h/z/�/�/�//�/ :/�/.??R?@?b?d? v?�?�/�??�?O�? *OONO<O^O�?�?�O �?�O�O�O_�O&__ J_�Oq_�O:_�_6_�_ �_�_�_�_"od_Io�_ o|ojo�o�o�o�o�o �o<o!`o�oTBx f�����8 �,��P�>�t�b��� ���я�������(� �L�:�p�����֏`� ʟ��ڟܟ�$��H� ��o���8�����Ư�� ֯د� �b�G���� z�h�����¿��ҿ(� N��^���R�@�v�d� �ψϾ� ���$Ϯ�� ��(�N�<�r�`ߖ��� ���φ�������$� J�8�n�ߕ���^��� ��������� �F��� m���6����������� ��N�3E���� f�����& J�>,NPb� ����"�// :/(/J/L/^/�/��/ ��/�/�/? ?6?$? F?�/�/�?�/l?�?�? �?�?O�?2Ot?YO�? "O�OO�O�O�O�O�O 
_LO1_pO�Od_R_�_ v_�_�_�_�_$_	oH_ �_<o*o`oNo�oro�o �o�_�o o�o8 &\J��o��p �l���4�"�X� ���H�����ď ֏���0�r�W��� � ��x���������ҟ� J�/�n���b�P���t� �������6��F�� :�(�^�L���p���� Ϳ��� ϒ��6�$� Z�H�~������n��� �������2� �Vߘ� }߼�F߰ߞ������� ���.�p�U���� v��������6�� -������N���r��� �������2���& 68J�n���� 
���"24 F|���l�� ��//./��{/ �T/�/�/�/�/�/�/ ?\/A?�/
?t??�? �?�?�?�?�?4?OX? �?LO:OpO^O�O�O�O �OO�O0O�O$__H_ 6_l_Z_|_�_�O�__ �_�_�_ ooDo2oho �_�o�oXozoTo�o�o �o
@�og�o0 �������� Z?�~�r�`����� ��������2��V��� J�8�n�\��������� ��.�ȟ"��F�4� j�X���П����~�� z�����B�0�f��� ��̯V������ҿ�� ��>π�eϤ�.Ϙ� �ϼϪ��������X� =�|��p�^ߔ߂߸� ������������� 6�l�Z��~������ ������ �2�h� V��������|����� 
��.d��� ��T����� l�c�<�� ����/D)/h �\/�l/�/�/�/�/ �//?@/�/4?"?X? F?h?�?|?�?�/�?? �?O�?0OOTOBOdO �O�?�O�?zO�O�O_ �O,__P_�Ow_�_@_ b_<_�_�_�_o�_(o j_Oo�_o�opo�o�o �o�o�o Bo'fo�o ZH~l���� �>�2� �V�D� z�h�����׏��� 
���.��R�@�v��� ��܏f�Пb������ *��N���u���>��� ��̯��ܯ��&�h� M������n�����ȿ ��ؿ��@�%�d��X� F�|�jϠώ������ �ϴ��ϰ��T�B�x� fߜ�����ߌ����� ���P�>�t�ߛ� ��d���������� �L���s���<����� ����������T�z�K ��$~l���� �,P�D�T zh����( �/
/@/./P/v/d/ �/��/ /�/�/�/? ?<?*?L?r?�/�?�/ b?�?�?�?�?OO8O z?_OqO(OJO$O�O�O �O�O�O_RO7_vO�A��$SERV_M�AIL  �E�vP�\XOUTPU}TkX�@}@`TRV 22 V;  yP (QF_<�_`TSAVE�\zY�TOP10 23>�Y d |O2o DoVohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r� ��������̏ޏ���0�&� UeYP�_]S�FZN_CFG ;4 UyS{D��Q�Uf�GRP 2�5p��Q ,B �  A���AD;�� B���  B�4&cRB21��VHELLi�6 U�V�P�_���(�%RSR(�)�;� t�_����������˯ ݯ��:�%�^�I���������  �Q%��Կ濡�������@���)�zG��2�@d��쿾ۖHK 17� ϚϕϧϹ��� �����*�%�7�I�r� m�ߑߺߵ�����՜?OMM 8�)��ڒFTOV_EN�BkT�Q�YHOW_?REG_UII�^R�IMIOFWDL��9~�WAITF�Ɉ���Pj��T��TIMj�����VAjP��~�_UNITE���Y�LCc�TRYj�Z�U`PMEi�:����Q	���f�;r�[ ������<����X�@Đ `	P?�  �����_�'P@6��V�VMON_ALIAS ?e��Phe1_��� ��
�%7� [m��N�� ��/�3/E/W/i/ {/&/�/�/�/�/�/�/ ??/?A?�/e?w?�? �?�?X?�?�?�?OO �?=OOOaOsO�O0O�O �O�O�O�O__'_9_ K_�Oo_�_�_�_�_b_ �_�_�_o#o�_GoYo ko}o(o�o�o�o�o�o �o1CU y ����l��	� �-��Q�c�u���2� ����Ϗ�󏞏�)� ;�M�_�
��������� ˟v����%�П6� [�m����<���ǯٯ �����!�3�E�W�i� �������ÿտ���� ��/�ڿS�e�wω� ��FϿ�������߲� +�=�O�a�s�ߗߩ� ����x�����'�9� ��]�o����P��� ���������5�G�Y� k�}�(����������� ��1C��gy����Z�$SM�ON_DEFPR�OG &����� &�*SYSTEM�*���RECA�LL ?}�	 �( �}/cop�y mdb:*.�* virt:\�tmpback\�=>192.16�8.56.1:11320 \mܑ�}3x5fr:\>�Pbi�(//�4�a���]�{/�/�/ }8��s:orderfil.datA X/�/�/?�4�/X �/{?�?�?�E/R?� �?OO0/�?�?f/wO �O�O�/�/I?�/�O_ _,?@O�Ob?s_�_�_ �?�?OO�?�_oo(O :O�_^Ooo�o�o�O�O A_Xo�o�o$_6_�o Z_�o}�"�_Go�_ j���2o��ho�y������q75vho�me.tpAuemp\��U�k����� �o�oM�y�����0 K�Tf���	���A� S��u�����,�=�O��b����*�\��:�ipl_fanu�c_smplgr�p_close.lsŉ=�O�կ믠� 3�E�Ο��n�ܿϤ� ��ѿڟ�Q��"�4� ǯX�j�|ώ�߲���������Xߑߤ�tpdisc 0}߀�R�d�v߈����tpconn 0 ����������*� ��=�O�a�s����� ��D�߿�����'�9� T�]�o����Ϸ�J� ����V!#�5�F�� k�� ����?� ��17�1}O as�/)�;���_� �/�/����T/��o/ �/?%7�[�/V? !?��F?�k?�?�?  O3/E/�/i?�?O�O �/LO�/gOyO�O_/���$SNPX_A�SG 2<����@Q� �P 0 '%�R[1]@1.Y1!_kY?�-�%k_ �_z_�_�_�_�_�_�_ 'o
oKo.o@o�odo�o �o�o�o�o�o�o G*kN`��� �����1��;� g�J���n�������ˏ ��ڏ����Q�4�[� ��j��������ğ� ���;��0�q�T�{� ����˯������� 7��[�>�P���t��� ǿ���ο�!��+� W�:�{�^�pϱϔϻ� ������� �A�$�K� w�Zߛ�~ߐ��ߴ��� ���+�� �a�D�k� ��z���������� '�
�K�.�@���d��� ������������ G*kN`��� �����1; gJ�n���� ��/�/Q/4/[/ �/j/�/�/�/�/�/�/ ?�/;??0?q?T?{? �?�?�?�?�?O�?O�7OD3TPARAM� =@UJQ ��	�;JP�D�@�H�D� ���3POFT_K�B_CFG  �zCFU0SOPIN_�SIM  @[��F�O�O_�@Q@RV�NORDY_DO�  �E�E%RQSTP_DSB�N��Bi_uHQ@SR �>�I � &� IPL_FA�NUC_SMPL�GRP_OPEN�u]yD�@Q@TO>�PN_ERR2_OB~�QPTN �E�
`�D�RRING_PRM�_�DRVCNT_GP� 2?�E�A�@x 	e_do|@Ro�ovo�o�WVD9`RP 1@`I�@�a�I�g �o�o 2YVh z������� ��.�@�R�d�v��� ����������� *�<�N�`�r������� ��̟ޟ���&�8� J�q�n���������ȯ گ����7�4�F�X� j�|�������Ŀֿ�� ����0�B�T�f�x� �Ϝ������������ �,�>�P�b߉߆ߘ� �߼���������(� O�L�^�p����� ��������$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@gdv�����bPRG_�COUNT�F�
b�ENBo�M�#�D/_UPD �1A�[T  
 �{Bf/x/�/�/�/�/ �/�/�/??C?>?P? b?�?�?�?�?�?�?�? �?OO(O:OcO^OpO �O�O�O�O�O�O�O _ _;_6_H_Z_�_~_�_ �_�_�_�_�_oo o 2o[oVohozo�o�o�o �o�o�o�o
3.@ R{v����� ����*�S�N�`� r����������ޏ�� �+�&�8�J�s�n��� ������ȟڟ������_INFO 1=BT%: \�	 3�w�b������?*&�?����>Y�L=�n-������h>F�d?9��]/�����>�@ ?��)��<@� D�&t����D�)�´ ��E�³��*��<��YSDEBU)G�U �*�d=)e�SP_PASS��B?w�LOG �CQ�^!  r*�#�0�  �9!�*�UD1:\x��7���_MPC���T%%�7�T!�U� �T!�SAV D���!��̱�$���SV��TEM_TIME 1E���_  0  ���#����ù�MEMBK  T%�9!̰̿9�K�[�7X|: � �'��}ߢ߲�v�����Y��r� ��@�� �,�>�P��h�z��0������� ����� ��0�B�T�f�x����e���������� *<N`r�� �������SK���$�Tf�xl�n*�X�2(�߷#� ��p)�� ��������</N/`/x7.e�*�� ��/ �$���/�/�/���2�?;?M?_?q?�?*�U�?�?���?'� ��?�?O"O4OFOXO jO|O�O�O�O�O�O�O��O__0_@�T1SVGUNSPD��� 'w��HP2M�ODE_LIM #F��{�DT2QPqQ�G��CUABUI_DCS J7w�F�'�_�$�$G��6_�\o�WG�*���9a 
?`�9o'�ISh��Scɼ�UEDIT K�_��XSCRN L��R�G M�[�U�:�eSK_?OPTIONl���{��b_DI��EN�B  �%w��aB�C2_GRP 2�N�Y���o��0Cy��s<\BCCF�`P]{�� ����v`�����!�G� 2�k�V���z�����׏ ԏ���1��U�@� y�d�������ӟ���� ���?�Q�g^�p� ������0�ٯį�� ��3�a�N��#�V�|� j�����Ŀ���ֿ�� ���B�0�f�Tϊ�x� �ϜϾ��������,� �P�>�`�b�tߪߐ� �`������ ���6� $�F�l�Z����� �������� ��0�2� D�z�h����������� ����
@.dR �v����� ��0N`r�� �����//� 8/&/\/J/�/n/�/�/ �/�/�/�/�/"??F? 4?V?|?j?�?�?�?�? �?�?�?�?OBO0OfO ~O�O�O�O�OPO�O �O_,__P_b_t_B_ �_�_�_�_�_�_�_�_ o:o(o^oLo�opo�o �o�o�o�o �o$ H6XZl��� |O��� �2��V� D�f���z���ԏ�� ����
�@�.�P�R� d����������П� ���<�*�`�N���r� ��������̯��&� �>�P�n�������� ��ƿ�ڿ�"�4�� X�F�|�jϠώϰϲ� ��������B�0�f� T�vߜߊ��߮����� �����,�b�P�� <����������p�� �&�L�:�p�����b� �������� �� $ZH~l��� ���� D2 hVxz���� ���/./@/R/�v/�d/�/�/�/�/�&� ��$TBCSG_G�RP 2Q�%�  ��!� 
 ?�   ?+??O?9?s?]?o?@�?�?�?�;�"�#S <�d�HA?��!	 HA�����5>���>�=�q?�\�5AT��A 2HOTHJ��ff?aG�?IL G>BpTOVN�t@B#E� @wA� 6J��O��M@��RjI>�#33*A�5�ABCO�OD�H�BPOQY�,_.^��HBY�ArBU�PB�t_.^�H�6�H �U�_�_�_ o=ooo�ho�o�kjh��a	�V3.002	'crx�c�`*�`�d8�"8T�O ?�S� Hqji p�m7  �3C�oY�`s�!J2�#T =�`lxCFG V��%
1 0�z���r,r��x����� �E� 0�i�T���x�����Տ ��ҏ���/��S�>� w�b�������џ���� ����=�(�:�s�^� ������ͯ2+ د� ����/��?�e�P��� t�����ѿ����¿ +��O�:�_υ��!�/ �϶/�ϼ������(� �L�:�p�^߀ߦߔ� �߸������ �"�$� 6�l�Z��~����� �������2� �V�h� (/����<��������� ��
@.Pv� �X����� *<Nr`�� �����//8/ &/\/J/l/�/�/�/�/ �/�/�/�/??"?X? F?|?j?�?�?�?�?�? �?��O$O6O�?fOTO vOxO�O�O�O�O�O_ _,_>_�Ob_P_�_t_ �_�_�_�_�_�_oo :o(o^oLo�opo�o�o �o�o�o �o$H 6X~l���� �����D�2�h� V�����HO��ȏ���� 
���.��R�@�b�d� v�����П������� *��N�`�r���>��� ��̯��ܯ��&�� J�8�n�\�~�����ȿ ���ڿ���4�"�D� j�Xώ�|ϲϠ����� ������0ߪ�H�Z�l� ߜߊ߬��������� ��>�P�b�t�2�� ������������ ��L�:�p�^������� �������� 6$ ZHjl~��� ��� 0VD zh����~�� ��ߺ@/./d/R/�/ v/�/�/�/�/�/?�/ �/<?*?`?N?�?�?�? �?t?�?�?�?�?O8O &O\OJO�OnO�O�O�O �O�O�O�O"__F_4_ V_X_j_�_�_�_�_�_ �_o�_oBo0ofo� /�o�oLozo�o�o �o,P>t�� �h�����(� :�L�^����p����� ʏ��ڏ܏�$��H� 6�l�Z���~���Ɵ�� �؟���2� �B�D� V���z�����ԯ¯�� 
��o"�4�F��v�d� �������������� *�<�N��r�`ϖτϜ�Ϥ�  ����� �������$T�BJOP_GRP� 2W����  ?����C��	��Y������X  ���Y� �,� � �x��� �@��?}�	 ��A��͔�C� G D�ǌь�>0�?>\?�е�aG�:�o���;ߴAT���Ռ�A��Ӭ�����ߦ�>�я\)?w��D�8Q��>��L��>������;iG�Ҍz�A�p�Љ� ��A�ff��0��m�������/:VM��ҹR��x��)���@��RD�Cр��щ�i�e��H�Q��ff��:��6/D�33��B   �����D�V��h�Q�Q�x���:�S1���}�,B�6?Q@��Hd��r�����d�=m�<#��
���0�;/��2d���B��� ��ٰ��"�� :kF ���� ����/4//,/XZ/�/��C��Ɛ�!���	V3.00�5�crx�#� *�� i�������* �C�  E$`� E�h Eܨ� F� F3�� FV4 Fx�� F�� F� F�X F�0��� F�F F��� Gs G� G� G�k G&�#��� Y? E@ E��� E�� E�� F� F�2 FN� F�j� F�� F��� F� F��H F�| Fʰ 9�IR�1t,H�5 *���?�2���3?���`-��ED_TCH cZ��(�#����h���d$�(�O�O���� �TESTPARS  ���SC�HR�@ABL�E 1[�  @��fւҞG�:�G��H�H�����G	��H
�H�HU����H�H�H�FRDI�O(�__%_7_I_[U�TO�_�[�_ �_oo/n�BS�_&� �Z�o&8J \n������ ���"�4�F���` �o'� W��po�o�o�o R_d_v_�_�_�X�Bm��NUM  ��U(�p��� �@��P�B_CFG �\V����@�IM?EBF_TT�A��:PE��VER�Sf�z����R 1]�KO 8zO����2� ����  �� �)�;�M�_�q����� ����˯ݯ���%� 7���[�m��������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/�x�S�e� �߉ߛ߱߿�������H�:Bۑ_P�Ŗ@ϕ�<@LIF ^&V��0ʑ����t�"��( 0
��@���@� d��W�M�I_CHAN�� �ϕ ��DBGLV�L��PF��ETHERAD ?�E
����0��7�I����ROUT!�HJ!}�����SN�MASK�ϓ$�255.���#��������#<@OOLOFS_DI�@R0�����ORQCTRL C_�K;c�?yTh ������	 -?Qcu������g��/9CPE_DETAI���>
PGL_CON?FIG eV�f����/cell�/$CID$/grp1/�/�/�/�/�/6c�d�??%?7? I?[?�/?�?�?�?�? �?h?�?O!O3OEOWO �?�?�O�O�O�O�O�O vO__/_A_S_e_�O �_�_�_�_�_�_r_�_�o+o=oOoaoso��} o�o�o�o�o�o�/+
}�o`r� ���o���� &�8��\�n������� ��ȏW�����"�4� F�Տj�|�������ğ S������0�B�T� �x���������үa� ����,�>�P�߯t� ��������ο�o�� �(�:�L�^��ϔ� �ϸ�����k� ��$��6�H�Z�l�g ��User Vie�w |)}}1234567890�� ������������2�}������2����a� s������,��3D�	��-�?�Q�c����2�4�������@��v�82�5�� q�����*�2�6`%7I[m��2�7����/!/3/�T/2�8 ��/�/�/�/�/�/F/�?2 l?Camera�ڄ/�M?_?q?�?�?�?�bE @?�?�?�>��O!O3O0EOWOiO_	  '6C� <?�O�O�O�O__�? 7_I_[_�O_�_�_�_�_�_ ?�'6��p_%o 7oIo[omoo&_�o�o �oo�o�o!3E �_�W���o���� ���o�!�3�~W� i�{�������X�W�K J����#�5�G�Y� � }������şן��� ��Ə(5��i�{� ������ïj����� V�/�A�S�e�w���0� �W� �տ����� /�֯S�e�w�¿�ϭ� �������Ϝ��W{)�� A�S�e�w߉ߛ�BϿ� ����.���+�=�O�a���9�ߢ���� ��������2�D��� U�z�����������c*	)50Z�!3E Wi����X�� ��/����.0 0;������� �//*/uN/`/r/ �/�/�/O)5�K?/�/ ??*?<?N?�r?�? �?�/�?�?�?�?OO �/��k�?`OrO�O�O �O�Oa?�O�O_MO&_ 8_J_\_n_�_'O9Et{ _�_�_�_oo&o�O Jo\ono�_�o�o�o�o �o�o�_9E���o8J \n��9o��� %��"�4�F�X��o 9EL������ȏڏ� ���"�4�F���j�|��������ğk�  o����)�;�M��_�q���������  � ə?fffB �Pߡk�����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��� �2�D�V�h�z� �ߞ߰���������
���.���
k�(  ���( 	  ;�q�_������� �������7�%�[�I�t���� �� ������[�0B Tfm�������� ��� 2yV hz������ �?/./@/�d/v/ �/�/�/�///�/? ?_/<?N?`?r?�?�? �/�?�?�?%?OO&O 8OJO\O�?�O�O�O�? �O�O�O�O_"_iO{O X_j_|_�O�_�_�_�_ �_�_A_o0oBo�_fo xo�o�o�o�oo�o�o Oo,>Pbt� �o�o���'�� (�:�L�^�������� �ʏ܏� ��$�k� H�Z�l���������Ɵ ؟�1�C� �2�D��� h�z�������¯	�� ��
�Q�.�@�R�d�v� ��ϯ����п������*�<�Nϕ�u�@ Ap�}Ϗϡ�p�w��[��� frh:�\tpgl\ro�bots\crx���10ia.xml]���� �2�D�V��h�zߌߞ߰�  ����������� �2� D�V�h�z���߯� ������
��.�@�R� d�v������������ ��*<N`r �������� &8J\n�� ������/"/ 4/F/X/j/|/�/��/ �/�/�/�/??0?B? T?f?x?�?�/�?�?�? �?�?OO,O>OPObO�tO�O�N��� �w���<< �� ?��K�O�O�O �O#_	_+_Y_?_q_�_ u_�_�_�_�_�_o�_�%oCo)o;o]o�o�����(�$TPGL�_OUTPUT sh�����`� �jfffB4  �a���o
 .@Rdv��� ������*�<��N�`�r����� ���`cell/fl�oor/wall� rite 34�56789012 ��ʏ܏� �����` �/�A�S�e�w��!������џ������} �6�H�Z�l�~��(� ��Ưد������� D�V�h�z���$���¿ Կ���
Ϣ���@�R� d�vψϚ�2Ϩ����� ���߰�&�N�`�r� �ߖ�.�@�������� �&��4�\�n��� ��<���������"� ����X�j�|������� J�������0�� >fx���F�b? $$zb�� ��:,^P �t������ //6/(/Z/L/~/p/��/�/�/�/�/�/?} �A(?:?L?^?p?�?�=�@�O�?�?�J ( 	 ?�?�?"O OFO4OjOXOzO|O�O �O�O�O�O_�O0__ @_f_T_�_x_�_�_�_ �_�_�_�_,ooPo����  << ?�o�o�`to�o�o�o �o��qo7I�oU Yk��%�� ��3�E��i�{�� c���K������ӏ� /����e�w������ �����A�S��+�ş 3�a�;�M������ͯ ߯y�˯���K�]� ��e���-��ɿۿ�� ���o���G�Y��}� ��iϗ���#ϭ���� ��1�C��/�y����� ����[���������-� ?��C�u��a��� ������Q���)���� _�q�K���������� ����%��1[�� ����=���� !EW�C��gy��gb)WGL1.XML�?�
-�$TPOFF_LIM l`�0ha��&N_�SV    �4�2*P_MON Mide4$�0�0�2)STRTCHOK jde2&%?�"VTCOMPA�TG(�!6&VWVA/R kg-�(K$� �/ ?�0�z"!_DEFP�ROG %�)�%IPL_FA�NUC_SMPL�GRP_CLOS�E�/?0ISPLA�Y' �.<2INST�_MSK  �<� x:INUSE9R�/~4LCK�<�;�QUICKMEN��?~4SCRE@�de�"tps�c~4�1.@3I2"D@_�HIST�*2)RAC�E_CFG l�g)�$0	4
�?��HHNL 2!mK:D`�A�+ !2�O �O__/_A_S_e_wZ��EITEM 2n��K �%$12�34567890<�_�U  =<�_�_<�_c  !
ok0�_Wo3�_xo�_ �o�oo�o6oHolo ,�o<b�o�o�o�o  �D��(�� L����N����ʏ ܏@��d�v����Z� ��~���􏜟�*�� N��r�2�D���Z�̟ ����¯&�ү��
� n��������0�گ�� ����"��F�X�j�� Ϡ�`�r�ֿ~���� ��0���T��&ߊ�<� ���ω��Ϥ�ߴ��� `�P�b�tߎߘ��� h������(�:�L� ��p��B�T���`��� �� �����6���l� ����k������ � �D�z: �Jp���
 .�R�$/6/�Z/ ���f/~//�/�/ N/�/r/�/M?�/h?�/ �?�??�?&?8?O�D�S�Bo�OJ� 3 �RJ �A]OT9
 jO�OwO�O~5JUD1:\�L���AR_GRP� 1p�[� 	 @�@_[_@>_,_b_P_�_t^��P �_�Z�Q�O�_�_	o�U?�  $o6k oVo Dozoho�o�o�o�o�o �o�o
@.dRt�	�5��C�SCB 2q"K o��0�B�T��f�x�����LUTORIAL r"K��O�GV_CON?FIG s"M�A�ZO�OF���OUTP�UT t"I7���R�������̟ ޟ���&�8�J�\� n�4���������̯ޯ ���&�8�J�\�n� �������ȿڿ��� �"�4�F�X�j�{��� �ϲ����������� 0�B�T�f�x߉Ϝ߮� ����������,�>� P�b�t�ߘ����� ������(�:�L�^� p��������������  $6HZl~ ��������  2DVhz�� �����
//./ @/R/d/v/��/�/�/ �/�/�/??*?<?N? `?r?�? �2����?�? �?�?
OO.O@OROdO vO�O�O�/�O�O�O�O __*_<_N_`_r_�_ �_�O�_�_�_�_oo &o8oJo\ono�o�o�o �_�o�o�o�o"4 FXj|���o� �����0�B�T� f�x��������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ����� ����
��.�@�R�d��v߈ߚ߬ߏ8��������Ѷ��? ,�>�P�b�t���� �����������(�:� L�^�p����������� ���� #�6HZ l~������ �2DVhz �������
/ ./@/R/d/v/�/�/ �/�/�/�/�/??)/ <?N?`?r?�?�?�?�? �?�?�?OO%?8OJO \OnO�O�O�O�O�O�O �O�O_!O4_F_X_j_ |_�_�_�_�_�_�_�_ oo/_BoTofoxo�o �o�o�o�o�o�o +o>Pbt����������%���$TX_SCRE�EN 1u����М}i�pnl/Y�gen.htm%�x����������/pPan�el setupČ}�ď��)�;�M�_��鏖����� ̟ޟ�g����8�J� \�n�����	��ȯگ ����"���ǯ��j� |�������Ŀ;��_� ��0�B�T�f�ݿ� �Ϯ���������mϛ� ��>�P�b�t߆ߘ�� ��3�������(�:����(�UALRM_�MSG ?E��R� S�(z����� ���������;�A��r�e�������n�SEoV  |����l�ECFG wvE�O�  (u�@�  A  w B�(t
 �� /sE�Oas����������G�RP 2x 0(v	 9[n��I_BBL_NO�TE y
T?��l/rJ��/q nDEFP�ROx�%|� (%���2p��� / /D///h/S/y/�/�/��/�/�/dFKEYDATA 1zE��Ep (v�HK?]?4?�?�?j:,�(�?�?(t([ ?INST ]�?�>�  ��� ��Z���?�>:OLOE��һ�� e��b�vRO�:[E�DCMD�?�O8@���� Əڂ����O,O�O�O�O#_ 
_G_Y_@_}_d_�_�_��_�_�_�_f>���/frh/gui�/whiteho?me.pngoIo�[omoo�o�"finst4o�o�o�o�o��g  FRH/�FCGTP/wz?cancel�oN `r��%s��������%nex��oS�e�w������d>"fedcmdC�F��ڏ����"�-�#earwrgB�Y�k�}� �����şן���� ���C�U�g�y����� ��>�ӯ���	��-� ��Q�c�u�������:� Ͽ����)�;�ʿ _�qσϕϧϹ�H��� ����%�7�o��m� ߑߣߵ��������� �!�3�E���i�{�� �������d����� /�A�S���w������� ����`���+= Oa������� �n'9K] �������� |/#/5/G/Y/k/� �/�/�/�/�/�/x/? ?1?C?U?g?y??�? �?�?�?�?�?�?O-O�?OQOcOuOl�K}�`����O@�O�M�O�O_�F,�_ 5_�_Y_@_}_�_v_�_ �_�_�_�_o�_1oCo *ogoNo�o�o�o�o�o �o�o	?&c uTߙ����� O�)�;�M�_�q��� �����ˏݏ���� %�7�I�[�m����� ��ǟٟ������3� E�W�i�{������ï կ������/�A�S� e�w�����*���ѿ� ���Ϩ�=�O�a�s� �ϗ�&ϻ�������� �'߶�K�]�o߁ߓ� ��4����������#� ��G�Y�k�}���� ���������1�8� U�g�y���������P� ����	-?��c u����L�� );M�q� ����Z�// %/7/I/�m//�/�/ �/�/�/h/�/?!?3? E?W?�/{?�?�?�?�? �?d?�?OO/OAOSO eO�?�O�O�O�O�O�O rO__+_=_O_a_�O �_�_�_�_�_�_�_����[������o.o@mobotoNf,`�oX�o�o�o �o�o#
GY@} d������� �1��U�<�y���r� ����ӏ���	��-� ?�Q�c�r_�������� ϟ�󟂟�)�;�M� _�q� �������˯ݯ �~��%�7�I�[�m� ������ǿٿ��� ��!�3�E�W�i�{�
� �ϱ���������ߚ� /�A�S�e�w߉�߭� ����������+�=� O�a�s���&���� ��������9�K�]� o�����"��������� ��#��GYk} �������� 1�Ugy�� �>���	//-/ �Q/c/u/�/�/�/�/ L/�/�/??)?;?�/ _?q?�?�?�?�?H?�? �?OO%O7OIO�?mO O�O�O�O�OVO�O�O _!_3_E_�Oi_{_�_ �_�_�_�_d_�_oo /oAoSo�_wo�o�o�o �o�o`o�o+=hOa8 c{�8 ������}����v,Џ�ȏ 9� �]�o�V���z��� ɏ���ԏ�#�
�G� .�k�}�d�����ş�� ������C�U�4 y���������ӯ�o�� 	��-�?�Q�c�򯇿 ������Ͽ�p��� )�;�M�_�ϕϧ� ��������~��%�7� I�[�m��ϑߣߵ��� ����z��!�3�E�W� i�{�
��������� ����/�A�S�e�w� ������������� ��+=Oas� ������' 9K]o��j�� ����/5/G/ Y/k/}/�/�/0/�/�/ �/�/??�/C?U?g? y?�?�?,?�?�?�?�? 	OO-O�?QOcOuO�O �O�O:O�O�O�O__ )_�OM___q_�_�_�_ �_H_�_�_oo%o7o �_[omoo�o�o�oDo �o�o�o!3E�o i{����R� ���/�A��e�w�@��������я�Ӌ���������� ���B�T�.�, @���8�����͟ߟƟ ��'�9� �]�D��� ��z�����ۯ�ԯ� ��5��Y�k�R���v� ��ſ������1� C�R�g�yϋϝϯ��� ��b���	��-�?�Q� ��u߇ߙ߽߫���^� ����)�;�M�_��� ���������l�� �%�7�I�[������ ����������z�! 3EWi����� ���v/A Sew���� ���/+/=/O/a/ s//�/�/�/�/�/�/ ?ڿ'?9?K?]?o?�? �/�?�?�?�?�?�?O �?5OGOYOkO}O�OO �O�O�O�O�O_�O1_ C_U_g_y_�_�_,_�_ �_�_�_	oo�_?oQo couo�o�o(o�o�o�o �o)�oM_q ���6���� �%��I�[�m���� ����D�ُ����!� 3�W�i�{������� @�՟�����/�A��0C��0���l�~���h���į��,������� � =�O�6�s�Z������� Ϳ�����'��K� ]�Dρ�hϥό����� ������#�5�?Y�k� }ߏߡ߳������� ��1�C���g�y�� �����P�����	�� -�?���c�u������� ����^���); M��q����� Z�%7I[ ������h �/!/3/E/W/�{/ �/�/�/�/�/�/v/? ?/?A?S?e?�/�?�? �?�?�?�?r?OO+O =OOOaOsOJߗO�O�O �O�O�O�?_'_9_K_ ]_o_�__�_�_�_�_ �_�_�_#o5oGoYoko }oo�o�o�o�o�o�o �o1CUgy� �����	�� -�?�Q�c�u�����(� ��Ϗ������;� M�_�q�����$���˟ ݟ���%���I�[� m������2�ǯٯ� ���!���E�W�i�{�Ѝ������@���>�@���ܿ�  �ؿ"�4��, �e� ߉�pϭϿϦ����� �� �=�$�a�s�Z� ��~߻��ߴ������ ��9�K�2�o�V��� �O���������#�2� G�Y�k�}�������B� ������1��U gy���>�� �	-?�cu ����L��/ /)/;/�_/q/�/�/ �/�/�/Z/�/??%? 7?I?�/m??�?�?�? �?V?�?�?O!O3OEO WO�?{O�O�O�O�O�O dO�O__/_A_S_�O w_�_�_�_�_�_�_�� oo+o=oOoaoh_�o �o�o�o�o�o�o�o '9K]o�o�� ����|�#�5� G�Y�k�}������ŏ ׏������1�C�U� g�y��������ӟ� ��	���-�?�Q�c�u� �������ϯ��� ��)�;�M�_�q����� $���˿ݿ��Ϣ� 7�I�[�m�ϑ� ϵπ���������!��P�#���P���L�^�p�Hߒߤ�~�,���߈������/� �S�:�w��p��� ���������+�=�$� a�H���l��������� ���_9K]o ���Ϸ���� #�GYk}� �0����// �C/U/g/y/�/�/�/ >/�/�/�/	??-?�/ Q?c?u?�?�?�?:?�? �?�?OO)O;O�?_O qO�O�O�O�OHO�O�O __%_7_�O[_m__ �_�_�_�_V_�_�_o !o3oEo�_io{o�o�o �o�oRo�o�o/ AS*w���� ��o���+�=�O� a����������͏ߏ n���'�9�K�]�� ��������ɟ۟�|� �#�5�G�Y�k����� ����ůׯ�x��� 1�C�U�g�y������ ��ӿ������-�?� Q�c�u�ϙϫϽ��� ����ߔ�)�;�M�_� q߃�ߧ߹������� ��%�7�I�[�m�ﴑ�hp���hp��������������, E���i� P��������������� ��AS:w^ ������� +O6s�d� ����/�'/9/ K/]/o/�/�/"/�/�/ �/�/�/?�/5?G?Y? k?}?�??�?�?�?�? �?OO�?COUOgOyO �O�O,O�O�O�O�O	_ _�O?_Q_c_u_�_�_ �_:_�_�_�_oo)o �_Mo_oqo�o�o�o6o �o�o�o%7�o [m���D� ���!�3��W�i� {�������Ï���� ��/�A�H�e�w��� ������џ`����� +�=�O�ޟs������� ��ͯ\����'�9� K�]�쯁�������ɿ ۿj����#�5�G�Y� �}Ϗϡϳ������� x���1�C�U�g��� �ߝ߯�������t�	� �-�?�Q�c�u��� �����������)� ;�M�_�q� ���������������$UI�_INUSER � ���"��  �_MENHI�ST 1{"  (/ �ڀ)/SOFT�PART/GEN�LINK?cur�rent=men�upage,1133,1A����({�5�5GHYk��'�8%�����~��2$5�B/T/f/�/�71�6w/�/�/��/��,�/�edi�t�DEFAUL=T�PICK�Q?�c?u?��z ?HOME@0ON_<?�?�?��?��<�?!>IPL�_FANUC_S�MPLGRP_CLOS�1SOeOwO�L����v�A�O�O�O�O�O�O_ �O6_H_ Z_l_~_�__�_�_�_ �_�_o�_2oDoVoho zo�o�o-o�o�o�o�o 
�o@Rdv� �)������ *��N�`�r������� �Ȍޏ����&�8� ;�\�n���������E� ڟ����"�4�ßX� j�|�������įS�� ����0�B�ѯf�x� ��������O����� �,�>�P�߿tφϘ� �ϼ��Ϲ�����(� :�L�^�aςߔߦ߸� ����k� ��$�6�H� Z���k�������� ��y�� �2�D�V�h� �������������u� ��.@Rdv �������ύ *<N`r��� ����/�&/8/ J/\/n/�/�/!/�/�/ �/�/�/?�/4?F?X? j?|?�??�?�?�?�? �?OO�?BOTOfOxO �O�O+O�O�O�O�O_�_�$UI_P�ANEDATA �1}���KQ�  	��}  ttp:/�/127.0hP1�:3080/fr�h/jcgtp/�flexdev.�stm?_wid�th=0 &_l�ines=15&�_columns�=40&_fon�t=24&_pa�ge=whole��P'_)  rim�_�_  \P
oo .o@oRodo�_vo�o�o �o�o�o�o�o�o< N5rY������ �  }�p%#t\o 	��-�?�Q�c���� �_����Ϗ���l� )�;�"�_�F�����|� ����ݟ�֟���7�I�0�m��y��MS�� ����ѯ����Z�+� ��O�a�s�������� Ϳ߿ƿ��'�9� � ]�Dρ�hϥϷϞ��� ����߄���G�Y�k� }ߏߡ�����8����� ��1�C�U��y�`� ������������� -��Q�8�u���n��� �0�����); ��_q�ߕ��� ��V�7I0 mT������ ��!//E/����� �/�/�/�/�/�/:/? ~/?A?S?e?w?�?�/ �?�?�?�?�?OO O =O$OaOHO�O�O~O�O �O�O�Od/v/'_9_K_ ]_o_�_�O�_?�_�_ �_�_o#o5o�_Yo@o }odo�o�o�o�o�o�o �o1UgN� �O_����	�� n?�Q��_u������� ��Ϗ6��ڏ�)�� M�4�q���j�����˟�ݟğ��%���}�6�o���������ɯ)]��a�ݯ�,�>� P�b�t�ۯ������� ���ٿ���:�L�3� p�WϔϦύ���Z��s��{�$UI_PO�STYPE  ��u� 	� ��-���QUI�CKMEN  ���0���RESTORE 1~�u�  ���a��ߴӢ�a�m������1�C� ��g�y����R��� ����	����(�:�L� �����������r��� );M��q� ���d����\ %7I[m�� ���|�/!/3/ E/��d/v/��/�/ �/�/�/?�//?A?S? e?w??�?�?�?�?�? �/�?OO�?OOaOsO �O�O:O�O�O�O�O_ _�O9_K_]_o_�_;�oSCREK�?P�u1sc��Wu2�T3�T4�TU5�T6�T7�T8�Q�STAT�� x_Ӵu��USER�P��_�RTPSC�Sk�s�SWd4Wd5Wd6�Wd7Wd8Wa��ND�O_CFG ��F�E���OP_C?RM5  A��f���PD�Q9i�?None>�0`�_INFO 2�j�up]�0%�_ Z�
K.o�d ���������5�G�*�k�4��aOFFSET ��qx�"S��*_��Ώ �����(�U�L�^� ��b��������ܟ� ��$�6���`߂�p����
��ʯV�a�aW�ORK ��m�������z�/`UF�RAME�o�RTOL_ABRTi���c��ENB��{�G�RP 1���\�?Cz  A��ޱ�"Q޿���&�8�B�T�y�J�U���a��?MSK  ��qڙ�Nf�%�i�%xR��ϛ�_EVN��b���f֑b3����
 h�aUE�V��!td:\�event_usger\��M�C7R�d���`F׭F�SPK��P�spotwe{ld��!C6���ߚ߾P��!��a�� T��ו��C�1��� g�y����������� ^�	���-�?�u����� ��������6%Z �;��q���� ��
"�W�3�:i��8�� r����/� '/9//]/o/J/�/�/ �/�/�/�/�/?�/5?�G?"?X?}?�?�$V�ALD_CPC {2��� k?�?�a O��Q<�@*�O7OIO��"S&BdpJm@j��IlD[�O V�?�O�?�?_O/_ A_S_bOtO�O�O�_�O �_�O�O(_oo=oOo ^_p_�_�_�_�_�o�o �_ o$o9K�olo ~o�o�o]�o��o�o � �G�Y�hz� ���׏b��
�� .�C�U�d�v������� ��Џ����*�+� Q�c�r���������̟ ����)�8�M�_� n���������˿گ� ���%�4�I�[�m�|� ����Fϴ�ֿ����� �3�B�W�i�xϊϜ� ������������/� >�S�e�w�ߘߪ߼� ��������L�=�,� a�s���������� ���$�9H�]o ������������  �D6k}� ������� .C/Rg/y/��� ���/�	?/*/? N/O?u?�?�/�/�/�/ �?�/O?&?8?MO\? qO�O�?�?�?�?�?�O �?_"O4OI_XOm__ �_�O�O�Oj_�_�Oo _0_B_Wof_{o�o�_ �_�_�_�_�oo,o >oSbow���o�o �o�o��(:p a�P��������� � ��'�6�H�]�l� ����*���Ə؏ꏥ� �#�2�D���h�Z��� ����ԟ����
�� ��@�R�g�v������� ��Я���	��-�<� N�5�r�sϙϫϺ�̿ ޿����)�8�J�\� q߀ϕߧ߶������� ���"�7�F�X�m�|� ���������ߎ��� �3�B�T�f�{���� �����������,� AP�b�w����� ������(=L ^��t���� � $&/K/Zl �/��/�/N/��� /�/2/G?V/h/"?�/ ~?�?�?�/�/�/??�.;�$VARS_�CONFIG �i0PA�  FP53��4LCMR_GRPw 2�PK�8��1	a0\@  %�1: SC130EF2 *�O�@54ə.5i0��8�0�5�`0`1?�  A�@�@p
@�.N 	&OX_.8<_N_�{_�Av_�_UA��@�Q�52�_�_52 B����Q 51�U�_ og_Dooho So�owo�o�o�o�o=o �oRov��<DIA_WORKW �PE�pz0�6,		j1PE�>�wG�P ��pY9��qRTSYNCS_ET  PI�PA��WINURL 3?�b0��X��j�|��������vSI?ONTMOU�53�<� �ʅ_C�FG �S۳�S۵PZ@� FR:\̃\�DATA\�� �� UD1�wLOG�  1��EX=�51' ?B@ ���P��=?��P���ş.7 �� n6  ���.6|��<���A  =�����54�Q�TRAIN�f���&� 
�7p��v�]4#��|B�PK (?qg��� 7y����ӯ���-�� Q�?�Y�c�u��������Ĉ_GE�PK�``0�
z0x2�c�RE���PE�8H�LEX�PLa01�-e��VMPHA�SE  PE�3��P=CRTD_FILTER 2�PK ��E�_���� ����,�>�P�b�t� .7�Ϣߴ����������� �2�D�7ISHI�FTMENU 1��PK
 <k<%����݂������� ���������K�"�4� Z���j�|������������	LIVE/�SNA`C%vs�flive���̃ �U`@4menuJO������r`��5�Y�MO��Q��@@@ZD���.�51<Y��P��$WAITDINEND׈`1�HOK  �IcՊr~S�eTIMׅ���GO�q�+�����cRELE|�'�Hҏ<�J_ACT' (t�qc_� ��y��%�?9F�"RD�IS`@�.�$X�VR��Q��$oZABC{B1�+' ,Y�Bu2?2M�!� VSPT q�Q͚E�
�
���?�
�?O�7D�CSCHG ���{�@�04GBph0IP$�+A�O�O��O�:MPCF_G' 1��IA�0�7,_�OMPn3��I���p���?o_=���  3~� ��w�?����vԿ�P�R����~�lD&t�����D)���?^U�����Q�w@t_�W� �U��]��X�]�S �_�Y
i�Vo<o^_�o��e�Y´ ²�E�³��l�*�`��b��k��P�o �o&P{�_�_�_��R0�_8od4�@�����O�t_CYLINuD����K �}f ,(  *��&���O�6�s�Z� �o����͎���_� ����J���n����� Տ��Q�7��ӟ��� e�F�X��|����G�! �_�����3�o�ܯǯ �婓�0�姖�J�A��tSPHE_RE 2��}̪� ����������(�;� �(Ϥ�L��ѿ��i� �ύ�������5�G�$� ��H�/�A�~��Ϣߴ�l��h0ZZ�& ��