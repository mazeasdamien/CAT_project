��   v��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@���&�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	>4SUSRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  wXKaIRTs1�	o`'2 L1���L2�R�	 %,��?���b1`Q�c�c~a����? � �`�c<�o��
 ��a�o@�o1CU �o z�����c� 
��.�@�R��v��� ������Џ�q��� *�<�N�`������ ��̟ޟm���&�8� J�\�n���������ȯ گ�{��"�4�F�X� j���������Ŀֿ����`TPT�X��ʊ�)�� �s �Ƅ�$/�softpart�/genlink�?help=/m�d/tpmenu.dg���ϨϺ���r��&a�s�pwd�� �+�=�O߄�s߅ߗ� �߻���\�����'� 9�K����߁����X�������a�f9�b�� ($p�-�@���T�?�x���a��a��c���c����Dl��k
���a�ah�a�ah��h�	.f���������q�`���`  ���|f ep��Jh#h�F�bc Xc�B 1)hR �\�`_�� �REG VE�D]���who�lemod.ht}m�	singl	�doub �trip8browsQ��� ��u���//�@/���dev�.sl�/3� 1�,	t�/_�/;/i/ ??/?�/S?e?w?�?�?�?� ��?�? OO%O7OIO[OmOO�E @�?�O�O�O�O �O_�F�	�?�?;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo oM'�o�o�o�o�o�o +=Oas� ��������? >�P�b�t��������� Ώ���O�����L� ^�_'_�������ş �����6�1�C�U� ~�y�����Ư��ӯ�o ���-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�-��Ϭ� ����������*�<� 7�`�r�A�Sߨߺ�q� ��i�����!�J�E� W�i��������� ����"��/���O�I� w��������������� +=Oas� ������, >Pbt���߼ ���//����� ^/Y/k/}/�/�/�/�/ �/�/�/?6?1?C?U? ~?y?�?Y��?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _�R_d_v_�_�_�_ �_�_�_�_�o*o�_�o`oro�j�$UI�_TOPMENU� 1K`�aR 
d�a�*Q)*defa�ult5_]*�level0 * [	 �o�0��o'rtpio�[23]�8tpst[1[x)w9��o	�=h58E�01_l.png���6menu5�y�p�13�z��zb	�4���q��]� ��������̏ޏ)Rr����+�=�O�a����prim=�pa�ge,1422,1h�����şן����1�C�U�g����|�class,5�p�����ɯۯ�����13��*�<�N�`�4r���|�53�������ҿ�����|�8 ��1�C�U�g�y�����@����������"Y�` �a�o/��m!ηq�Y��w�avtyl}Tfqm�f[0nl�	��c�[164[w��59@[x�qG���/��29� �o�%�1���{��m� �!�����0�B��� f�x���������O������,>����2 P�����\�� '9K�������������1���/$/6/H/Z/��~|�ainedi'���/�/�/�/�/��c�onfig=si�ngle&|�wintp���/$?6?H?�Z?	�ߐ??ٷ�gl�[�<��?�߲08@��
A���?,OH2�ڀDO�?cO�O�z �� �4s�x�O�O� $��Ol�E_W_i_{_�_ �_���_�_�_�_oo /o�_Soeowo�o�o�oz�$;�$doub5�o��13��&du�al�i38��,4�o&�o9�o�n�o �a8���Ao�� ��&�8��\�n��� ������m�����
� �.�@�K�d�v���������Z{?�;�M� sc�_;���s��X�}���e�u��0�����O_ �J�p�^�6e�u7�����ｿϿ ���P�)�;�M�_� qσ�ϧϹ�������(���"�1�M� _�q߃ߕߠϹ����� �����7�I�[�m� �������������!�����6(�]�o�`�������$��74��@����)�C�ߟ�T�	TPTX[c20�=Aw24#GJ���Bw1H�� ����8�"H���A0#��[�tv`�R���@2�K0�1�1���5S:�$tr?eeview3�f�3��o}381,26M/_/q/0�/�/ �/�/�/�/~/?%?7?@I?[?m?�o/܈5�o 5%���?�?�?
?#O5O�GOYOkO}O�?�? "2�?8"2K��O�O_�O��1�?�E�f_x_�_� �6_ڀedit�a>_P_�_�_oˉ /���_�Cooo�o�o B�o�o��oA�o� +=Oas� �o������� (�9���Q�x������� ��ҏO����,�>� P�ߏt���������Ο ]�����(�:�L�^� ퟂ�������ʯܯk�  ��$�6�H�Z��l� ������ƿؿ�y��  �2�D�V�h����Ϟ� �������ϕo�o��o @ߧE�c�u߇ߙ߬� ������O����)�<� M�_�q���W����� ����&�8���\�n� ��������E������� "4��Xj|� ���S�� 0B�fx��� �O��//,/>/ P/�t/�/�/�/�/�/ ]/�/??(?:?L?�� ߂?1ߦ?���?�? �?�?O$O5OGO�?SO }O�O�O�O�O�O�O�O ��2_D_V_h_z_�_�_ �/�_�_�_�_
oo�_ @oRodovo�o�o)o�o �o�o�o*�oN `r���7�� ���&��J�\�n� ��������E�ڏ��� �"�4�ÏX�j�|��� ����a?s?蟗?�sO _/�A�S�e�w����� ����������,� =�O�a�#_������ο ��=��(�:�L�^� pς�Ϧϸ�������  ߏ�$�6�H�Z�l�~� ߐߴ���������� ��2�D�V�h�z��� ����������
���� @�R�d�v�����)����������ƚԔ�*default�%��*level8�ٯw���?� tpst[�1]�	�y�t?pio[23����u���J\�menu7_l.�png_|13���5�{�y4�u6���//'/ 9/K/]/���/�/�/�/ �/�/j/�/?#?5?G?�Y?k?�"prim�=|page,74,1p?�?�?�?�?��?�"�6class,13�?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_�B_T_f_x_{?�218 �?�_�_�_�_�__B6o9oKo]ooo�o`��$UI_USE�RVIEW 1�֑֑R 
���o��o�o[m�o'9K ] �����l ���#�5��oB�T� f������ŏ׏鏌� ��1�C�U�g�
��� ������ӟ~����� v�?�Q�c�u���*��� ��ϯ�󯖯�)�;� M�_�
��~������ ݿ���%�ȿI�[� m�ϑ�4ϵ������� �Ϩ�
��.ߠ�i�{� �ߟ߱�T�������� �/���S�e�w��� Fߨ����>���+� =�O���s��������� ^�����'���� FX��|���� ��#5GY� }����p�� �h1/C/U/g/y// �/�/�/�/�/�/�/? -???Q?c?/p?�?�? ?�?�?�?OO�?;O MO_OqO�O&O�O�O�O �O�O�?�O_ _�OD_ m__�_�_�_X_�_�_ �_o!o�_EoWoio{o �o0h