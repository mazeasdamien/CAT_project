��   :�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����FSAC_L�ST_T   �8 $CLNT�_NAME �!$IP_ADD�RESSB $A�CCN _LVL  $APPP � ���$8 A~O  ���z�����o VER�SIONw�  XK�IRTUALw�'�DEF\ � � �� ���ENA'BLE� �������LIST 1 ��  @!ȁ,��)���� (yL^���� ���-/ /Q/$/u/ H/Z/�/~/�/�/�/�/ �/?�/:? ?q?D?V? h?�?�?�?�?�?O�? 7O
OOmO@O�OdO�O �O�O�O�O_�O3__ _T_<_z_`_�_�_�_ �_�_�_�W