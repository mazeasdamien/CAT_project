��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  � QA> �1
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1�TU4QQER�AR�x1R� � /$TIT91� �� � �Td�T0�ThP�TU5�V6�V7�V8�V9�W0�W�WOQ�U�W�gQ�U�W1�W1�W1��W1�W2�R!SBoN_CF�!@$<!J� ; ;2�1�_CMNT�$�FLAGS]�C�HEK"$�b_O�PTJB � ELL�SETUP � `@HO8@9 P�R�1%�c#�aREPR�hu0D+�@���b{uHM9 MN��B;1��AUT�OBJ U��0 49DEVIMC�STI/@�� ��@b3�4pB�d�"V�AL�#ISP_UsNI�tp_DOcv<7�yFR_F�@|%�u13��A0s�C_�WA�t,q�zOFFu_T@N�DEL��Lw0dq�1�Vr?1^q�#S?�o`Qb"U�t#*�QTB����MO� �E' � [M������REV�BI�L���XI� v�R_  !D�`~��$NOc`�M�|��0��ɂ/�#ǆ� ԅ��!X��@Ded p �E RD_E��h��$FSSB6�`K�BD_SE�uAG*� G�2Q"_��2b�� V!�k5p`(��C��@0q_ED� �� � t2�$!SL�p-D%$� �#r�B�ʀ_OK1��0] P_C� ʑ0tx��U �`LACI�!��a�Y�� �qCOsMM� # $D
�� ��@���J_\R_M��BIGALLOW� (Ku2-B�@VAR���!�AƮ#BL�@� � !,K�q���`S�p�@�M_O]˥��CCFS_UT��0 "�A�Cp'��+pqXG��b�0 4� OIMCM ��#S�p �9���i �_�"tO?  ��M�1� h$�IMPEE_F�s��s��0� t����D_���J��D��F����q_����0 T@L��L�DI�s@G�^� �Pć$I�'���Fned X@GRU@���Mb�NFLIx�\Ì@UIRE�xi42� SWITn$�`0_N�`S 2CFz�0M� �#u�D��!��v`���J�`J�tV��[ E���.p�`�ʗELBOF� �շ�p@`0���3����� F�2�T��A`�rq1J1,��z _To!��pЩ�g���G� }�r0WARNM�p�#tC�v`�ç` � C�OR-UrFLT�R��TRAT9 T|%p� $ACCVq���� ��r$OR�I�_&�RT��S\<��@CHG�0I�E��TW��A�I'��T�m�D���� �202�a1��HSDR�2��2�2J; �S���3��4��5���6��7��8��9�KD׀
 �2 @.� TRQ�$vf��4'�1�<�_U<�G�z�Oec  <� �P�b�t�53>B_�LL�EC��!~�MULTI�4�"u�Q;2ПCHILD��;1 t_��@T� "'�STY92	r��=���)2���ױ��ec# |r056$J ���`���uTOt���E^	EXTt�����2��22"(�0����$`@D	��`&��+����� %�"��`%�ak����N�s��?���&'�E�Au��Mw�9 ��% ��TR�� ' L@U#9 ����At�$JOB`����PM�}IG��( dp������^'#j�~�x�pO�R�) t$�F�L�
RNG%Q@�TBAΰ �v&r�*`1�t(��0 �x!�0�+P��p�%���*��@͐U��q�!�;2J�S_R��>�C<J�T8&<J D`5CF9����x"�@?��P_�p�7p+ \@RaO"pF�0��IT�s�0NOM��>Ҹ4s(�2�� @U<PPgў�P8,|Pn��0�1P�9�͗ RA���pl�?C�� �
$TͰ.tMD3�0T��pQU�`�΀+AHlr>�T1�JE�1\�J����PQ��\Q��hQCY�NT�P��PDBG�D̰�0-���PU�6$$Po�|�u�AX�����TAI�sB�UF,�\��B�1. �����F�`PI|�U-@PvWMuXM�Y��@�VFvWSIMQ�STO�q$KEE�SPA��  ?B�BP>C�B�A��/�`�ˏMARG�u2�F�ACq�>�SLEW *1!0����
�4s��CW$0'���pJqB�Ї�qDECj��e�s�V%1 �Ħ�CHNR�MP�s�$G_@�gD�_x�@s��1_FP�5�@TC�fFӓC�Й���qC��+�VK�*��"�*�JRx���SEG�FR$`IOh!�0S�TN�LIN>�csPAVZ�z�Ц@�D2�� ��r 2��hr�rWQ��?3` +^?�� �եq�`��q|`����p�t��|aSIZ#�!� �T�_@%�I��qRS�*s��2y {�Ip{�pTpLF�@��`��CRC����CCTѲ�Ipڈ�a���b��MIN��a1�T����D<iC �C/����!uc�OP4�n j�E�Vj���F��_!uF��N����|a��=h?KeNLA�C2�AOVSCA�@A�U�r1�4�  �cSF�$�;�Ir ��3�a�05��	 D-Oo%g��,,m�P���ޟ� VQRC�6� n���s���U��R�0HANC��$LG��ɑDQ�$t�NDɖ��AR۰N��aqg��ѫ�X�ME��^�Y�[PS�3RAg�X�AZ�П�t��rEOB�FCT��A��`�2t!Sh`0ADI��O��y�s"y��n!�������~#C�G83t!��BMPmt@�qY�3�afAES$�삓��W_;�BAS~#XYZWPR��R*�m!��	�I7_7  ƀI@dd���8\�p_C:T8���#�cR_L
 � �9 ���C�/�,(zJ�LB�$�3��D��5�FORC��b�_AV;�MOIM*�q�SaԫBP`�@��y�HBP�ɀE�F��~��AYLOAD&$ER�t&3�2��Xrp�!*z�R_F}D�� : T`�I�Y3��E�&��Clt��MS�PU
a$(kpD��9 �rb�;�B�	EVId��
�!_IDX�$���B@X��X<&�SY5� M�_HOPe�<��ALARM��2W�r��2R_�0= h�b P�q�`M\qJ@�$PL`A&�M#�$�`��� 8�	���V�T]�0�VQU�PM{�uU��>�TITu��
%�![q�BZ�_;���? �B �pQk��6NO_HEADE^az��}ѯ� �`􂳃���dF�ق�t� ���@�@��uCIRTR�`��ڈ�L��D�CB@4�RJ`��� \P���A�2L>���OR�r��O��<��F`UN_OO�Ҁ$����T������I�VaCx�PX�WOY���B�p$�SKADR�DBT��TRL��C���րfpbDs��~�DJ$j4 _�DQ}�։PL�qwbWA����WcD�A��A�=�2�UMMY9���10�~pDBd����D;[QPR��? 
9�D�Z����E O�Y1$��a$8��L�)F!/�2����0G�G/���PC�1H�f/�PENEA@T�f�I�/Y#�REC�OR`"JH �@ �E$L�#F$#PR���+jp���q��_D$�qPROSS]�
���R�r�` u�$TRIG96P�AUS73ltETU�RN72�MR:�U2 0Ł0EW$��?SIGNALA�QR�$LA�З5�1G{$PD�H$Pİ"�AI�0�A�C�4�C��DO�D�2�!��6GO_AWAYF2MOZq�Z�� {CS��CSCBg��K Իa#���ERI�0Nn�T�`$������FCBPL�@QBGAGE���P��ED|B0D�wA[CD�OF�q[F�0�FoC��MPMA�B0XoC�$FRC�IN��2Dk��@���$NE�@�FDL|8�� L� ��@��=��Rw�_��P� OVR10���l�~��$ESC_�`>uDSBIO����pTe�E�VIB�� �`s��Z��V��pScSW��$�VL�:�Lk��X���ѣ�bQ�����USC�P��A8=�	Q��MP1%e&S�*`�(bt`'c5۳ESUd��-cWg&SWg ?cWd����Wd��Wd.���AUTO$�Ya҃�ac�SB����-d���&SwB[��GB�f$/VOLT�g ��  �GAOD!�qr���@:�ORQҀ�Kra�$DH_THE&0�Rgp� qtnwALPHnt��o���w0 Vp]�$�.�R a�[��s�5�`r�CQ#RBUD�S� F1M�B�sV
��;��Lb��tk���BRTHR���L��T`�Z���Vɖ��DE  �1��2�⋅�� ������kѯ�aәT t0V�ꆸ������̈ Я�-�"�N~��sxS2����INHB��ILTG0ɡ�T?��3 $�w��E��PqQxQ�ThqPe��0Y�AF}�O�ນ��ڗ�� qPڳē����bPܙ����PL?���3���TMOU��ēS���� ���s�/�S18���O�A�ܙ��I����CDI8Ƒ˩o�STI��գ��O:ҋ�,0���AN��Qg�S��+r��#x$�����w�_�����PRA�P`pvC����MCNeQ�e�����VERSP��r�oPIw�FP�åǲШ۷G.�DN"��G>�����F�2ŤǷ�M�7�F��_
�MN�D̠,����d �{ƭa����OB��`�U˱z���DI�� ��#���3�����A����w�Fx���3�ONp�5��Q��VAL�{CR[�_SIZ��8b�;Qn�REQ�Rb�`�=2b���CHq� ΂�ڃ�Ռ�����:��n�S_U��X��wWF�LG���wU$�CV�iMGP�QδFLXP�923R�u���&EAL�P-�C	��
+rT��W��� �R�cx���NDMS7�d ��K>S�P_M'0h�STWv�������AL�P���Q���pU���U�IAG,��o��d�U�-�T"A-`� ���A������H`��Q`��6��Pq_D&��1s��.�P��F�>2�T�� ?7 1A>��#�t#L��?_0=i @@>LD�cง�0�FRI�0 �`Ѐ��1}ѲI�V\1�*�>1�UP�`��a��C�LW��
`L=S&-c&&S�C.w�� L����!����d�Q$w�҇��$w���8�
�P�5RSM��(�V0h � r��d6^2AW�a_TRp}��8@NS_PEA�����< ��$�SAV�G�8�6G]%���CAR �`�!�$���"�CRa���$ d�#E8�@��"STD���!qFpo��'QOF���%��"RC���&RC۠�(F�2A�R#7��X�%, gMA�Q_�a���
QQ��al2��u4Ib�r7I�R�9wQH�7�8M/��!Cp�R�  �p�2F�<�SDN�a0 0�2W2QM P $Mi��s$cA� $C�cm�9���4�A�T�0CY_ wN LS!IG1x'�yB��y@@H2Y�N�O����SDEV�I�@ O@$n�RBT:VSP�3�CuT�DBY|�A	W|`3CHNDGDAwP H@GRP�H	E iXL�U��VS�F�x2� CL1p aQ6ROp��FB�\]�FEN�@��S���ChAR d�@DyOd�PMCSb���P薇P�R��HOT�SWz42�DMpEL�E�1/ex\8`�RS T�@���r� hf��`OL�GHA�Fk�Fs��C�A@T � $MDLUb/ 2S@�E���q��6�q	0�i�c�e�cJ��	uݢ�#~5t+w�PTO��� �byUހTSLAVS� wU  ��INP ��	V�ЊyA_;�EN�UAV $R�PC�_�q�2 1bL�w�aD�pSHO+� �W ���A�a�q�2кr�v�u�v�sCF�� X` ,f��r�OG gE��%XD�h��pC�Iߣ�i�MA��D�x AYr?�W� p�NTV	��D�VE�0@�SKIB��T�`g?Ň2��" JZs�! Cꆻ���f�_SV/ �`X�CLU��H���O�NL��'�Y�T��O=T:eHI_V,11 �APPLY��HI�4`;�U�_ML�� $VRFY8��	�U�M{IOC_�I���J 1/��߃O��@X�LSw"`@$?DUMMY4����ڑ�Cd L_TP����kC��^1CNF f���E��@T�y� 	D_#UQ_��ݥ�YPCP��=�� �����G�?$����џ Y +�
0R�T_;P�~T��C�Cb Z�r�TE ���=�פ�DG�@�[ D�P_BA�e`kc�!$��_��H���\�� \�pAb�=cARGI�!$����`[���c_SGNA] ��`U���IGN�Տ��� ���V������ANNUN��&�˳�EU�<J'�ATCH���J��y��t^ <`@g�����:c$Va������ᑴaE�F] I�� _ �@@FͲITb�	$TOTi �C�O��c�c@EM�@NIF�a`tB��c��ùA>���DAY@CLOAD�D\�n���� �EF7�X�I�Ra��K���O�%��a?�ADJ_)R�!@b��>�H2��"[�
 c�%��`a�͠MPI�J��D��qA��?�Ac 0� �х�� ��Z�ϡ��Ui ��CTRLܖ Yp d��TR�A8 ?3IDLE_�PW  �Ѡ��Q��V��GV_���`c ��o�;Q@e� �1$��6`<cTAC�-3��P�LQ�Z�Rdz\ A-u:ɰSW;�A\���/Jղ�`b�K�OH�(OsPP; �#IRO� ��"BRK��#AB  �O������� _ ���F���`d͠, j@�S�RQDW��MS��P6X�'z��IF�ECAL�� 10^tN��V��豊�V�(0}f�CP
��Nr� Yb�0FLA_#f�OVL ��HE��>�"SUPPO��ޑ�\�L�p��&2XT�$Y-
Z-
W-
���/��0GR�XZl�q�$Y2�CO�PJ�SA�X2R��*r�!���:��"!�I�0)��f `�@CACH�E��c��0�s0L}AZ SUFFI, C��q\��哹6oÀPMSW�g� 8�KEYIM[AG#TM�@S�àn
2j�r���aO�CVIE��~�h �aBGL����`�C?�@��P���i��m!`STπ!� ���������/EMAI�`N��`A��PZ�FAU� �jH�"�qa��U�3���� }�k< �$I#�US�� �IT'�BUF`�r�DNB���SUBu$��DC_���J"��"SAV�%�"k�������';��P�$�UOR	D��UP_u �%��8OTT��_B`��8@�LMl�F4��C7AX�@Cv���Xu 	��#_uG��
�@YN_��R�l6���D�E��UM����T��F���caC�DI`BED%T)@C��~�m�rI��G�!c�&��l`����Q�P��FZP n (�pSV� )d\��ρ��-�A��o�� ����>"$3C_R�IK��kB���hD{pRfgE.(AD�SP~KBP�`�II�M�#�C�Aa�A��UЂG���iCM! IP`��KC��� �DTH� ȷS�B*�T��CHS�3�CBSC��� ���V�dYVSP�#[T_D^rcCONV�Grc�[T� �Fu F�ቐd0�C�0j1��SC5�e�]CMER;dAFBgCMP;c@ETBc� p\FU D�Ui ��+�~�C�D�I%P702# �E	O���qWӏ�SQ��1QǀSU��MSS�1j�u�4`�T�aAa��A>�1r� "�Й��4$ZO@s���"l�U6�&��eP���e�CNc�l��l�l�iGGROU�W)��S c�MN�kNu�eNu�e NpR|b|�i�cH�pi�8�z
 �0CYC���s`�w�c��zDEL�3_D��RO�a�� �qVf���v{�O�2� ��1��t��:R�ua�.#�� ��AL� �1s@ˢI1¡�J0�PB��,���0ER^�T�Gbt ,!@��5��aG�I1LcR1s 
M!A������1u����H�����P����Cڠ	������2��J0��0vH *	�L U�1#J�Q��V
�[�7A z���z��z��z�Ѩz�Fz�7w�8w�9Pw���y���1��1��U1��1��1Ě1њU1ޚ1�2��2�����2��2��2��2�Ě2њ2ޚ2�3J��3��3����3��U3��3Ě3њ3ޚe3�4��BXTF��1w6�.(�0�f�0�U�0ŷ�e��FDR�5�xTU VE���?1���SR��REr�F���OVM~Cz)�A2�TROV2ɳDT� R�MXa�I�N2���Q�2�IND�p�r�
���0�0�0G@u1��[�G`��{�D_֎[�RIV�P��G�EAR~AIOr�K"N�0�y�p�5`�@�a�Z_MCM܀ �� �F��UR��Ryǀ��!?� ��p?nЋ�?n�ER�vёa�!��P��zI:�PXq�B�RI0%�ԩ�UP?2_ { ���##TDPR�%TBp������Վ��C�2| QT��"�4)�:%	`t^B��p�IFI���� Mc���.�PT���!FLUI��} � ��K UR �c!���B�1SPx E��EMP�p�2$��S.^�?x��Jق0�
3VRT���0x$�SHO��Lq�6 A�SScP=1��PӴBG_���-���x���FORC3"��i�d~)"FUY�1�2\�2�1�h�ܦ p� |��NAMV�a��������S!"��$VIS�I��#�SCM4SEP����:0E�V�O���$���M���$�I��@�F�MR2��� �5`�r�@ǀ� �2�I�9 F�"�_����LIMITy_1�dC_LM��|����DGCLF��6��DY�LD����!5�������M�Fc����u	 T�sFS0Ed� P���QC�0$EX_QhQ1i0�P�aQ53�5��GoQ��g� ����RSW�%�ON�PX�EBUG���'�GRBp�@U��SBK)qO1L� ��POY 
)�(�P��M��OXta`SM��E�"�a���`_E � �0�F���TERMZ%��c%=aORI�1_ �~c%me�SMepiO��_ �|'��`��(�c%�UP>� ?�� -���b����q#� ���G<�*� ELTOQ�p�0�PFIrc�1Y���P�$�$�$UFR�$��1L0e&� OTY7�PT4q��k3NST�pPATz�q4PTHJ�a�`EG`*C�p1AR�T� !5� y2$2R�EL�:)ASHFTPR1�1�8_��R�P�c�& � $�'@�@� ��s�1 @I�0�U�R G�PAY�LO�@�qDYN_�k���.b�1|��'PERV��RA��H��g7��p�2�J�E-�J�R�C���ASYMFgLTR�1WJ*7����E�ӱ1�I��aUT�pbA�5�F�5aP�PlC�Q1FOR�p�M�I!����W��/&�0F0�aels�H��Ed� �m2XN���5`OC1!>?�$OP�����c�����bRE�PR.3�1a�F��3e��R�5e�X�1>(�e$PWR��_���@R_�S�4��et6$3UD�� �R72w ���$H'�!�`ADDR�fH�L!G�2�a�a�a��R���U�� H��SSC����e-��e���eƪ�SEE���HS{CD��� $����P_�_ B!rP􍀌����HTT�P_��HU�� (�OBJ��b(�Qp��eLEx3Us��� � ���ะ_��T?#�rS�P��z�sKRN�LgHIT܇ 5��P���P�r������PL��PSS<�ҴJ�QUERY_FL�A 1�qB_WEBwSOC���HW��1U���`6PIN'CPU���Oh��q�����d���d����e��IHMI_ED^� T �RH�;?$��FAV� d�~Ł�IOLN
◓ 8��R�@�$SLiR$INoPUT_($
`���P�� CـS�LA� �����5�1��C��B�QI�O6pF_AS7��$L%�}w%�A��\b.1�����T@HYķ�����ah�wUOP4� `y� ґ�f�¤�������`PCC
`����#��>��IP_ME��7� Xy�IP�`�U�_NET�9����Rĳs�)��DS�P(�OqFO�BGȞ�`��M�A��� �l�:CTAjB�pAF TI�-U��Y ޥ��0PSݦBUY IDI�rF ��P������ �y0�,�����Ҥ�NQ�Y R���IRCA�i� ך ěy0�CY�`EA�����񘼀�CC����R�0�A�7Q�DAY_���NTVA����$��5 ����SCAd@��CL���� ������8�Y��2e�o�N_��PCP�q��ⱶ�� ,�N����
�xr����:p�N� 2� !؀��(ᵁ����xr۠LABy1��Y .��UNIR��Ë �ITY듭��e�R�#�5���R_U{RL���$AL0 �EN��ҭ� ;�T��T_U��ABKsY_z��2DISԐ��Al�Jg�����P�$���E��g�R���З A�/���J����FLs��7 Ȁ|���
�UJR� ���F{0G��E7��J7 O^ R$J8I�7�H�R�d�7��E�8{��H�APHIQ�S��DeJ7J8�B��L_KE*� � �K��LM�[� � <X�X�Rl�u���WATCH_VA��o@D�tvOFIELc��cyU L��4� � o1Vx@��-�CT[�9�m�q�LGH��� �$��LG_SIZ��t�z�2y�p�y�FD��Ix���+!��w� \ ����v��S���2 ��p�������\ ���A4�0_gCM]3NzU
RFQ\vv�rd(u�"B��2�p����I ��+ �\ ��v�RS���0  �Z�IPDUƣ�qLN=��ސ�p�z@6���f�>sD�PLMnCDAUiEAFp0���TuGH�RE��|�BOO�a�g� C��I�IT+����`��RE���ScCR� �s��DI���SF0�`RGIO"$D�����T("�t|�	S�s{�W$|�X���JGM^'MNCHL;�|�FN��a&K�'�uЅ)UF�(1@�(F�WD�(HL�)STP�*V�(%Г(��(�RS9HIP�+��C�[T�# R��&p:'^9U =q�$9'�H%C𜓚"Gw)�0PO�7�*�`�#W}$���)EX��TUI�%I���Ï����rCO#C� *�$S��	)��B@v�NOFANA|��Q
�AI|�t:��EDCS��c�C�c�BO�HO�GS���B�H9S�H(IGN�����!O���DDEV6<7LL����-�ҭЦ(�;�T�$@��2�p������#A���(�`�{�Y��PWOS1�U2�U3�Qp	��2�@�Ш ��{�PtD����&q`)��0�d��VSTӐ�R�Yl�\@ ` /�$E.fC.k�p�<p=fPf���4�ѩ LRТ� ��x�c�p���<�Fp�dY�@!�_ � ��7Lpx&���c �MC7�� ���CLD�PӐ��TRQLI0#ѽ�ytFL��,r��5s8�D�5wS�LqD5ut5uORG���91HrCRESERAV���t���t���c~�� � 	u095t5u��PTp���	xq�t�vRCLMC�������q�Y�M��k�������$DEBUGMA�S��ް��?U8$T�@��Ee�g���MFRQՔ� �� j�HRS_KRU��a��A���k5FREQ� �y$/@x�OVER�С�n��V#�P�!EFI�%�a��g�I9���t� \R�ԁ�d�$U�P��?��p�PS�P��	�߃C��͢a��U|\�l�?( 	��MISC� Yd@�QRQ��	��3TB � Ȗ0A�՘AX����ؗ�E�XCESj�5Ъ�M��\��W�����	����SC�P � 	H��̔_��Ƙǰ]�����MKHԳ�K�J� m�B_K�F�LIC�dB�QU�IREG3MO��O�˫3�R�L�`MGմ �`��T����aNDU�]���>��k�G�Df��I�NAUT���RSM>�a��@N�r]3x-�pP4�PSTL\�w� 4X�LOC�V�RI%��UEXɶA�NGuBu��qODA����������MFO����Y�b@p�e4�2k�SUP�evQ�FX��IGG� � ��p�c ���cQ6�dD�%�b|� !`��!`��|��3w�ZW&a�TI�V��XP�IN[�� t��MD��I�)֟@����HݰM��DIA�����W,!�wQt�1�D�)$L밸���]�� 0�C�U��VP��p�<�Or!_V��ѻ ��P0�S�X�5�����ءP��0N���P��KqES2���-$B� ����ND2�����2_TX�dXTR1A�C?�/��M�|q�`�Pv��XҰ�P�t SBq`�USW�CS��T��	���PgULS��A�NSޔ���R��JOIN@��H��~`j�=��b@��b�����P=��0$��b$���TA����S���S�HS�E��S�CF�aPJ��R��P�LQ� 
��L�O��н.���^�	 ��8���������RR2��� �1��eA�q d%$��Iΐ+�G�Ay2+/� �P�RIN�<$R� SW0"�a/�A;BC�D_J%�¡\u��_J3�
�G1SPܠe�u�P�B�3��р`u���J/���r�qO8QI<F��CSKP"zH{�{�J���Q�L2LBҰ_AZ�r�~ELQ��OCMPೕ�T���cRT�����1�+�����P1��>@�Z��SMG0��=�J�G�`SCL�͵S'PH_�@��%V�zu� RTER` � �< A_�@G1�"�A�@c��\$DIܔ
"23UDF�  ǀ~ LW�(VELqIN�b)@� _BL�@u��$G�q��$�'�'�%`<�� E�CHZR/�TSA_,`� ���E}`<�!���5�Bu�1}`_�� �)5D2d&�L@5I��N9t&��D�H�A���ÀP$aV `�#>A$�X�Ͳ�$Q�p�R}ӆ��H ��$BELvᵆ<!_ACCE�!c��7/���0IRC_] ��pNTT��S$P	S�rL� d�/Es ��F{�@F
��9gGDCgG36B���_�Q��2�@�A���1_M�GăDD�A]"ͲFW�`���3�EC�2�H�DE�KPPABN<>G��SPEE�B�Q %_pB�QY�Y��11�$USE_��,`P.k�CTReTYP�0Z�q P�YN��Ae�V)хQM���ѷ��@O� YA�TINC o�ڱ�B�DՒ�WG֑ENC����u�.A�2�Ӕ+@INPOQ�I06Be��$NT�#�%NT23_�"�2IcCLO� �2_`��I� _�if� _�k�? �` e�j�C400fMOSI��A���ОA䃔�PERCH  �c��B" �g��c��lb=���@��oUu@�@	A6B(uLeT	~�1eT�8ljgv�fTRK@%�AY��"sY��q6B�u��s۰�]��RU�MO1Mq�ՒY�MP�^���C�s�CJR��D�UF �BS_BCKLSH_C6B)��� �f���St�H��RR��Q>DCLALM-d��8�pm0��CHK��>�GLRTY����d��Y��)Üd_U	M]�ԉC��A!�n=PLMT� _L�0��9��E�.� � �#E)�#H� =��Q3pLo�xPC�axHW�8頿EׅCMCE��@.�GCN_,ND�Ζ&�SF�1�iVoR���g<!��6B���CATގSH)�,�Df Y��f��7A���܀3PAބ�R_P݅�s_ �v���s����JG�T]���Y�|����TORQUaP0��c�yPOU��b��P%�_W�u�t�@�1D��3C��3C�IK�IY�I�3F�6��X���@VC�00RQ�t��1���@ӿ��ȳ�JRK�����UpDeB M��UpMC� sDL�1BrGRVJ�`Cĭ3Cĳ3$�H_��8"�j@q�COS~˱~�LN���µ�ĭ0 �����u����̓��1Z���f$�MY��������>�THET=0reNK23�3h�l�3��CBm�CB�3C! AS� ��u����3��m�SB�3��x�'GTS$=QC������������$DU��Kw�B�%(��%Qq_��a��x�{�AK���b(��\�A`�����p�{�{�LPH~�g�Aeg�Sµ���� ����g������֚�EV��V��0��V��UV��V��V��V	�V�V%�H������P��G�����H��H��UH	�H�H%�O��O��OV	��O��O���O��O��O	�O
�O�Fg���	������SPBALA�NCE_-�LE6��H_`�SP!1���A��A��PFUL�CElTl��.:1=��UTO_�����T1T2��22N ���29`�\1�qnL�(=B�3�qTXpOv 
A>4�INSEG�2�a�REV��`aDI�F�uS91�8't"1�tpOB.!t�M��w�2�9`��,�LCHgWARRCBAB�� ��#�`-ФQ 5�X�qPR��&��2��� 
�""��1eROB͠CR6B5��_ 
�C�1_���T � x ?$WEIGH�P`#$��?3àI�Qg`sIFYQ�@LAG�R�q�S�R �RBIL�x5OD�p�`V2ST�0V2P!t�W0�11�&1/0�30
�P�2�Q�A  2řd[6D�EBUg3L_@�2��MMY9&E N8z�D`$D_A�a�$�0��O� �!0DO_@A.1� <B0�6�m�Q�IB�2�0N-cdH_p`�P �2O�� �/� %��T`"a���T/!�4)@TICYKh3| T11@%�C� ��@N͠�XC͠R�?��Q�"�E�"�E8@P�ROMP�SE~� $IR��Q��8R;pZRMAI)��Q4�R4U_r02S; t�q�PR8�COD�3sFU�Pd6ID_[��vU R!G_SU;FFu� l3�Q;Q�BDO�G �E�0�FGRr3�"�T�C �T�"�U�"�Uׁ�T8D��0�B0Hb _FIv�19*cORD�13 50�236V�+b|�Q1@$ZDT}U�s0�1;E�4 *:!L_NAmA�@�b>�EDEF_I�h�b �F�d�E�2�F�4�F�c�E�e�FISP��PAKp�Ds�C�d��44בi��2D�"�It��3D�O#OBLOCKEz��S�O�O�Gq�R�PUM�U�b�T �c�T�e�T!r�R�s�U �c�T�d�R�6�q�S � ���U�b�U�c�S�Z��X�@P` t�@q�e�)@W�x���s����TE�<D��( l1LOM�B_��ɇ0V2VI]S;�ITYV2A��}O�3A_FRI���a SIq�QR��@��@�3�3V2WB��W�4����_e��QEAS^3�Rϡ��P_�[p:R�4�5��6_3ORMULA�_Iz���THR.^2�Gtg�30f���<8�5COEFF�_O�A	 ��A��GdR�^3Sg0BCAn�O/C$��]3���0G�RP� � � �$�p�YBX�@TM~w���u�B�s��bC�ER, Tttsd�0ɛ  �LL�TSpS~�_SVNt�ߐ����0����0� ވ�SETUsMEA*P�P��W0�1+b/0�� � h��  @ڐo�l�o�cqz�"�b�@cqq`tP�AG��R�� Q\p*q�[p��>�c NPRE�C>at�5@MSKy_$|�� PB1?1_USER�e"��{ ���VEL@���{ 0�$Ō!I]`���MT�ACFG>���  �@@ =O�"NORE-0l@,o�V�SI.1�d��6��"UXK�fP!��D�E�� $KE�Y_�3�$J3OG��0SV���0���!��}�SW�"�ah\aS�ՐT|�GI����| ^�� 4 �h��'d2�!XYZ�c���3� ��_7ERR#�� 8Ԡ�AfPV�d��1����_$BUF��X��ܴ��MOR|�� HB0CUd�lA�!���GQ\aB�,"!a	$� ���a�����?�G~�� � �$SIՐ���VOx��T�0OBJE_���ADJU)B��EGLAY���%�DR�OU.`=ղВQ0b=��T���0���;BDIR���; I�"0DYNW�#���	T��"R���@�0�"�OPWORK����,%@SYSB9Uy�SOP��$ޑ�U�; P�pN�<�PA�t�>�"��+OP�PUd!0�`!z��l�IMAGw�1B0y�2IM�Õ��INe�d��RGO�VRD��-��o�P q��0��J�Os���"�L�pBa���o�PMGC_Ee`���1Ny M A�21�2U����SL_��� � ?$OVSL�ǫň?q�`��2�" -�_ ��k�P��k�Pu���2�C� �`�Ź����_ZER�D��$G�� 1�>���� @*���%MO~PRI��� 
�JP8+��=!/�L���ح�T� �0AT�US��TRC_T���sB��}fs��9s�1Re`��� DFAm����L���"��00a� ޱ��XEw{�����C0vcUP��+p	qPXPȝj�43 ���PG\���$S�UBe�%�qe9J?MPWAIT z�}%LO��F�A�R�CVFBQ�@x"�!R��� �x"ACC� R�&�B�'IGNR_{PL9DBTB�0Pqy!BWbP�$w��Uy@�%IGT�PI���TNLN�&2R���rL�NP��PE�ED \HADO!W�06�w��E[q4�jO!�`SPDV!� LbAz�`�07��3UNIr��0"!R��LYZ`� o���PH_PK��~e�RETRIE9�{�q����0'PFI�"�� �G`�0D �2�g�DBGL�V�#LOGSIZ,��EqKT�!U��VD�D�#$0_T�G�MBՐCݱ��|@eMRvC|}�3�CHECK0����PO�V!�k��I��LE(!��PA�rpT�2K�W��@P�2V!� h $ARIBiR� c�a/�qO�P8�ӐATT�� 2�IF|@z�Aq4S�3�UX���oaPLI�2V!� $g���I�TCHx"[�W �A�S9�2xRLLB�V!�� $B�A�DYs��BAM�!���Y9�PJ5Ƚ�Q��R6�V�Q_KGNOW�Cb��U��#AD�XV��0D�+i?PAYLOAt��BIc_��Rg�RgZOc�L�q��PLCL_�� !7��b�Q�B��d���fF�iC�֠�js��d�I�hR�ؠ�g�ҢdB����JL��q_J�a#���AND��Ĳ.t�b�a�L!q�PL0AL_ �P�0���Q�րC��DNcE���sJ3CpWv� TPPDCK������P��_ALPHgs�sBaE��gy|�K�|1�� � ����HoD_1Oj2ydDP�AR�*��;�&�^��TIA4U�5U�6��MOM��a����n���{�Y�B� AD�a���n���{�PUB��R��҅n�҅{����2�Wp��W �  �PMsbT� ����S���� e$PI��81��TgPJ��niJ�IV�Id�Ir��[��3!��>!���r�Ӫ�U3HIG�SU3�%�4얎4 �%� ���"����!
�<�!�%SAMP����^��_��%�P4s ю���[ 	ӝ�3  ���0���&�C�����^��Sp��H&0	�IN�SpB����뤕"���6��6�V�GAM�M�SyI�� ET�ْ��;�D�tA�
$NZpIBR!62IT�$HIِ_���C�˶E��ظAҾ���LWͽ�
���7����rЖ,0�qC�%CHyK��" �~I_A�����Rr�Rq�ܥ�Ǚ��ԥ���Ws ��$�x 1����I7RCH_5D�!� RN{��#�LE��ǒ!,��x����90MSWFL��$�SCR((100��R@��3]B��ç���a����َ0��PI�3A9�METHO�����%��AXH��XX0԰62ERI���^�3��R�0$u	D��pF{�_���?���1�L�L�_�a�OOP����wᲡ��'APP:���F���@0{���أRT�V�OBp�0T����;��� 1�I��� ��r����RA�@MGA1��B&�SV-��P�_@CURg�;�GRyO[0S_SA�QX��Y�#NO�pC! "�tY��Zolox��������!b����&�DO�1A���A����Х ��A���A"�WS��c P�QM)��o � ��YLH�qܧ��SrZ�]B��o�����ĵq_r�C1��M_W��B�g���c�M�  �`Vq�$p�x1�o�3"�PMJ�,�� !�'A� 9�!Wi:�$�LWQ|ai�t g�tg�tg{t� �AN`���S��SpX�0	O�sRqZ��P� *�W� ���M���� ����������X��� �N�@���P�q_~R� |�q#(Y����& n��&{�Y�Z��'�&t���Q�� &�"0����0}`�$PQ�P�MON_QUc� �� 8�@QCO�U��%PQTH��H�O�^0HYS:PES�R^0UEI0O��@]O|T�  �0PG�õz�RUN_TO��eOْ.�� �PE`�5C��A<�I�NDE�ROGR�AnP� 2g�NEg_NO�4�5IT���0�0INFO�1�C �Q�:A�Ȓ!�OIB� (��SLEQݖFAѕF@�6�POSy�T� =4�@ENAB��0�PTION.S%0E�RVE���G��wFG�CF�A� @R0JX$Rq�2���R�H��O�G "�EDI�T�1� �v�K��ޓʱE�NU�0W*XAUTu�-UCOPY�ِN\�����MѱNXP\[q�PR�UT9� _RN�@O;UC�$G�2�T>� �$$CL`� ���� ��a�&a� �P�S�@�Xw�PXK�Q�IRTU��_�PA�� _WRK 2 �e�@ 0  �5�QMoYh�Jo|m |l	 �`�m�oa�`��o�o�f�e�l}�a0I[ct'`BS�*�� 1�Y� <7���� ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������sr;CC��LMT� ����s  dѴI�Nڿ�дPRE_EXE��)�Ƅ0`jP��za'`DV���S�@e)�%�select_macro����kϤ�>qtIOCNVVB��k ��P��US�x�w���0V 14kP $$p��a�|�`?���߰>�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p ������� ���$�ѰLARMRECOV ^������LMDG ��Ь�LM?_IF ���d  YST-0�40 Opera�tion mod�e AUTO S���ed P) h�ang�(L:3)������)�;�M��_�q��, 
 ����#�>TEL�EOP ǘLIN�E 0ǑقABO�RTEDǘJOI�NT 100 %�����$���@��$�A��ATA�ǒؑ3��גؒ�� ? clear䀪����ί��NGTOL�  @� 	 �A |���ѰPPINFO �� f�L�^�p����  ������k��� ۿſ�����5��Y�0C�iϏ�%���ٯ�� ��������'�9�K��]�o߁ߓߙ�PPL�ICATION �?t���|�Hand�lingTool�ǖ 
V9.4�0P/17����
883ǀ����F90�	�549����|����7DF5�м��ǓNone���FRA�� �69��_ACTI�VE1�  �� � s ��ڀMOD���������CHGAoPONL�� �oOUPL[�1	��� >�B�T�f����CUREQ 1
���  Tp�p�p�	��������l��� ����������i3�l�p���^H��A�t
HTTHKY� FXv|�� *<N`���� ����//&/8/ J/\/�/�/�/�/�/�/ �/�/�/?"?4?F?X? �?|?�?�?�?�?�?�? �?OO0OBOTO�OxO �O�O�O�O�O�O�O_ _,_>_P_�_t_�_�_ �_�_�_�_�_oo(o :oLo�opo�o�o�o�o �o�o�o $6H �l~����� ��� �2�D���h� z�������ԏ��� 
��.�@���d�v���0��������TO������DO_CLEA�N���E�NM  �� p������ɯۯv�DSPDgRYRL���HI��o�@��G�Y�k�}��� ����ſ׿�������MAX��,�呿��=�X,�<�9�<���PLUGG,�-�9���PRC��Bm�"q�6�(ϗ�O���^�SEGF�K�� �� �m��G�Y�k�}�8������LAP$�7� �������+�=�O�a�s����� �T�OTAL_ƈ� �U�SENU$�1� �������RGDI_SPMMC�d��C�O�@@�1�O�"�D��-�_STRING 1��
�M��S���
��_ITE;M1��  n��� ������ $6H Zl~��������I/O SIGNAL���Tryout� Mode��I�npNSimul�ated��Ou�t`OVER�R!� = 100���In cyc�lT��Prog� Aborj��~JStatus���	Heartbe�at��MH F�aul��Aler�!/!/3/E/W/�i/{/�/�/�/  (���(����/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO�/WORИ�~A�/ XO�O�O�O�O�O __ $_6_H_Z_l_~_�_�_�_�_�_�_�^PO ���"`�KoEoWoio {o�o�o�o�o�o�o�o /ASew��bDEV%n�p9o ����#�5�G�Y� k�}�������ŏ׏������1�C�PALT�-j��OD����� ��ȟڟ����"�4� F�X�j�|�������į֯X�GRIB���� ���6�H�Z�l�~��� ����ƿؿ���� π2�D�V�h�z�����R �-��&���������� "�4�F�X�j�|ߎߠ� �������������PREGn�W���0� ~������������ � �2�D�V�h�z���������$�$AR�G_~@D ?	������  	$�$	[]��$:	��SBN_CONFIG�X�WqRCII�_SAVE  �$zm��TCEL�LSETUP �
%  OME�_IO$$%M�OV_H� ��R�EP��#��UTOoBACK� 	�tFRA:\�D� .D�z '�`�D�w� ��s  2�5/11/29 �20:26:16D�;D���#//h��C/j/|/�/�/�/�/D�X/�/?? (?:?L?�/p?�?�?�? �?�?�?g? OO$O6O HOZO�?~O�O�O�O�O��O�O���  c_�F_\ATBCK?CTL.TM�)_�;_M___q_8INI�m��j~CMESSAG� �Qz >�[ODE_D� ��j�XO�p�_@PwAUS6` !�� , 	��; :oHg,		 2oloVo�ozo�o�o�o �o�o�o 
D.P�z}d`TSK  �mw}_CUPD�T�P�Wd�p�VXWZD_ENB�Tf
�vSTA�U�u���XISX UNT� 2�vwy � �	 ����J �Ѽ �V�'��� G%��D�R��������M��l��K��_�m�����z�I���;�f)���x`t�:���s���p���4�MET���2@��y PQ�B�Ec�A�_yB�ߤBWl�B-��B�x���?;��>����?)"�?��W�?���@ K��5�SCRDCFG� 1Y; ��� ���%�7�I�pD�Q �	ܟ������ϯ�� Z��~�;�M�_�q���`����6���FGR9���p�_ԳPNA� �	FѶ_ED��P1��� 
 ��%-PEDT�-¿ R�v���E��<�GE�D�;�9/�>���  ����2�����B� ��ˀ�{�����j�����3 ��#� �G�Y���G����6�����4�W������Zݨ��Z�l������5K��ߘ�� Y�t���&�8���\���6��d��Y�@� ���(��7�S 0wY�w��f����8����{�I Z��C/��2/���!9{/��//LZݤ/�?V/h/�/�/��CR ���?�?Tn?�? ?�2?�?V?԰!�NO_�DEL�ҲGE_�UNUSE޿дI�GALLOW 1��   (�*SYSTEM�*��	$SER�V_GR[�@`REG�E$�C���@�NUM�J�C�MP�MU?@��LA�YK���PM�PAL�PUCYC10 N3^P!^YSULSU_�M5Ra�CLo_�TBOX�ORI�ECUR_��P�MPMCNV6V�P10I^�PT4DLI�p�_�I�	*PROGRA��DPG_MI!^Ko]`AL+ejoTe�]`B�o�N$F�LUI_RESU`9W�o�O�o�dMR�N�@�<�?�;M_ q������� ��%�7�I�[�m�� ������Ǐُ�����!�3�E�W�2BLAL_OUT �K����WD_ABO�R:PcO��ITR_�RTN  �$��빸�NONSTO��� lHCCF�S_UTIL ��̷CC_AU�XAXIS 3$� h}�j�|������ƽCE_RIA3_I`@�נ���FCFG �$�/�#��_L�IM�B2+� ��� � 	��B\T���$� 
Ԡ��)+�Z���/�����[�����.R���!�����L��(
5������PA�`GP 1H�����A�SϨe�w�6�CC� CU7��J��]��p��}����� C���U������������Ué�̩�ձ�ߩ�U�������;����PCk���������������������Ա��������� D� D!��!�!�!� ���&?��HE@O�NFIpC�G_�P�P1H�  +EH��ߟ߱�����������C�KPAUSf�Q1H�ף IR �S�H�A��e��� ������������E��+�i�{�a���A�?Iץ�MؐNFO� 1���� �3��$4�A��Y���[��2�#�@"��Nl,�*�����B����C�_��0C+��r�|�2��hPb�O� �� ��LLECT_��!�����EN�+`�ʒ���NDEַ#�/��1234567890�"�A��/ҵHw��#)j��< i{��;��/� �/`/+/=/O/�/s/ �/�/�/�/�/�/8?? ?'?�?K?]?o?�?�?@�?�?O�?��$�� ��IO #&��"S▒O��O�O�O`GTR�2'DM(��^�?�NN��(oM Z��_M[OR)q3)H��7� �U3��Y�_�_�_�_�_��[bR�kQ*H�CI?<�<Ѡ<cz�KFd����P,�� ;ϒo�o�o˿�o�oœh�UY@E�oS� �sja.�PDB.���4�cpmidbg03��Рs:��>uq�pz��v  E��>x��}.���}�`��|�<�m!gP���t��~f��������@ud1:��?��XqDEF �-��zC)*�c�O�buf.txt�J��|K�[`�/DM��>���R�A���MCiR20_{RCdX���hS21�����G���CzA�d4�E�I�jC%�eC�6� G/X"D�O[oF]�H��j�F� F��TWJ��iG�JI؂��LڒYJ4�JN�N��mKE�NMSo��d�����f23DL�D�	>z�!� 2���}��yc
�@�x9� C�Ĵ g D4G�E����  E%q�F�� E�p�u��F�P E���fF3H ��GM��Ъ5�>�33��?�x�n9�q@�Q5�����RpA?a��=L_��<#�QU�@�,�Cϒ���RSMOFST +i������P_T1Ɠ4�DMA =ք�MO�DE 5dm�@���	Q�M;���%��?���<��M>��Ͷ�T�ESTc�2i�`�R��6�O�K�CN�A(B���n� 8��\��n�CdB���C�pp�����p:d�QS ��� P������4�I7>�)��>B8m5$��RT_c�PROG %j%��d�1�>h@NUSER��x��KEY_TBL � e�����	
��� !"�#$%&'()*�+,-./(:;�<=>?@ABC�c�GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����>���͓��������������������������������������������������?������4A8��LCK��F�y��S�TAT��2�X�_�ALM�����_A�UTO_DO��E�FDR 3:�i�2h&q[~��� BUOS�YST-322 �Auto sta�tus chec�k time o�ut ���i�$?TELEO8��i� ��)qA��ʜ@Ĭ������?�ڛ��MsB�õ��?*?��?�Mf=�o��TR��-����D.�B����C���B��N�*p�4�N4m�J5Hj5H��H>�i�BJ�d�BF�z�pZ��[~�bb�t����5/�M�*F�B�GA�+$���@�R��J�}B�Q�H����������2>���@�@����&�C�BxHCKH<B��6>Tbt���/��[��+ ���g?/$/�?�'�lS�!���rA��7�A��y��x��&߇BC��!@��?�1�?�*���0��0&����@ڒ�����Ba��5�&�-�tO�tD�:O���/�/?�u�AUS�O�O�Oi�$�O _:�c@m� _J_p�� N_8_�_�_V_�_�_�_ �]�Oo)o;o�OLoqo _�o�o�_�o�o�o�o �o�oFXo� �No���o�� ��@�N�$�b�x��� ��n������A� �b�\�z�|�n����� ��ʟ���(�֏O�a� s������T�ʯį� �֯����2�H�~� ��>���ɿۿ���� ��2�,�J�L�>�xφ� \Ϛϰ����Ϧ��1� C��T�y�$Ϛߔ߲� �ߦ���������N� `�߇���V߼��� ��������H�V� ,�j�������v��� ��$I��jd�� �v����� 0��Wi{&�� \�����/&/ �:/P/�/�/F�/�/ �/��/?�:?4?R/ T?F?�?�?d?�?�?�?  O�/'O9OKO�/\O�O ,?�O�O�?�O�O�O�O �O
_ _V_h_O�_�_ �_^O�_�_�O
oo"_ $ooPo^o4oro�o�o �o~_�o	�_,Q �_rl�o�~�� ���&�8��o_�q� ��.����dڏԏ� �� �.��B�X��� ��N�ǟٟ럖���!� ̏B�<�Z�\�N����� l����������/�A� S���d���4�����¯ Ŀ�����Կ�(�^� p���ϩϻ�f����� ����*�,��X�f� <�zߐ����߆���� #���4�Y��z�t�� ������������.� @���g�y���6���� l�����������(6 J`��V��� ���)��JDb dV��t��� /�7/I/[/l/�/ <�/�/��/�/�/? �/?0?f?x?&/�?�? �?n/�?�?�/OO2? 4O&O`OnODO�O�O�O �O�?__+_�?<_a_ O�_|_�O�_�_�_�_ �_�_ o6oHo�Ooo�o �o>_�o�ot_�o�oo �o0>Rh� �^o����o�1� �oR�L�jl�^����� |���Џ���?�Q� c��t���D�����ҏ ԟƟ ���"�8�n� ��.�����˯v�ܯ� ��"��:�<�.�h�v� L�����ֿ迖��!� 3�ޯD�i���τϢ� �ϖ����ϴ����>� P���w߉ߛ�FϬ��� |�����
����8�F� �Z�p���f����� ����9���Z�T�r� t�f�����������  ��GYk�|� L������� �*@v�6�� �~�	/�*/$/B D/6/p/~/T/�/�/�/ �/�?)?;?�L?q? /�?�?�/�?�?�?�? �?�?OFOXO?O�O �ON?�O�O�?�O�OO __@_N_$_b_x_�_ �_nO�_�_o�OoAo �Obo\oz_|ono�o�o �o�o�o(�_Oa so��To���o �����2�H�~� ��>��ɏۏ��� �2�,�J�L�>�x��� \�����������1� C��T�y�$������� ������į��N� `��������V���� ��������H�V� ,�jπ϶���v���� ߾�$�I���j�d߂� ��v߰߾ߔ������ 0���W�i�{�&ߌ�� \������������&� ��:�P�����F���� ��������:4R� TF��d���  ��'9K��\� ,������� �
/ /V/h/�/�/ �/^�/�/�
??"/ $??P?^?4?r?�?�? �?~/�?	OO�/,OQO �/rOlO�?�O~O�O�O �O�O�O&_8_�?__q_ �_.O�_�_dO�_�_�O �_�_ o.ooBoXo�o�tc�$CR_FD�R_CFG ;�re�Q
�UD1:�W�P:�PJ�d  �`�\��bHIST 3<�rf  �`  w?�R@tuAtB�bC�PUYpDtEtItUg�Ppotw�_���bINDT_E�N6p�T��q�bT1_D�O  �U�u�sT�2��wVAR 2m=�gp hq�  -�t���t�R��4�����m[��RZ�`ST�OP��rTRL_�DELETNp�t ���_SCREE�N re�r�kcsc�rUw�MMENU 1>���  <�\% �_��T��R��S/� U���e�w�ğ������ џ�	�B��+�x�O� a�����������ͯ߯ ,���b�9�K�q��� ����࿷�ɿ���� %�^�5�Gϔ�k�}��� �ϳ��������H�� 1�~�U�gߍ��ߝ߯� ������2�	��A�z� Q�c��������� ��.���d�;�M��� q������������Y�Ӄ_MANUAL�{��rZCD�a?x�y�rG ���R��f"
�"
?|�(��PdTGRP� 2@�y�B1� � s��� ��$DBCO�pR�IG���v�G_E�RRLOG A���Q�I[m ��NUMLIM��s��u
�PXWORK 1B�8���//�}�DBTB_�� !C%���S"� ��aDB_AWAYz��QGCP �r�=�ןm"_AL(�F�_�Yz���p�p�vk  1D� , 
��/"�/%?/(_M�pqw,�@�=5ONTIM6����t�_6�)�
�0�'MOTN�ENFpF�;REC�ORD 2J�� �-?�SG�O� �1�?"x"!O3OEOWO �8_O�O�?�OO�O�O �O�O�O(_�OL_�Op_ �_�_�_A_�_9_�_]_ o$o6oHo�_lo�_�o �_�o�o�o�oYo}o 2�oVhz��o� �C�
��.�� R��K��������Џ ?��ߏ�*�����+� b�t�㏘�����Ο=� O�����:�%���p� ߟ񟦯��O�ǯ�]� �����H�Z����� ����#�5����ϩ��i"TOLEREN�Cv$Bȿ"� L���� CSS_CC�SCB 2K�\0"?"{ϰϟ� ��7��
����@�R� d�3߈ߚ�"�x��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy���� �������R�LL]�La��m1T#2 C��C��F�^ +A�C�pC���#�0�� 	 A����B���?�  �$�����\0袰�0��B� �`#s�K/]/o/�ϓ/�/�/s/�/�/��K{�0Le��>5�1�r��9Kr�Ȧ�/��/`?;
�@��O?�?�?�?�Ȏ0AF��?{F�A OO�7�1���9M	AB
AZOdBAE�9�$O�O�O�Oi:P��`^�@0�DJCA�� @��
qX-.
[#_   M?�>O�ڴ�q_�_�_�_:W�A<o:[@<ǲ/o�/�_+o`Poboto�eACHC�jV�WB$�Dz�cD�`�a=/�o�oo�oHW�a.+!��2=t ,y�J?�.s�s�js �w�yj�������Q�Qs�@`�� $�����A����Bމ �o��'�9��_]�o� N���r���ɟ۟_�B��ʄ��YZ>`�>���A��zB��@��6>V?�y��X0�Z�l�~����`_м ¯���
���̯9�,� ]�o��� �H�����ٿ 뿊��ƿ3�E�W�i� ����$ϱ����� Ϟ� ���/�A�S߶�w�V߀h߭ߌ��S���ߐ�_�f	��H�?�Q� ~�u��������� ���D��-�g�q� ������������
 @7Icm�����  ���� �)M@qdv �������/ /I/P�m/�v/�/�/ �/�/�/�/�/?3?*? <?i?`?r?�?^/�?�? �?�?�?O/O&O8OJO \O�O�O�O�O�O�O�O��g	  QU�P�s �PWC4p*p�p�6U6P\C9p/�p�� ]V^PM]Ê6P�:P�>P�VJ_�^P�bP�fP�Vr]&v���p Q
k���_oo�id1Q&oNo ;o_co�oˏUU�A   �o�k1Q@��  �o�k�b�.�����p �� 1��6�01C����C�cPfL��?#~�c>�{���`�cP�@@�d��r��`B�cP>�s�qC���p����b�t<��o?�PH�)S�B�tq�q�p�r�`B���eI"C�&�Q�4( �oz��UU�:��9��@����>V�^��/Q�-R@`����W�c���Bg�)�b�<�`ځ`  ?�p�x��U�[?���}t���$���$DCS�S_CLLB2 {2M��p��P�^?�NSTCY� 2N���  ����� ��ʟ؟���� �2� D�Z�h�z�������¯�ԯ��SA�DEVI_CE 2O��!�$��4&V�h����� ��˿¿Կ���
�7� .�[�R�ϑϣϵ������4(A�HNDGDg P��*�Cz�A�LS 2Q�� _�Q�c�u߇ߙ߽߫����?�PARAM �RP��1�`�&�R�BT 2T�� �8�P<C�'p# �qi�l��s@"��R��(qI�X��y0�pB CW  ��B\x�N��`Z����%��)���X�j� �p����zq�����B 	�(s,�F�p�V���q���b��B ��4&c �S�e�l�4+�����H1~���{�D�C�$Z���b���A,� 4��u@�X@���^@w���]Bߣ��B�cP%���C4�C3:_^C4��nЬ ���p8�-B�{B��A������ l��C��C3�JC4�jC3��yn+��3 Dff 2��A PB W4+@ :�]o�W��� ��/�/P/'/9/ K/]/o/�/�/�/�/? �/�/�/?#?5?�?Y? k?�?�?�o�?�?O�? 6O!OZOlOWO�O�Es �?�?�?�O�O_�O�O L_#_5_G_Y_k_}_�_ �_�_ o�_�_�_oo 1o~oUogo�o�o�o�o �owO D/Az e����O�o�o
� �o��R�)�;���_� q����������ݏ� <��%�r�I�[�m��� �����ǟٟ&�8�� \�G���k�������گ ů�����F��/� A�S�e�w�Ŀ������ ѿ�����+�x�O� aϮυϗϩϻ����� ,���b�t�ﯘ߃� �ߧ���������:� �C�U߂�Y�k��� ���������6��� l�C�U�g�y������� ���� ��	-? Q������� @+dvQ� �������*/ //%/r/I/[/�// �/�/�/�/�/&?�/? \?3?E?�?i?{?�?�? U�?�?"O4OOXOCO |OgO�O{��?�O�? �O�O0___f_=_O_ a_s_�_�_�_�_�_o �_oo'o9oKo�ooo �o�o�o�o�o�O: %^I�������H�$DCSS�_SLAVE �U���	����z_4D � 	��AR_M�ENU V	�  �j�|�������ď�B�Y�� ��~?�SH�OW 2W	� � �b�aG�Q�X� v���������П֏���� @�:�d�a�s� ���������߯�� *�$�N�K�]�o����� ��̯ɿۿ���8� 5�G�Y�k�}Ϗ϶��� ��������"��1�C� U�g�yߠϝ߯����� ���	��-�?�Q�c� ��s����������� ��)�;�M�t���� ������������ %7Ip�m���� ������!3 ZWi���J� ���//DA/S/ e/��/��/�/�/�/ �/?./+?=?O?v/p? �/�?�?�?�?�?�?? O'O9O`?ZO�?�O�O �O�O�O�OO�O_#_ JOD_nOk_}_�_�_�_ �_�O�_�_o4_.oX_ Uogoyo�o�o�o�_�o �o�ooBo?Qc u���o:����CFG X)��3�3q5p�_FRA:\!�L+��%04d.CSVj|	p}� �q[A g�CHo�zv��	����3q������́܏� ���4���JP����q�p1� �RC_O�UT Y���C��_C_F�SI ?i� .������� ͟�����>�9�K� ]���������ίɯۯ ���#�5�^�Y�k� }�������ſ���� �6�1�C�U�~�yϋ� �����������	�� -�V�Q�c�uߞߙ߫� ���������.�)�;� M�v�q������� �����%�N�I�[� m��������������� ��&!3Eni{ ������� FASe��� �����//+/ =/f/a/s/�/�/�/�/ �/�/�/??>?9?K? ]?�?�?�?�?�?�?�? �?OO#O5O^OYOkO }O�O�O�O�O�O�O�O _6_1_C_U_~_y_�_ �_�_�_�_�_o	oo -oVoQocouo�o�o�o �o�o�o�o.); Mvq����� ����%�N�I�[� m���������ޏُ� ��&�!�3�E�n�i�{� ������ß՟����� �F�A�S�e������� ��֯ѯ�����+� =�f�a�s��������� Ϳ�����>�9�K� ]φρϓϥ������� ����#�5�^�Y�k� }ߦߡ߳��������� �6�1�C�U�~�y�� �����������	�� -�V�Q�c�u������� ��������.); Mvq����� �%NI[ m������� �&/!/3/E/n/i/{/ �/�/�/�/�/�/�/3��$DCS_C_�FSO ?����71 P ??T?}? x?�?�?�?�?�?�?O OO,OUOPObOtO�O �O�O�O�O�O�O_-_ (_:_L_u_p_�_�_�_ �_�_�_o oo$oMo HoZolo�o�o�o�o�o �o�o�o% 2Dm hz������ �
��E�@�R�d��� ������ՏЏ��� �*�<�e�`�r����� ����̟�����=��8�J�\�������?C/_RPI4>F?�� �����3?�&�o�X���� >SLү@d� �����%�7�`�[� m�Ϩϣϵ������� ���8�3�E�W߀�{� �ߟ����������� �/�X�S�e�w��� ����������0�+� =�O�x�s��������� ����'PK ]o������ ��(#5Gpk }�����Q��� /6/1/C/U/~/y/�/ �/�/�/�/�/?	?? -?V?Q?c?u?�?�?�? �?�?�?�?O.O)O;O MOvOqO�O�O�O�O�O �O___%_N_I_[_ m_�_�_�_�_�_�_�_ �_&o!o3oEonoio{o �o�o�o�o�o�o�o FASe������>�NOCO�DE ZU���?�PRE_?CHK \U��p�A �p�< ��pU�]�o�U� 	 <Q������ ��ۏ�Ǐ�#���� Y�k�E�����{�şן ��ß����C�U�/� y�����s���ӯm��� 	���?��+�u��� a�������ɿ�Ϳ߿ )�;��_�q�K�}ϧ� �������ω���%��� �[�m�Gߑߣ�}߯� �߳����!���E�W� 1�c��g�y������ �������A�S�-�w� ��c����������� ��+=asM_ ������' �]o	�� ����/#/�G/ Y/3/e/�/i/{/�/�/ �/�/?�/?C?9K y?�?%?�?�?�?�?�? 	O�?-O?OOKOuOOO aO�O�O�O�O�O�O�O )_____q_K_�_�_ a?�_�_�_�_o%o�_ Io[o5oGo�o�o}o�o �o�o�o�o�oEW 1{�g���_� ���/�A��M�w� Q�c����������Ϗ �+���a�s�M��� ������ߟ���'� ��3�]�7�I������ ɯۯ�������G� Y�3�}���i���ſ�� ������1�C���+� yϋ�eϯ��ϛ����� ����-�?��c�u�O� �߫߅ߗ�������� )��M�_�U�G��� A������������� I�[�5����k����� ��������3E Q{q���]� ���/Aew Q������� /+//7/a/;/M/�/ �/�/�/�/��/?'? ?K?]?7?�?�?m?? �?�?�?�?O�?5OGO !O3O}O�OiO�O�O�O �O�O�/�O1_C_�Og_ y_S_�_�_�_�_�_�_ �_o-oo9oco=oOo �o�o�o�o�o�o�o __M_�ok�o �������� I�#�5����k���Ǐ ��ӏ��׏�3�E�� i�{�5c���ß��� ��ӟ�/�	��e�w� Q�������ѯ㯽�ϯ �+��O�a�;����� ���Ϳ߿y���� !�K�%�7ρϓ�mϷ� �ϣ���������5�G� !�k�}�W߉߳ߩ��� ���ߕ��1���g� y�S�������� ���-��Q�c�=�o� ��s��������� ����M_9��o �����7 I#mYk�� ����!/3/)/ i/{//�/�/�/�/�/ �/�/?/?	?S?e??? q?�?u?�?�?�?�?O O�?%OOOE/W/�O�O 1O�O�O�O�O__�O 9_K_%_W_�_[_m_�_ �_�_�_�_�_o5oo !oko}oWo�o�omO�o �o�o�o1Ug AS������ 	����Q�c�=��� ��s���Ϗ�o���� ��;�M�'�Y���]�o� ��˟����۟�7� �#�m��Y������� �����!�3�ͯ?� i�C�U�������տ� ������	�S�e�?� �ϛ�uϧ��ϫϽ�������$DCS_SGN ]	��E��-����01-DEC-�25 19:20� ��29-N�OVV�20:27�_�x�x� [}�t��q�т�x���ك�JѨ�EƼÞ� ��ǖ��  1�HOW �^	� �x�/�VERSI�ON =��V4.5.2��E�FLOGIC 1�_���  	������C��R�%�P�ROG_ENB � ��:�{�s�U?LSE  X���%�_ACCLI�M�����d���WRSTJNT��E��-�EMO�|�zя�$���INIOT `2�����OPT_SL ?�		�	�
 	�R575��]�74jb�6c�7c�50���1���C���@�TO  L��� �]V�DEX��dE��x�PATH ;A=�A\k�}��HCP_CL?NTID ?�:� D�ռ���IAG_GRP �2e	�����z�	 @� � 
ff?aG���B�  �2��/�8[I@�c�ς!�7@��z�@^�@�
�!��mp�2m15 8901234567�����  ?���?�=q?���
?޸R?��Q�?��?������(�?Ǵz���x�@�7  A_�Ap !�7A�88_�B4�� ��L�x��
�@�@���\@~�R@x�Q�@q�@j��H@c�
@\���@U�@Mp��//'$�; |�O)H��@Ct }>d 9��@4�_/\)@)� #t {@��/��/�/�/�/P'?�̗�?���_ ?�}p�?u?on{?s ?\�Q�? ?2?D?V?�h8�
=?����0w5�z�H?�p�h��?^�R�?�?�?�?�?h8�U�t0���@�?��0�;@&O 8OJO\OnOP'�$_� _Y_k_�O?_�_�_�_ �_�_s_�_�_1oCo!o goyoo�o��Bj"� ��2{1�@"?����f�t0�d"5!=�
u4V��u"��B3t�A>u��?@�[q��@`,=q��=b��=�E�1>�J�>�n��>��H"<�;o �z�s�q���� �x�C�@<(��Uz� 4��� ����A@x�? *�o��m*�P�b�� �tn���2���Ώ�����i>J��&��bN2�"��G��N��o@�@v���0����@ffr!�l ��33���({��"C�� ƒ�I�CH�)C.dBت"8"����'���"~��A?�&"K����pf�B��@�p�������p���?5���3|�Y=�y�2��/�6�B��6�5=���6
*��~�`C���B���C�_�xВ������3���N�T������0C+�r�|�2�G#�����ȿ�� �׿����?,�<��o��CT_CON�FIG f�|�|�egY���STBF_TTS��
����О�}�:��1�MAU����~��MSW_CF���g�  # ��OCoVIEW��h!�-���s߅ߗߩ� ���ߟ�a�����,� >�P���t����� ��]�����(�:�L� ^�������������� k� $6HZ�� ~������y  2DVh��������v�RC�i���!���/ S/B/w/f/�/�/�/���SBL_FAUL�T j*6��!G�PMSK���'��TDIAG k���-�������UD1: 6789012345I2��=1�Ǥ�P\υ?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�Od6�96���r
t?�O|�TORECP"?4:
B4 4_[7��s?p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�O�O�O��o7�UMP_OP�TIO=��.�aT�R����)uPM�E��Y_TEM�P  È�3�BC�gp�B�QtU�NI����gq�YN_BRK lL�~7�EDITOR�a��a@�r_
PENT� 1m)  �,&TELEO�[p���&SET_WCp,��l�pPSNAP^PX�?�MTPG�pW�i� �/��IĦ��ʏ�� �=�$�a�H�����~� ����ߟ�؟���9�  �2�o�V���z���ɯ ���ԯ�#�
�G�D���pMGDI_ST�AzuV�gq�uNC_INFO 1n!��b���X�����غ���n�1o!� ���o����
�d �oU�g�yϋϝϯ��� ������	��-�?�Q� c�u߇ߙ߽߫��� u ����
��*�B�*�P� b�t��������� ����(�:�L�^�p� ��������2������� 9�CUgy� ������	 -?Qcu��� �����//1;/ M/_/q/�/�/�/�/�/ �/�/??%?7?I?[? m??�?�?�?��?�? �?O)/OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�_ �_�?�?�_�_o�_3O =oOoaoso�o�o�o�o �o�o�o'9K ]o����_�_� ���+o5�G�Y�k� }�������ŏ׏��� ��1�C�U�g�y��� �����ӟ���	�#� -�?�Q�c�u������� ��ϯ����)�;� M�_�q���������˿ ݿ����7�I�[� m�ϑϣϵ������� ���!�3�E�W�i�{� �ߟ߹���������� %�/�A�S�e�w��� �����������+� =�O�a�s��������� �������'9K ]o������ ��#5GYk }�	������ /1/C/U/g/y/�/ �/�/�/�/�/�/	?? -???Q?c?u?�?�?� �?�?�?�?/O)O;O MO_OqO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�?�_�_�_�_ O�_!o3oEoWoio{o �o�o�o�o�o�o�o /ASew��_ �_����o�+� =�O�a�s��������� ͏ߏ���'�9�K� ]�o�������ɟ۟ ���#�5�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�q߃ߝ��߹��� �������%�7�I�[� m����������� ���!�3�E�W�i�{� �߇���������� /ASew�� �����+ =Oas������ ����//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? ���?�?�?�?��? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�?�_�_ �_�_�?�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ m�_u����_� ��!�3�E�W�i�{� ������ÏՏ���� �/�A�S�e���� ����u������+� =�O�a�s��������� ͯ߯���'�9�K� ]�w���������ɿ� ����#�5�G�Y�k� }Ϗϡϳ��������� ��1�C�U�g߁��� �߯���ۿ����	�� -�?�Q�c�u���� ����������)�;� M�_�y߃��������� ����%7I[ m������ �!3EWq�c ���������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?i{�?�?�?�? ��?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_�?s? }_�_�_�_�?�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qk_u��� �_�����)�;� M�_�q���������ˏ ݏ���%�7�I�c Q���������ٟ� ���!�3�E�W�i�{� ������ïկ������/�A�[� �$E�NETMODE �1p����  k�k��f�����j�OATC�FG q�����Ѵ��C����DATA 1r�w�Ӱ���*	�*��'�9�K�]�l�dlύ�e��ϻ� ��������'ߡϳ� ]�o߁ߓߥ߷�1��� U����#�5�G�Y��� �ߏ����������� u��1�C�U�g�y��� ���)�������	 -����cu������j�RPOST�_LO��t�[
�׶#5Gi�RR�OR_PR� %�w�%L�XTAB_LE  w�ȟ�����RSEV�_NUM ��  ���  ��_AUTO_EN�B  ���X_;NO5! uw���}"  *�x ��x �x �x + +�w �/�/�/Q$FLT9R=/O&HIS#]��J+_ALM 1]vw� �[x,e�+�/Q?c?u?�?ș?�?�/_"W   �w�v!���:j�T�CP_VER �!w�!x�?$EX�T� _REQ�&9�H)BCSIZKO=D�STKhIf%�~?BTOL  ]{Dz�"�A =D_BWD�0�@�&�A쟲�CDI�A w�ķ���]�KSTE�P�O�Oj�POP_�DO�Oh�FDR_?GRP 1xw��!�d 	�?�_��yP�s�Y�Q'�M�"���l���T� ����VyS�_�]�TA8���AU��@�d��_�_ okGo2oWo�}oho�o�o�om?����@p�?���=����n
? L��z$b�` �o���3:�o^I��hA@`�t@S3	3�uh}@�q�g�<�yPF@ ��|�yPG�  @�Fg?�fC�8RL��}�?��`i��~6�X�����875t���5���5`+���~��� ������� Z�k�� �����FEATUROE y���@���Handl�ingTool ��]Engl�ish Dict�ionary�4�D St��ard���Analog� I/O>�G�gle ShiftZ��uto Soft�ware Upd�ate�mati�c Backup����ground� Edit ��C_ameraU�FY��CnrRndIm����ommon �calib UI���nˑ�Monoitor$�tr�?Reliabn���DHCP �[�at�a Acquis�3�\�iagnos���R�v�ispla�yΑLicens�Z�`�ocument Viewe?��^�ual Che�ck Safet�y��hance�d���s�Fr�ܐ�xt. DI�O /�fi��@�e�nd�Err>�L(��\�4�s[�rP�K�� �@
�FCTN /Menu��vZ����TP In��faycĵ�GigE־��Đp Mask� Exc�g=�H�T԰Proxy �Sv��igh-wSpe�Ski��� Ť�O�mmuni�c��onsV�ur໰��q�V�ײcon�nect 2��n{crְstru!�$�ʴ�eۡ��J��X��KAREL Cmod. L�ua�~��Run-Ti<��Env�Ȟ�el u+��s��S/W��ƥ���r�Book�(System)�
�MACROs,~M�/Offseu��p�HO���o�u�MR�8�4���MechStop+�t����p�im�q���x�R������odo�witc�h�ӟ�.��4�O�ptmF��,�fi�l䬳�g��p�ul�ti-T�Γ�P?CM fun�Ǽ��o��������Regeie�rq���riݠ�F���S�Num �Sel��/�:� Adjua�*�W�q�h�tatu��ߪ��RDM Robo}t�scove'���ea��<�Fre�q Anlyq�Rem��O�n5�����ServoO�!��?SNPX b-�v�;SN԰Cliܡ?r�Libr&�_��Q ��q +oJ�t���ssag��X�@ 0����	�@/Iս��MILIB��P� Firm���Pλ�AccŐ͛TPsTXk��eln���������orq}uo�imula=�4�|u(�Pa&���ĐX�B�&+�ev.̸��ri��TU�SB port ��iPf�aݠ&R� EVNT� n?except�����%5��VC�rl�c���V���"�%4q�+SR SCN�/gSGE�/�%UI	�?Web Pl��>���A43��ۡ��ZDT Applj�<
�{1EOAT�����&0?�7Gridp�񾡬=�?iR�"�.5� F���/גRX-10iA/L�?�Alarm Caouse/��ed(��All Smoo�th5���C�sciyi+�V�Load�ΌJUpl�@w�to�S ��rityA_voidM(�s7�1t�@�ycn��0���_�CS+���g. c��XJo� ��-T3_H�.RX��U����Xcollabo����RA�:�.9�D��in���N�RTHI
�On��e Hel����ֿ������1trU�ROS Eth$��A� �����;,�G �B�,|HUpV�%�W�3t ԰�_iRS�ݐ��64MB DRsAM�o�cFRO8���L8F FlD���d��2M �A:�opm�bԕex@V�
�sh�qD��wce�u��p��|tyn�sA�
�%�Ar����J��^�.v� P)Q/sbS�`���8O�N��mai��U����R�q�T1��^FC+Ԍ%̋Fs�9�ˌk̋��Typ߽FC%�hױV�N Sp�ForްK��Ԇ��lu!����cp�P'G j�֡�RJ�[L`Sup"}���֐f��crFP��lu� ��al�����r��i�
q�4@�ް�uest,IMPLE ׀6*|H�Z���c0�BTeap(�|���$rtu���V�9HMI�¤��wUIFc�pono2D�BC�:�L�y�p� ��������ʿܿ	� � �?�6�H�u�l�~ϫ� �ϴ���������;� 2�D�q�h�zߧߞ߰� �������
�7�.�@� m�d�v������� �����3�*�<�i�`� r��������������� /&8e\n� �������+ "4aXj��� �����'//0/ ]/T/f/�/�/�/�/�/ �/�/�/#??,?Y?P? b?�?�?�?�?�?�?�? �?OO(OUOLO^O�O �O�O�O�O�O�O�O_ _$_Q_H_Z_�_~_�_ �_�_�_�_�_oo o MoDoVo�ozo�o�o�o �o�o�o
I@ Rv����� ����E�<�N�{� r�������Տ̏ޏ� ��A�8�J�w�n��� ����џȟڟ���� =�4�F�s�j�|����� ͯį֯����9�0� B�o�f�x�����ɿ�� ҿ�����5�,�>�k� b�tφϘ��ϼ����� ���1�(�:�g�^�p� �ߔ��߸������� � -�$�6�c�Z�l�~�� �����������)� � 2�_�V�h�z������� ��������%.[ Rdv����� ��!*WN` r������� //&/S/J/\/n/�/ �/�/�/�/�/�/?? "?O?F?X?j?|?�?�? �?�?�?�?OOOKO BOTOfOxO�O�O�O�O �O�O___G_>_P_ b_t_�_�_�_�_�_�_ oooCo:oLo^opo �o�o�o�o�o�o	  ?6HZl�� �������;� 2�D�V�h�������ˏ ԏ���
�7�.�@� R�d�������ǟ��П �����3�*�<�N�`� ������ï��̯��� �/�&�8�J�\����� ������ȿ�����+� "�4�F�Xυ�|ώϻ� ����������'��0� B�T߁�xߊ߷߮��� ������#��,�>�P� }�t��������� ����(�:�L�y�p� �������������� $6Hul~�����  ?H552���21R785�0J614AwTUP'545'�6VCAMC�RIbUIF'2�8cNRE52�VR63SCH�LIC�DOC�V�CSU86�9'02EIOC��4R69VEgSET?UJ7U�R68MASK^PRXY{7OCO#(3?+ �&3j&J6%53��H�(LCHR&O�PLG?0�&MH�CRS&S�'MCS�>0.'552MD�SW+7u'OPu'M�PRv&��(0&PCMzR0q7+ 2l� �'51J51�8�0JPRS"'69�j&FRDbFRE�QMCN93�&SNBA��'SHLBFM1G�8�2&HTC>TMsIL�TPA�oTPTXcFELF�� �8J9�5�TUTv'95�j&UEV"&UEC�R&UFRbVCC�
XO�&VIPnFC;SC�FCSG���IWEB>HTT>R6��H;RV�CGiWIGQWIP�GS�VRCnFDGvu'H7�7R66J�5'R�8R51*
(6�(2�(5V�)J8�86�L=I%� �84g662R�64NVD"&R�6�'R84�g79ڎ(4�S5i'J7�6j&D0�gF xR�TSFCR�gCR�Xv&CLIZ8IC�MS�Sp>STY:nG6)7CTO>���7�NNj&ORqS�&C &FCB��FCF�7CH>F�CR"&FCI�VF�C�'J�PO7GBfMv�8OLaxENDS&�LU�&CPR�7L�WS�xC�STxT�E�gS60FVmR�IN�7IHaF �я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� !3EWi{� ������ /ASew��� ����//+/=/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]? o?�?�?�?�?�?�?�? �?O#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �_�_�_�_�_	oo-o ?oQocouo�o�o�o�o �o�o�o);M _q������ ���%�7�I�[�m���������Ǐُ��  H55�2��21�R7�8�50�J61�4�ATUP7�5�457�6�VCA�M�CRI��UI�F7�28��NREv�52v�R63�wSCH�LICƚ�DOCV�CSU��8697�0F�E�IOCǛ4�R6=9v�ESETW�u��J7u�R68�M�ASK�PRXY���7�OCO��3�W����6�3�J6�5�536�H$�LC�HƪOPLGW�0^�MHCRǪS���MCSV�0��55�F�MDSW���OP��MPR���6��06�PCM��R0`E˓�F���6�51f��51��0f�PRSv��69�FRD���FREQ�MCN��936�SNBA�כ%�SHLB�M�E��ּ26�HTC�V�TMIL�6�T{PAV�TPTX��#ELړ�6�8%�#���J95��TUTv��95�UEV��wUECƪUFR���VCCf�O��VI�P��CSC��CS�Gƚ$�I�WEBnV�HTTV�R6՜���S���CG��IG���IPGS'�RC���DG��H7��RK66f�5�u�R��WR51f�6�2�I5v�#�J׼��6���LU�5�s�v�4��6�6F�R64�NV�D��R6��R84֦79�4��S5n�J76�D0u�FRTS&�CR�CRX��CLI&�e�CMSV�sV��STY��6�CT�OV�#�V�75�NN��ORS����6�F�CBV�FCF��C�HV�FCR��FC-IF�FC��J#�˵G
M��OL�E�NDǪLU��CPUR��Lu�S�C$��StTE�S60n�FVRV�IN��IH���m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s�@��������͏ߏ��STD�LANG���0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰����RBT
�OPTN������'�9�K� ]�o�����������DPN	���)� ;�M�_�q��������� ������%7I [m����� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	-?Qcu� �������� )�;�M�_�q������� ��ˏݏ���%�7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w� ��������ѿ���� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� ������1�C�U�g� y���������������@	-?Qc�f�������9�9��$FEAT�_ADD ?	����  	�#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������DEMO y?   �L� B�T߁�xߊ߷߮��� ��������G�>�P� }�t��������� ����C�:�L�y�p� �������������� ?6Hul~� �����; 2Dqhz��� ��� /
/7/./@/ m/d/v/�/�/�/�/�/ �/�/?3?*?<?i?`? r?�?�?�?�?�?�?�? O/O&O8OeO\OnO�O �O�O�O�O�O�O�O+_ "_4_a_X_j_�_�_�_ �_�_�_�_�_'oo0o ]oTofo�o�o�o�o�o �o�o�o#,YP b������� ���(�U�L�^��� ��������ʏ��� �$�Q�H�Z���~��� ����Ɵ����� � M�D�V���z������� ¯ܯ��
��I�@� R��v���������ؿ ����E�<�N�{� rτϱϨϺ������ ��A�8�J�w�n߀� �ߤ߶��������� =�4�F�s�j�|��� ����������9�0� B�o�f�x��������� ������5,>k bt������ �1(:g^p ������� / -/$/6/c/Z/l/�/�/ �/�/�/�/�/�/)? ? 2?_?V?h?�?�?�?�? �?�?�?�?%OO.O[O ROdO�O�O�O�O�O�O �O�O!__*_W_N_`_ �_�_�_�_�_�_�_�_ oo&oSoJo\o�o�o �o�o�o�o�o�o "OFX�|�� �������K� B�T���x�������ۏ ҏ����G�>�P� }�t�������ןΟ�� ���C�:�L�y�p� ������ӯʯܯ	� � �?�6�H�u�l�~��� ��Ͽƿؿ����;� 2�D�q�h�zϔϞ��� �������
�7�.�@� m�d�vߐߚ��߾��� �����3�*�<�i�`� r������������ �/�&�8�e�\�n��� ��������������+ "4aXj��� �����'0 ]Tf����� ���#//,/Y/P/ b/|/�/�/�/�/�/�/ �/??(?U?L?^?x? �?�?�?�?�?�?�?O O$OQOHOZOtO~O�O �O�O�O�O�O__ _ M_D_V_p_z_�_�_�_ �_�_�_o
ooIo@o Rolovo�o�o�o�o�o �oE<Nh r������� ��A�8�J�d�n��� ����яȏڏ���� =�4�F�`�j������� ͟ğ֟����9�0� B�\�f�������ɯ�� ү�����5�,�>�X� b�������ſ��ο�� ��1�(�:�T�^ϋ� �ϔ��ϸ������� � -�$�6�P�Z߇�~ߐ� �ߴ���������)� � 2�L�V��z���� ��������%��.�H� R��v����������� ����!*DN{ r������� &@Jwn� ������// "/</F/s/j/|/�/�/ �/�/�/�/???8? B?o?f?x?�?�?�?�? �?�?OOO4O>OkO bOtO�O�O�O�O�O�O�__0]   'XF_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o o&o8oJo\ono�o�o �o�o�o�o�o�o" 4FXj|��� ������0�B� T�f�x���������ҏ �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ����������
��.�  /�)�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?V?h?z?�?�? �?�?�?�?�?
OO.O @OROdOvO�O�O�O�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|� �������� 0�B�T�f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�\�n� ���������������� "4FXj|� ������ 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<N `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������P ��$�4�8�+� N�`�r߄ߖߨߺ��� ������&�8�J�\� n����������� ���"�4�F�X�j�|� �������������� 0BTfx�� �����, >Pbt���� ���//(/:/L/ ^/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?l? ~?�?�?�?�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�o&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�`�r����������� ����&8J\ n������� �"4FXj| �������/ /0/B/T/f/x/�/�/ �/�/�/�/�/??,? >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO ^OpO�O�O�O�O�O�O��O __$_6Y�$F�EAT_DEMO�IN  ;T��fP�<PNTIND�EX[[jQ�NPI�LECOMP �z����Q�iRIU�PSETU�P2 {�U~�R�  N �Q��S_AP2BCK� 1|�Y  #�)7Xok%�_8o<P�P&oco9U�_�o o�oBo�o�oxo�o 1C�og�o��, �P�����?� �L�u����(���Ϗ ^�󏂏�)���M�܏ q������6�˟Z�؟ ���%���I�[��� �����D�ٯh���� ��3�¯W��d���� ��@�տ�v�Ϛ�/� A�пe����ϛ�*Ͽ� N���r���ߨ�=��� a�s�ߗ�&߻���\� �߀��'��K���o� ��|��4���X����� ��#���G�Y���}�� ����B���f������1�Y�PP�_ 2>�P*.VR8���*��������l PC���OFR6:�2�V�TzPz�w�]PG���*.Fo/��	�:,q�^/�STMi/ �/ /�-M/�/�H�/?�'?�/�/g?�GIFq?�?�%��?D?V?�?�JPG �?O�%O�?�?oO�
#JSyO�O��5C�O�MO%
JavaS�cript�O�?C�S�O&_�&_�O %�Cascadi�ng Style SheetsR_���
ARGNAMOE.DT�_��� �\�_S_�A�T�_�_>�PDISP*�_���To�_�QLaZoo�CLLB.ZIXwo2o$ :\�a\�o��i�AColla�bo�o�o
TPEINS.XMLƱ_:\![o�QCu�stom Too�lbarbiPA?SSWORDQo��?FRS:\�d�B`Passwor�d Config ���/��(�e��� �����N��r��� ��=�̏a������&� ��J���񟀟���9� K�ڟo�������4�ɯ X��|���#���G�֯ @�}����0�ſ׿f� �����1���U��y� �ϯ�>���b���	� ��-߼�Q�c��χ�� �߽�L���p��ߦ� ;���_���X��$�� H�����~����7�I� ��m���� �2���V� ��z���!��E��i {
�.��d� ���S�w p�<�`�/� +/�O/a/��//�/ 8/J/�/n/?�/�/9? �/]?�/�?�?"?�?F? �?�?|?O�?5O�?�? kO�?�OO�O�OTO�O xO__�OC_�Og_y_ _�_,_�_P_b_�_�_ o�_oQo�_uoo�o �o:o�o^o�o�o) �oM�o�o��6 ��l��%�7�� [����� ���D�ُ h�z����3�,�i� �������ßR��v�������$FIL�E_DGBCK �1|������ < ��)
SUMMA�RY.DG!�͜�MD:U���ِ�Diag Sum�mary����
C?ONSLOG��n����ٯ���Con�sole log����	TPACC�N�t�%\������TP Accou�ntin;���F�R6:IPKDM�P.ZIPͿј
��ϥ���Exception"�ӻ���MEMCHECKЏ�������-�Me�mory Dat�a����:n )��RIPE�~ϐ��%ߴ�%�� Packet L:����L�$�c���S�TAT��߭�� %A�Sta�tus��^�	FTAP����	��/��mment TB�D2�^� >I)ETHERNEw��
�d�u�﨡Et�hernJ�1�fi�guraAϩ��DCSVRF&����7����� verify all:���� 44��DIFF/��'���;�Q�diff��r�d���CHG01������`A����it�2���270���fx�3���I ��p�VTR�NDIAG.LS�u&8���� �Ope��L� ��n�ostic��Y�)VDEV�DAT�������Vis�Dev�ice�+IMG@��,/>/�/:�i$�Imagu/+U�P ES/�/FORS:\?Z=���Updates OListZ?��� �FLEXEVEN���/�/�?���1 ?UIF EvM�M����-vZ)CRSENSPK�/�˞�\!O���C�R_TAOR_PE�AKbOͩPSRB?WLD.CM�O͜�E2�O\?.�PS_ROBOWELS���:GIG��@_�?|d_��GigE�(�O��N�@�)>UQHADOW__D_�V_�_��Shad�ow Chang�e����5dt�RRCMERR�_�_�_�oo��4`CFG �Erroro ta�ilo MA��k�CMSGLIB goNo`o�o|R�e��z0�ic�o�a�)�`ZD0_O�os��7ZD�Pad�l{ �RNOTI��Rd���Not�ific����,�AG��P�ӟt��� ������Ώ]����� (���L�^�폂���� ��G�ܟk� ����6� şZ��~������C� د�y����2�D�ӯ h��������¿Q�� u�
�ϫ�@�Ͽd�v� Ϛ�)Ͼ���_��σ� ߧ�%�N���r�ߖ� ��7���[�����&� ��J�\��߀���3� ����i����"�4��� X���|������A��� ��w���0��=f �����O�s �>�bt �'�K���/ �:/L/�p/��/�/ 5/�/Y/�/ ?�/$?�/ H?�/U?~??�?1?�? �?g?�?�? O2O�?VO �?zO�OO�O?O�OcO �O
_�O._�OR_d_�O �__�_�_M_�_q_o o�_<o�_`o�_mo�o %o�oIo�o�oo�o 8J�on�o��3 �W�{�"��F� �j�|����/�ď֏�e������0��$F�ILE_FRSP�RT  ��������?�MDONLY �1|S�� 
� �)MD:_�VDAEXTP.�ZZZ1�⏹�ț�6%NO B�ack filey ���S�6P�� ���>��K�t����� '���ί]�򯁯�(� ��L�ۯp������5� ʿY�׿ Ϗ�$ϳ�H� Z��~�Ϣϴ�C��� g���ߝ�2���V��� cߌ�߰�?�����u� 
��.�@���d��߈����C�VISBCK�q�[���*.VD�����S�FR:\���ION\DAT�A\��v�S�V�ision VD ���Y�k����y� ��B�����x���1 C��g���,� P����?� Pu�(��^ ��/��M/�q/ �/>/�/6/�/Z/�/? �/%?�/I?[?�/??�?2?D?�?9�LUI�_CONFIG �}S����;O $ �3v�{S� ;OMO_OqO�O�O�I#@|x�?�O�O�O__ %\�OH_Z_l_~_�_'_ �_�_�_�_�_o�_2o DoVohozo�o#o�o�o �o�o�o
�o.@R dv����� ���*�<�N�`�r� �������̏ޏ��� ��&�8�J�\�n���� ����ȟڟ쟃���"� 4�F�X�j�������� į֯����0�B� T�f�����������ҿ �{���,�>�P�b� ���ϘϪϼ�����w� ��(�:�L�^��ς� �ߦ߸�����s� �� $�6�H���Y�~��� ����]������ �2� D���h�z��������� Y�����
.@�� dv����U� �*<�`r ����Q��/ /&/8/�\/n/�/�/ �/;/�/�/�/�/?"? �/F?X?j?|?�?�?7? �?�?�?�?OO�?BO TOfOxO�O�O3O�O�O �O�O__�O>_P_b_ t_�_�_/_�_�_�_�_ oo�_:oLo^opo�o|�o$h  x�o��c�$FLUI_�DATA ~�����a�(a�dRESUL�T 3�ep� �T�/w�izard/gu�ided/ste�ps/Expert�o=Oas���������z��Continue with Gpance�:�L�^� p���������ʏ܏� � �b-�a�e�0 �0`��cl�a?��ps� ��������ҟ���� �,�>�P��0ow��� ������ѯ����� +�=�O�a�?�1�C�U�=e�cllbs�ֿ �����0�B�T�f� xϊϜ�[��������� ��,�>�P�b�t߆߀�ߪ�i�{��ߟ�]�e�rip(pſ-�?� Q�c�u������� ������)�;�M�_� q���������������@������`�e��#pTimeUS/DST	���� ���!3E�?Enabl(�y �������	/P/-/?/Q/�b�`)�/M_q24| �/�/??)?;?M?_? q?�?�?Tf�?�?�? OO%O7OIO[OmOO �O�Ob/t/�/�/Z�~"qRegion�O 5_G_Y_k_}_�_�_�_��_�_�_�America!�#o5oGo Yoko}o�o�o�o�o�o�o��Ay�O�O3�O�_qEditor �o����������+�=� � To�uch Pane�l rs (rec_ommenp�)K� ������Ə؏���� �2�D�|�%���I[qacces oܟ� ��$�6�H��Z�l�~�����Co�nnect to� Network ��֯�����0�B�@T�f�x�����x��@!��}����,!��s �Introduct!_4�F�X�j�|ώ� �ϲ���������� 0�B�T�f�xߊߜ߮�0�������� ɿ ��"�i�{��� ������������/� A� �e�w��������� ������+=�H�3��+�O� ����� 2 DVhz�K��� ���
//./@/R/ d/v/�/�/Yk}�/ �??*?<?N?`?r? �?�?�?�?�?�?��? O&O8OJO\OnO�O�O �O�O�O�O�O�/_�/ 1_�/X_j_|_�_�_�_ �_�_�_�_oo0oBo S_foxo�o�o�o�o�o �o�o,>�O_ !_�E_����� ��(�:�L�^�p��� ��So��ʏ܏� �� $�6�H�Z�l�~���O ��s՟���� �2� D�V�h�z�������¯ ԯ毥�
��.�@�R� d�v���������п� ���ş'�9���`�r� �ϖϨϺ�������� �&�8���\�n߀ߒ� �߶����������"� 4��=��a��Mϲ� ����������0�B� T�f�x���I߮����� ����,>Pb t�E��i���� (:L^p� ������� // $/6/H/Z/l/~/�/�/ �/�/�/����/? �V?h?z?�?�?�?�? �?�?�?
OO.O�RO dOvO�O�O�O�O�O�O �O__*_<_�/?? �_C?�_�_�_�_�_o o&o8oJo\ono�o?O �o�o�o�o�o�o" 4FXj|�M___ q_��_���0�B� T�f�x���������ҏ �o���,�>�P�b� t���������Ο��� ��%��L�^�p��� ������ʯܯ� �� $�6�G�Z�l�~����� ��ƿؿ���� �2� �S��w�9��ϰ��� ������
��.�@�R� d�v߈�G��߾����� ����*�<�N�`�r� ��Cϥ�g���ύ�� �&�8�J�\�n����� ������������" 4FXj|��� �������-�� Tfx����� ��//,/��P/b/ t/�/�/�/�/�/�/�/ ??(?�1U?? A�?�?�?�?�? OO $O6OHOZOlO~O=/�O �O�O�O�O�O_ _2_ D_V_h_z_9?�?]?�_ �_�?�_
oo.o@oRo dovo�o�o�o�o�o�O �o*<N`r ������_�_�_ �_#��_J�\�n����� ����ȏڏ����"� �oF�X�j�|������� ğ֟�����0�� ��u�7�������ү �����,�>�P�b� t�3�������ο�� ��(�:�L�^�pς� A�S�e��ω��� �� $�6�H�Z�l�~ߐߢ� ���߅������ �2� D�V�h�z������ ���������@�R� d�v������������� ��*;�N`r ������� &��G	�k-�� ������/"/ 4/F/X/j/|/;�/�/ �/�/�/�/??0?B? T?f?x?7�?[�? �?�?OO,O>OPObO tO�O�O�O�O�O�/�O __(_:_L_^_p_�_ �_�_�_�_�?�_�?o !o�OHoZolo~o�o�o �o�o�o�o�o �O DVhz���� ���
���_%o�_ I�s�5o������Џ� ���*�<�N�`�r� 1������̟ޟ�� �&�8�J�\�n�-�w� Q���ů������"� 4�F�X�j�|������� Ŀ�������0�B� T�f�xϊϜϮ���� �������ٯ>�P�b� t߆ߘߪ߼������� ��տ:�L�^�p�� ���������� �� $������i�+ߐ��� ���������� 2 DVh'���� ���
.@R dv5�G�Y��}�� �//*/</N/`/r/ �/�/�/�/y�/�/? ?&?8?J?\?n?�?�? �?�?�?��?�O� 4OFOXOjO|O�O�O�O �O�O�O�O__/OB_ T_f_x_�_�_�_�_�_ �_�_oo�?;o�?_o !O�o�o�o�o�o�o�o (:L^p/_ ������ �� $�6�H�Z�l�+o��Oo ��sou����� �2� D�V�h�z������� ����
��.�@�R� d�v���������}�߯ ����ٟ<�N�`�r� ��������̿޿�� �ӟ8�J�\�nπϒ� �϶����������ϯ ��=�g�)��ߠ߲� ����������0�B� T�f�%ϊ������� ������,�>�P�b� !�k�Eߏ���{����� (:L^p� ���w���  $6HZl~�� �s�������/��2/ D/V/h/z/�/�/�/�/ �/�/�/
?�.?@?R? d?v?�?�?�?�?�?�? �?OO���]O/ �O�O�O�O�O�O�O_ _&_8_J_\_?�_�_ �_�_�_�_�_�_o"o 4oFoXojo)O;OMO�o qO�o�o�o0B Tfx���m_� ����,�>�P�b� t���������{oݏ�o ��o(�:�L�^�p��� ������ʟܟ� �� #�6�H�Z�l�~����� ��Ưد����͏/� �S��z�������¿ Կ���
��.�@�R� d�#��ϚϬϾ����� ����*�<�N�`�� ��C���g�i������ �&�8�J�\�n��� ���u��������"� 4�F�X�j�|������� q�������	��0B Tfx����� ����,>Pb t������� /����1/[/�/ �/�/�/�/�/�/ ?? $?6?H?Z?~?�?�? �?�?�?�?�?O O2O DOVO/_/9/�O�Oo/ �O�O�O
__._@_R_ d_v_�_�_�_k?�_�_ �_oo*o<oNo`oro �o�o�ogOyO�O�O�o �O&8J\n�� �������_"� 4�F�X�j�|������� ď֏�����o�o�o Q�x���������ҟ �����,�>�P�� t���������ί�� ��(�:�L�^��/� A���e�ʿܿ� �� $�6�H�Z�l�~ϐϢ� a���������� �2� D�V�h�zߌߞ߰�o� �ߓ��߷��.�@�R� d�v��������� ����*�<�N�`�r� �������������� ��#��G	�n�� ������" 4FX�|��� ����//0/B/ T/u/7�/[]/�/ �/�/??,?>?P?b? t?�?�?�?i�?�?�? OO(O:OLO^OpO�O �O�Oe/�O�/�O�O�? $_6_H_Z_l_~_�_�_ �_�_�_�_�_�? o2o DoVohozo�o�o�o�o �o�o�o�O_�O%O _v������ ���*�<�N�or� ��������̏ޏ��� �&�8�J�	S-w� ��cȟڟ����"� 4�F�X�j�|�����_� į֯�����0�B� T�f�x�����[�m�� ��󿵟�,�>�P�b� tφϘϪϼ������� ���(�:�L�^�p߂� �ߦ߸������� ￿ ѿ�E��l�~��� ����������� �2� D��h�z��������� ������
.@R �#�5�Y��� �*<N`r ��U�����/ /&/8/J/\/n/�/�/ �/c�/��/�?"? 4?F?X?j?|?�?�?�? �?�?�?�??O0OBO TOfOxO�O�O�O�O�O �O�O�/_�/;_�/b_ t_�_�_�_�_�_�_�_ oo(o:oLoOpo�o �o�o�o�o�o�o  $6H_i+_�O_ Q����� �2� D�V�h�z�����]o ԏ���
��.�@�R� d�v�����Y��}ߟ 񟵏�*�<�N�`�r� ��������̯ޯ𯯏 �&�8�J�\�n����� ����ȿڿ쿫���ϟ �C��j�|ώϠϲ� ����������0�B� �f�xߊߜ߮����� ������,�>���G� !�k��Wϼ������� ��(�:�L�^�p��� ��S߸�������  $6HZl~�O� a�s����� 2 DVhz���� ����
//./@/R/ d/v/�/�/�/�/�/�/ �/���9?�`?r? �?�?�?�?�?�?�?O O&O8O�\OnO�O�O �O�O�O�O�O�O_"_ 4_F_??)?�_M?�_ �_�_�_�_oo0oBo Tofoxo�oIO�o�o�o �o�o,>Pb t��W_�{_��_ ��(�:�L�^�p��� ������ʏ܏��� $�6�H�Z�l�~����� ��Ɵ؟꟩��/� �V�h�z�������¯ ԯ���
��.�@��� d�v���������п� ����*�<���]�� ��C�EϺ�������� �&�8�J�\�n߀ߒ� Q������������"� 4�F�X�j�|��Mϯ� q��������0�B� T�f�x����������� ����,>Pb t�������� ����7��^p� ������ // $/6/��Z/l/~/�/�/ �/�/�/�/�/? ?2? �;_?�?K�?�? �?�?�?
OO.O@ORO dOvO�OG/�O�O�O�O �O__*_<_N_`_r_ �_C?U?g?y?�_�?o o&o8oJo\ono�o�o �o�o�o�o�O�o" 4FXj|��� ����_�_�_-��_ T�f�x���������ҏ �����,��oP�b� t���������Ο��� ��(�:����� A�����ʯܯ� �� $�6�H�Z�l�~�=��� ��ƿؿ���� �2� D�V�h�zό�K���o� �ϓ���
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� ������������ ��#���J�\�n����� ������������" 4��Xj|��� ����0�� Q�u7�9��� ��//,/>/P/b/ t/�/E�/�/�/�/�/ ??(?:?L?^?p?�? A�?e�?�?�/ OO $O6OHOZOlO~O�O�O �O�O�O�/�O_ _2_ D_V_h_z_�_�_�_�_ �_�?�?�?o+o�?Ro dovo�o�o�o�o�o�o �o*�ON`r �������� �&��_/o	oS�}�?o ����ȏڏ����"� 4�F�X�j�|�;���� ğ֟�����0�B� T�f�x�7�I�[�m�ϯ ������,�>�P�b� t���������ο��� ��(�:�L�^�pς� �Ϧϸ����ϛ����� !��H�Z�l�~ߐߢ� ����������� �߿ D�V�h�z������ ������
��.����� �s�5ߚ��������� ��*<N`r 1������ &8J\n�?� �c������/"/ 4/F/X/j/|/�/�/�/ �/�/��/??0?B? T?f?x?�?�?�?�?�? ��?�O�>OPObO tO�O�O�O�O�O�O�O __(_�/L_^_p_�_ �_�_�_�_�_�_ oo $o�?EoOio+O-o�o �o�o�o�o�o 2 DVhz9_��� ���
��.�@�R� d�v�5o��Yo��͏� ���*�<�N�`�r� ��������̟��� �&�8�J�\�n����� ����ȯ��я����� �F�X�j�|������� Ŀֿ�����ݟB� T�f�xϊϜϮ����� ������ٯ#���G� q�3��ߪ߼������� ��(�:�L�^�p�/� ���������� �� $�6�H�Z�l�+�=�O� a��������� 2 DVhz���� ����
.@R dv������� ����/��</N/`/r/ �/�/�/�/�/�/�/? ?�8?J?\?n?�?�? �?�?�?�?�?�?O"O ��/gO)/�O�O�O �O�O�O�O__0_B_ T_f_%?w_�_�_�_�_ �_�_oo,o>oPobo to3O�oWO�o{O�o�o (:L^p� �����o� �� $�6�H�Z�l�~����� ��Ə�o珩o��o2� D�V�h�z������� ԟ���
���@�R� d�v���������Я� ����׏9���]�� !�������̿޿�� �&�8�J�\�n�-��� �϶����������"� 4�F�X�j�)���M��� �߅�������0�B� T�f�x������� ������,�>�P�b� t���������{��ߟ� ����:L^p� ������  ��6HZl~�� �����/�� ��;/e/'�/�/�/�/ �/�/�/
??.?@?R? d?#�?�?�?�?�?�? �?OO*O<ONO`O/ 1/C/U/�Oy/�O�O_ _&_8_J_\_n_�_�_ �_�_u?�_�_�_o"o 4oFoXojo|o�o�o�o �o�O�O�O	�O0B Tfx����� ����_,�>�P�b� t���������Ώ��� ���o�o�o[��� ������ʟܟ� �� $�6�H�Z��k����� ��Ưد���� �2� D�V�h�'���K���o� Կ���
��.�@�R� d�vψϚϬϾ�Ͽ�� ����*�<�N�`�r� �ߖߨߺ�y��ߝ��� ��&�8�J�\�n��� �������������� 4�F�X�j�|������� ����������-�� Q������ ��,>Pb !�������� //(/:/L/^// A�/�/y�/�/ ?? $?6?H?Z?l?~?�?�? �?s�?�?�?O O2O DOVOhOzO�O�O�Oo/ �/�/�O_�/._@_R_ d_v_�_�_�_�_�_�_ �_o�?*o<oNo`oro �o�o�o�o�o�o�o �O_�O/Y_�� �������"� 4�F�X�o|������� ď֏�����0�B� T�%7I��mҟ �����,�>�P�b� t�������i�ί�� ��(�:�L�^�p��� ������w��������� $�6�H�Z�l�~ϐϢ� ���������ϻ� �2� D�V�h�zߌߞ߰��� ������
�ɿۿ�O� �v��������� ����*�<�N��_� �������������� &8J\�}?� �c�����" 4FXj|��� ����//0/B/ T/f/x/�/�/�/m�/ ��/�?,?>?P?b? t?�?�?�?�?�?�?�? O�(O:OLO^OpO�O �O�O�O�O�O�O _�/ !_�/E_?	_~_�_�_ �_�_�_�_�_o o2o DoVoOzo�o�o�o�o �o�o�o
.@R _s5_��mo�� ���*�<�N�`�r� ������gȍޏ��� �&�8�J�\�n����� ��c��џ���"� 4�F�X�j�|������� į֯������0�B� T�f�x���������ҿ �������ٟ#�M�� tφϘϪϼ������� ��(�:�L��p߂� �ߦ߸������� �� $�6�H���+�=ϟ� a���������� �2� D�V�h�z�����]��� ������
.@R dv���k�}������$FMR2_GRP 1���� �C4  B��	 ��9K6/F@ a@�6�G�  �Fg��fC�8R�y?ǀ  ��66��X���875t���5���5`{+�yA�  /�+BH�w-%@S339%�5[/l-6@6!�/xl/�/�/ �/�/?�/&??J?5?�G?�?k?�?��_C_FG �TK��?�? OO�9NO {
F0FA� K@�<RM_CHKTYP  ��$&� ROM�a@_MINg@������@�R XS�SB�3�� 7�O���C��O�O�5TP_DEF_OW  ���$WIRCOM�f@_�$GENO�VRD_DO�F̾�E]TH��D dzbUdKT_ENB7_{ KPRAVCu��G�@ �Y �O�_�?oyo&onI* �QOU�NAIRI<�@��oGo�oX�o�o��C�p3���O:��B��+sL�i�O�PSMT���Y(�@
t�$�HOSTC�21���@�5 kMC��R{����  27.0z0�1�  e� ]�o�������K�ď֏���������	anonymous!� O�a�s����� �4��������D�!� 3�E�W�i��������� ï柀�.���/�A� S���课�П���� Ŀ����+�r�O�a� sυϗϺ������� ��'�n��������� ��ڿ����������F� #�5�G�Y�k���υ� ����������B�T�f� C�z�g��ߋ������� �����	-P��� ��u������ (�:�<)p�M_q ��������/ $ZlI/[/m//�/ ����//�/D!? 3?E?W?/?�?�?�? �?�/�?./OO/OAO SO�/�/�/�/�?�O? �O�O__+_r?O_a_ s_�_�_�O�?O�_�_�oo'o�t�qENT� 1�hk P!\�_no  �p\o �o�o�o�o�o�o�o �o:_"�F� j�����%�� I��m�0���T�f�Ǐ ��돮��ҏ3���,� i�X���P���t�՟�� ៼�
�/��S��w� :���^�������������ܯ=� �QUI�CC0J�&�!1�92.168.1'.10c�X�1��v�8��\�2�ƿؿ9��!ROUTER�:��!��a���PCJOG��e�/!* ��0��U�?CAMPRT�϶�c!�����RTS����x� !So�ftware O�perator PanelU߇����7kNAME !~Kj!ROBO�����S_CFG 1��Ki ��Auto-st�arted�DFTP�Oa�O�_�� �O����������E_� .�@�R�u�c�	����� ������cN:�L�^�; r���R������ ��%H�[ m���jO|O�O �O4!/hE/W/i/{/ �/T�/�/�/�/�// �//?A?S?e?w?�?� ���??�?</O+O =OOO?sO�O�O�O�O �?`O�O__'_9_K_ �?�?�?�?�O�_�?�_ �_�_o#o�OGoYoko }o�o�_4o�o�o�o�o f_x_�_g�o� �_�����o�� -�?�Q�tu������ ��Ϗ�(:L^`� 2��q����������� ݟ���%�H�ʟ[� m����������� � ί4�!�h�E�W�i�{� ��T���ÿտ�
�� ��/�A�S�e�w����_ERR �����ϗ�PDUSIZW  �^6�����>��WRD ?�(����  guestƀ��+�=�O�a���S�CD_GROUP� 3�(� ,��"�IFT��$PA��OMP�� n��_SH��ED��w $C��COM���TTP_AUTH� 1��� <!�iPendan�m�x�#�+!KAREL:*x���KC�������VISION SET��(����?�-�W�R���v������������������G�CT_RL ���a��
��FF�F9E3��F�RS:DEFAU�LT�FAN�UC Web Server�
td G����/� 2�DV��WR_CONFIG ��՗�����I�DL_CPU_P5C� �B����w BH�MIN�����GNR_IO������ȰHMI�_EDIT ���
 ($/C/�� 2/k/V/�/z/�/�/�/ �/�/?�/1??U?@? y?d?�?�?./�?�?�? �?OO?OQO<OuO`O �O�O�O�O�O�O�O_�_;_�NPT_S_IM_DO�*�NSTAL_SC�RN� �\UQT�PMODNTOL8�Wl[�RTYbX��qV�K�ENB�W��ӭOLNK 1�����o%o7oIo�[omoo�RMAST�E��Y%OSL?AVE ��Ϯe�RAMCACHE��o�ROM�O_CF1G�o�S�cUO'�~�bCMT_OP� 8 "��5sYCL�ou�� _ASG 1����
 �o�� �����"�4�F��X�j�|����kwrNU�M����
�bIP��o�gRTRY_C�N@uQ_UPD��a��� �bp�b���n��M��аP�}T?��k �� ._������ɟ۟퟈S ���)�;�M�_�q� � ������˯ݯ�~�� %�7�I�[�m������ ��ǿٿ�����!�3� E�W�i�{�
ϟϱ��� �����ψϚ�/�A�S� e�w߉�߭߿����� ����+�=�O�a�s� ���&��������� ���9�K�]�o����� "������������� ��GYk}��0 �����C Ugy��,>� ��	//-/�Q/c/ u/�/�/�/:/�/�/�/ ??)?�/�/_?q?�? �?�?�?H?�?�?OO %O7O�?[OmOO�O�O �ODOVO�O�O_!_3_ E_�Oi_{_�_�_�_�_ R_�_�_oo/oAo�_ �_wo�o�o�o�o�o`o �o+=O�os �����\n� �'�9�K�]�����������ɏۏi�c�_M�EMBERS 2��:�  � $:� ����v���1���RC�A_ACC 2��� �  [�  )��s ]� ��` 6>@l��l��)B� �9p����  il����a�BUF001 �2�n�= �.�u0  u0�:��H�T�b�nz�{�  8���  ���Vu0��eJ�s�J��J��J��J���J��J��J��J��VJ������(���7��J��Yu0p����gu0(��L��tu0aohȽa�������������u0.�PF������u0_p�������u0	`k�{���0u ���V��2� 2�,2�U82�F2�R2�`2�Ul2�x2��2��2�Tq�4��2��2��2�U�2��2��2����	��#�ߙ2 ��������� �!��)��1��8� :�@�B�H�Z�l�~���ࢯ��ƣ��ѡ8L��ءc�p��-��G��a�h��@i�(�{p 0��p88�xJ�\�n��Y���t� x�����������ҡ��ҩ�u  x���ҹ�s�8�� ��ɰ�Ѱ�ٰ���ߙ3������� ��!�/��1�?�l� A�O�V�Z�V�b�V�j� V�r�V⑲�V��V� ��V��V��l����� ��������������� ɠ��Ѡ��٠��s��� �������������	� ��������!���)� l�0���Bҗ�Jҗ�R� ��Zҗ�bҗ�jҗ�r� ��q���y��Ё��Љ� ��>򙲧�>򩲗б� ��>������Ѳ�����ݖCFG 2��n� 4G�l�
l�<l�47M�a��HIS钜n� ��� 2025O-12-�l��� # )珢� ���� 2��ׁ�{q1}	6�4m���h   7 pD���xl�;s�14 ��l�7 ��9 ����������C�3 	 U��{ � *[~�qq1-3E����� &f  �' "�b/t/  P�X�`�����  �  $  >� 8 ����������� , (!�  8C�� d{�q4[}�R)'29}?1?C?U?g?�y?�?�?h�( %� C� -�RO  *C l��<B��?OO*O<ONO `OrO�O�O�O�?�?�O �O__&_8_J_\_n_ �_�O�O�_�_�_�_�_ o"o4oFoXoٚS���[m
-  L _o�o�o�o�o!3 EWEW7d\������ _�%C >��"��"��r>�  3��"���r �" �"C�:��a .�a%/7*8
 cI 8��"y����y/�s� �r� �r�+�  X� �X*�|c�,: J��"��0  Q�1� 
 R*�: b�(=�`??I�[�m���������ǟ�8�cH |9�,��01�\�_�_%�7�I�[�m� �������ǯ�_��� �!�3�E�W�i�{��� ��֯诬������ /�A�S�e�w�eowc���o�o
i������� �0�B�T�f�x�fxe3�����������rI:�q�pB�q�D�qB�H�q
�*��I�q�J�q�B�*�B� B��V��{��J�7*	
�qI �ߨ��& �� �⾀���p���p�G�+��2�;�C� "&� .[�6�� ��&�8�n� ���������������:T�[��0f���п N`r����� ��'9&8J\ n������ �/"/4/F/X/j/|/��/�/��I_CFG� 2��� H�
Cycle T�ime�Bus=y�Idl�"��min�+1�Up�&�Re�ad�'Dow�8?>� 1�#Co�unt�	Num	 �"����<�p�qaPROG�"힦����)/�softpart�/genlink�?current�=menupage,1133,}w�OO&O8O<b5leS�DT_ISOLCW  ���Ҁ�/�J23_DSP_�EN�vK0�@INC ��M�s�@�A   ?�=�?��<#�
�A�I:�o��N_�tX�O<_�GOB�0C�C���1�FVQG_GR�OUP 1�vK%�<��C�y�_D_?�x�?�_�pQ�_o.o@o�_dovoȈo�o�w,_NYG_IN_AUTO��>�MPOSRE^_pV�KANJI_MA�SK v�HqREL?MON ��˔?�ry_ox����(�.6r�3��7�C����u�o�DKCL_�L�`NUM��E�YLOGGING�������E�0LA�NGUAGE ���~��DEFAULT ��6��LG�!��:2k�� 80�2ଊ�'~�  �W 
��ћ��GO�UF ;��
��(UT1:�� � �-�?�Q�h�u����������ϟ�����(�g4�8i�N_DISP ��O8�_��_��LOCTOL����Dz A�A���GBOOK ����d�1
�
�۠ ������#�5�G�Y�`i���3{�W�	��@쉞QQJ¿Կ1���_BUFF 2��vK ������
�ڢVB&�7 C�ollaborativ�=�OΗώ� �ϲ���������'�� 0�]�T�fߓߊߜ��?DCS ��9�B �Ax���Rh�%�-�?�|Q���IO 2���� ���Q� ������������ �*�<�N�b�r����� ����������&�:e�ER_ITMsNd�o����� ��#5GYk }����������hSEV�`�M.dTYPsN�c/pu/�/
-�aRST5����SCRN_FLW 2�s��0��� �/??1?C?U?g?�/�TPK�sOR"��NGNAM�D��~�N�UPS_ACR� ��4DIGI�8~+)U_LOAD[P�G %�:%T_NOVICEt?���MAXUALR�M2��a���E
LZB�1_P�5�` ��4y�Z@CY��˭�O�+���ۡ�D|PP 2]�˫ �Uf	R/ _
_C_._g_y_\_�_ �_�_�_�_�_�_oo ?oQo4ouo`o�o|o�o �o�o�o�o)M 8qTf���� ���%��I�,�>� �j�����Ǐُ���� �!���W�B�{�f� ������՟����ܟ� /��S�>�w���l��� ��ѯ��Ư��+���O�a�D���p���RHD�BGDEF ��E�ѱO��_LDX�DISA�0�;c�M�EMO_AP�0E� ?�;
  ױ��3�E�W�i�{ύ���ϱ�Z@FRQ_C_FG ��G۳�A ��@��Ô�<��d%�� ������Bݯ�K���*i�/k� **:tҔ�g�y�ߔ��� �����������J� ���Es�J d������,(H���[���� �@�'�Q�v�]����� ����������*�NPJISC 1��9Z� ������ܿ������	Zl_MSTR �#-~,SCD 1�"��{����� ���//A/,/e/ P/�/t/�/�/�/�/�/ ?�/+??O?:?L?�? p?�?�?�?�?�?�?O 'OOKO6OoOZO�O~O �O�O�O�O�O_�O5_  _Y_D_i_�_z_�_�_ �_�_�_�_o
ooUo @oyodo�o�o�o�o�o �o�o?*cNl�MK���;�љ$MLTAR�M���N��r� ��հ��İM�ETPU��zr���CNDSP_A�DCOL%�ٰ0�C�MNTF� 9�F�Nb�f�7�FSTLqI��x�4 �;�ڎ�s����9�PO�SCF��q�PR�PMe��STD�1ݶ; 4�#�
v��qv�����r��� �����̟ޟ ��� V�8�J���n���¯������9�SING_CHK  ���$MODA����t�{�~2�DEV �	�	MC:>f�HSIZE��zp��2�TASK �%�%$1234?56789 ӿ��0�TRIG 1�; lĵ�2ϻ�0!�bϻ�YP�����H�1�EM_IN�F 1�N�`�)AT&FV0�E0g���)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ��2��H6� ^���Rφ��A�߶� q�������� ��5� �����ߏ�B߳��� ��������1�C�*� g��,��P�b�t��� ���R�?���u 0��������� ������M q�� �Z���/�%/ ��[/ 2�/�/ h�//�/�/�3?�/ W?>?{?�?@/�?d/v/ �/�/O�//OAOx?eO ?�ODO�O�O�O�O_��NITORÀG �?z�   	�EXEC1~s&R2*,X3,X4,X5,X���.V7,X8,X9~s 'R�2�T+R�T7R�TCR �TOR�T[R�TgR�TsR��TR�T�R�S2�X2��X2�X2�X2�X2��X2�X2�X2�X2*h3�X3�X37R2��R_GRP_SVw 1��� (�q�>�����F��=5�[����濢c�a���_D�B���cI_ON_DB<��@��zq  �zpORzpPY�1u�zp�>w+�ZpZpY��@�N �p{�p|>{���p5q�r-ud�1�����8�PG_JOG �ʏ��{
�2�:��o�=���?����0�B��~\�n��������H�?��C�@�ŏ׏����  �����qL�_NAME !�ĵ8��!De�fault Pe�rsonalit�y (from �FD)qp0�RMK_ENONLY��_�R2�a 1�L�XL�8�gpl d����ş ן�����1�C�U� g�y���������ӯ� ��	����
�<�N�`� r���������̿޿� :��)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+��<�Sew����������A�a��B�Bw��Pf���� ��/!/3/E/W/i/ {/�/�/�/���/�/ ??/?A?S?e?w?�? �?�?�?�?�?�?�/�/ +O=OOOaOsO�O�O�O �O�O�O�O__'_9_0&O�S���x_�]�rdtS���_�]�_�_ �W�����S"oe_oXoa ��qogoyo �o�o�o�o�ouP�p4"|����	`[oUgy8qK�A\����s� A ��y@hT�Q�Q��"���T�k\$��  ���P�PE�xC�  �I�@oa� <o��p�������ߏ
f��Q*�����0��P�Cr� � �3r �.� @D� M A�?�G�-�?.<I�.@I�A���~�  ;�	lY��	 �X  ������� �, �� �����uPK�o������]K���K]�K	�.��w�r_	����@
�)�b�1������I�Y������T;fY�{S=���3����I��>J���;Î?v��>��=@����	�E��RѯעZ��p�wp��u�� D!��3��7pg  ?�  �9�͏�W���	'� �� u�I� ��  ��u��:��È��È=��9ͱ���@��ǰ �3��\�3�E�&����N�pC�  ' Y�&�Z�i�b�@f�i�Fn�C����I�C��4��b��r��!�`����B�p����q���}ر�.Dz Ə<ߛ�`�K�pߖ���w������А 4P�����.z��d  ��Pؠ?�ff0�_��	�� 2p>��P���8.f�t�>L����U���(.��P���������
ĉ��� �x��;e�m���KZ;�=g;�?4�<<�����%�G��3����p?offf?ذ?&S����@=0e�?��q�+�rN�Z��� I���G���7���(��� ��!E0iT�`���+��F�p ���#��D�� w������ �//=/(/a/L/�/ p/��/�p�6�/Z #?�/ ?Y?k?}?��? �?>?�?�?�?�?�?1OD�����KD�y^KCOp�OO�O���ذO��O�O�Oai���J��}�DD1���.�D���@�AmQa��9N,�ȴA;�^@���T@|j@$��?�V�>��z�ý��=#��
>\)?���
=�G�-]��{=���,���C+��Bp��P��6��C�98R���?�N@��(��5���-]G�p�Gs�b�F�}�G��>.E�VD��Kn���I��� F�W�E���'E���D���;n���I���`E�G���cE�vmD���-_�oQ_�o�o�o  �o$H3X~ i������� ��D�/�h�S���w� �������я
���.� �R�=�v�a�s����� П����ߟ��(�N� 9�r�]���������ޯ ɯۯ���8�#�\�G� ��k�������ڿſ�� �"��F�1�C�|�g� �ϋ��ϯ��������z�P(�Q34�] �����Q�	�9�Oߵ5�3~�mm��aҀ�5Q�߫�aғ�x���ߵ1����� ��1��U�C�y�g��%%P�P���!�/���'���
���.������4�;�t�_����� ����������:�%��/�/d�������� 7%[Im���027�  B�XS@J@�CH#PzS@�0@ZO/1/C/U/g/y/�-�#��/�/�/��/�/�3?�3�� U@�3��0�0�13��5
  ?f?x?�?�?�?�?�? �?�?OO,O>OPO�Z�@1 ���ۯ�c�/�$MR_CA�BLE 2ƕ�_ ��TT�� ���ڰO���O�)�@�� �C_���_O_u_7_ I__�_�_�_�_�_o �_�_oKoqo3oEo{o �o�o�o�o�o�o�o�o Gm/�K!�"���O����ذ��$�6���*Y�*�* �COM ���I����  ��)�%%� 2345678'901���� ��Ï���� � !� �!
���Mn�ot sent �b��W��T�ESTFECSALGR  eg�*"!d[�41�
k�������$pB����������� 9UD�1:\maint�enances.�xmlğ���C:��DEFAUL�T�,�BGRP 2��z�  �� O���%  �%!1�st clean�ing of c�ont. v�i�lation 56��ڧ�!0�����+B��*������+��"%��mec�h��cal ch�eck1�  �Bk�0u�|��ԯ�����Ϳ߿�@���rollerS�e�w�ū��m�ϑϣϵ��@�Basic �quarterl!y�*�<�ƪ,\�)�`;�M�_�q�8�MJ�,�ߓ "8��� ���ߕ �����+�=��C�g�ߋ�ʦ�߹��������@��Overhaul�ߔ��?� x� I�P����}���������� $n������ �)l�ASew��� ��� �+ =O�s���� ���/R�9/� (/��/�/�/�/�// �/�/N/#?r/G?Y?k? }?�?�/�???�?8? OO1OCOUO�?yO�? �?�O�?�O�O�O	__ jO?_�O�Ou_�O�_�_ �_�_�_0_oT_f_;o �__oqo�o�o�o�_�o o,oPo%7I[ m�o��o�o�� ��!�3��W��� �����ÏՏ�6��� �l����e�w����� ����џ�2��V�+� =�O�a�s������ ͯ����'�9��� ]�������⯷�ɿۿ ���N�#�r���YϨ� }Ϗϡϳ������8� J��n�C�U�g�yߋ� �ϯ������4�	�� -�?�Q��u������� ����������f�;� ������������� ���P���t�I[ m������ :!3EW�{ ��� ���/ /lA/��w/��/��/�/�/�/X*�"	 �X�/?.?@?�)B  a/o?m/o%w?�?�?}? �?�?OO�?�?OOaO sO1OCO�O�O�O�O�O __'_�O�O]_o_�_ ?_Q_�_�_�_�_�_�\� Џ!?�  @�! M?HoZo�lo�&4o�o�o�o�(�*�o** F�@ �Q�V�`o'�9�o]o�����/^&�o���� �/�A�S�e���#� ����я�����+� q�����7�������k� ͟ߟ��I�[���K� ]�o���C�����ɯ���o$�!�$MR�_HIST 2���U#�� 
 \�7"$ 23456789013�;��
�b2�90/����[� ��./����ǿٿF� X�j�!�3ρϲ���{� �ϟ�����B���f� x�/ߜ�S����߉��� ���,���P��t���=��$�SKCF�MAP  �UK&��b
�� �����ONREL  �$#������EXCFENB�q
����&�FNC-���JOGOVLI�M�d#�v���KE�Y�y���_P�AN������RU�Ni�y���SF?SPDTYPM�����SIGN��TO1MOTk�����_CE_GRP 1��U��+�0 �ow�#d��� ���&�6\ �7y�m�� �/�4/F/-/j/!/ t/�/�/�/{/�/�/�/�?�+��QZ_ED�IT
����TCO�M_CFG 1����0�}?�?�? 
>^1SI �N�!���?�?���?$O�����?XO78T_/ARC_*�X��T_MN_MOD�E
�U:_SP�L{O;�UAP_C�PL�O<�NOCH�ECK ?�� �� _#_5_ G_Y_k_}_�_�_�_�_��_�_�_oo��NO_WAIT_L	lS7> NTf1�����%��qa_ERR&H2�������?o�o�o�o��OGj�@O�cӦm|)���GAA�Y����[��2#�@�"� Nl�,��<���?����)��n�bP�ARAM�b����tGO�8
�.�@� = n�]�o� w�Q�����������`Ϗ�)��7�[��m� �����ODRD�SP�C8�OFFSET_CARI0��OǖDISԟœS;_A�@ARK
T9�OPEN_FIL�E��1T6�0OPTION_IO�����K�M_PRG ;%��%$*�����'�WO��N�s�ǥ�� ���u����	� ����Ӧ������RG_DSBL'  ����jN����RIENTTO����C�����A� ��U�@IM_D�S���r��V��LCT �{mP2ڢȪ3̹��dҩ��_P�EX�@���RAT��G d8��̐UOP װ�:�����S�e�Kωϗ��$��r2G�L�X�LȚ�l 㰂�������'�9� K�]�o߁ߓߥ߷��� �������#�5�G���2��v������� ������e�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?�q1�~?�?�?�? �?�?�?�?O O2ODO�yA�a�tn?~M��~O�O�P�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�O�O o$o6oHoZolo~o�o �o�o�o�o�o�o  �_oVhz��� ����
��.�@�`R�d�QOES������B�d�ӏ�ʏ ��������Y�D�}�0��r��������� ԟڟ���p���=�M��q�	`������<��c�:�o�¯�ԯ����A� � �k�C�C�ڰ"�ڰ���O�_�  ���-����)�C�  � t�k���g�����Կ���ѿ
�5���_:�ĳ�O�U���6���6�H��n��� � ^�~\� @D�  p�?�v�\�?:px�:q�C4r�p�(��  �;�	l��	 ��X  ������� �, � ��������Hʪ�����H���Hw��zH���ϝ�8�B���B� � Xѐ�`�o�*��3����t�>u���fC�{ߍ��:pB\�
��Ѵ9:qK	�t�� ����p$���*��� DP��^��b�g  ?�  �h������)�	'� �� ��I� ��  ��'�=��������t�@�����!�b��^;b��t�U�(�N��r�  '��E�C�И�t�C�И��ߗ���jA�@C�����%�B��� ��,���H:qDz�k�ߏz���������А 4P����:uz:���	�f��?�ff0'�&8� ]�m��8:p��>L������$�(:p�P ��	������:�{ x�;e�m"��KZ;�=g;�4�<<���E/Tv��b����?fff?�?&�� )�@=0�%?��%_9��}!�� $�x��/v��/f'��W ,??P?;?t?_?�?�? �?�?�?�?O�?(OO LO�/�/�/EO�OAO�O �O�O�O_�O_H_3_ l_W_�_{_�_�_1��_ A���eO+o�ORooOo �o�o�oK/�o�omo��o*'`+�,�zt���CL�H��}?�����,
������u���F�D1�/n�t��p��q��@I�h~,�ȴA;�^@���T@|j@$��?�V�n��z�ý��=#��
>\)?���
=�G�����{=��,���C+��Bp���6��C�98R���?�}p��(��5�����G�p�Gs�b�F�}�G��>.E�VD��KL����I��� F�W�E���'E���D���;L����I���`E�G���cE�vmD���\�՟��ҟ��� /��S�>�w�b����� ��ѯ�������=� (�:�s�^��������� ߿ʿ�� �9�$�]� Hρ�lϥϐϢ����� ����#��G�2�W�}� hߡߌ��߰������ ��
�C�.�g�R��v� ��������	���-� �Q�<�u�`�r����� ��������'Mz�(�34�]O!���8h~�%�3~�m�����5Q�����x��!���   `N�r��	e%P@"P��Q�_/�V/9/$/]/H)����c/j/�/�/�/�/ �/�/�/!??E?0?i?�T?"&�_�_�?�?�8��?�?O�?OBO0O fOTO�OxO�O�O�O�O�2f?_  B�X�pyp$QCHR�z�p@�N_`_r_�_�_�_�]c�O�_�_o�o+o?�Bc� U@d4��QJc�D
  2o�o�o�o�o�o�o %7I[m���oa �����c�/�$PARAM�_MENU ?� � � DEFP�ULSE��	W�AITTMOUT��{RCV� �SHELL_W�RK.$CUR_oSTYL�p"��OPT8Q8�PTB�M�G�C�R_DECSN�p������� �������-�(�:��L�u�p��������qS�SREL_ID � ��̕US�E_PROG �%�z%���͓CC�R�pޒ��s1�_H�OST !�z!6�s�+�T�=����V�h���˯*�_TGIME�rޖF��p?GDEBUGܐ�{�͓GINP_FLgMSK��#�TR2��#�PGAP� ���_b�CH1�"�TY+PE�|�P���� ����0�Y�T�f� xϡϜϮ��������� �1�,�>�P�y�t߆� ���߼�����	���(�Q�L�^�p��%�W�ORD ?	�{
? 	PR�p#�MAI��q"SUd���TE��p#��s	1���COLn%h��!���L�� !՜�F�d�TR�ACECTL 1�� �q ��{ |#�����_�DT Q�� ��z�D ȿ � K` ��c`��_`�������� ��1CUgy �������	 -?Qcu�� �����//)/�;/M/ � b �@P"M`P"k`P" ��h/z/�/�/�/�/�/ �/�/
??.?@?R?T/ ~?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_�_��Z5oo*o <oNo`oro�o�o�o�o �o�o�o&8J \n������ ���"�4�F�X�j� |�������ď֏��� ��0�B�T�f�x��� ������ҟ����� ,�>�P�b�t������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�.�oP� b�tφϘϪϼ����� ����(�:�L�^�p� �ߔߦ߸������� � �$�6�H�Z�l�~�� ������������ � 2�D�V�h�z������� ��������
.@ Rdv����� ��*<N` r������� //&/8/J/\/n/D� �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�? �?�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� � 2�D�V�h�z�����������$PGTRA�CELEN  ���  ������Ά_UP �����������΁_�CFG ����烸�
���*��:�D�O���O�  ��O��DEFS_PD ��������΀H_CONFIG ����� ����d�Ĕ�݂ ��ǑP�^�a�㑹��΀I�N�TRL �d�=�8^���PE��;೗���*��ÑO�΀LID����	T�LLB 1}ⳙ ���BӐB4��O� �䘼����Q� �<< ��?� ������M�3�U� ��i���������ӿ��	�7�T�Ϣk�b� tϡ�诚��������~S�GRP 1爬����@A!����4I���A ��Cu�C�O_CjVF�/���Ȕa�zي�ÑÐ��t��ޯs���´�ӿߨ�B������������A�S�&�B34�_������j�������� �	�B�-���Q���M�x������  Dz�� ��.�����&L7 p[��������6!Zh)�w
V7.10_beta1*�Ɛ�@�*�@�) @�+A Ē�?��
?ff�f>����B�33A�Q�0�B�(��A���AK��h�����//'/9/P�p*��W�ӑ�n/�/�%����R�fh����*���P2�LR� �/�/�/�/�/H?�Ĕ	�I�u�&:���? ��x?�?A���P!\3� Bu�B��?�5B)H�3[4��o��4&��[45��/B\3x3Dx�?YO�?aOkO}O�<<�R@��O�C��O�O�O�O�DA�X�K�NOW_M  �Z�%�X�SV ���ڒ���_�_ �_?�_�_�_o�����W�M+�鳛 ���	@�3#����_�o�\A��
7]bV4�@u���u��e�o�l,�X�MR
+��JmT3?��W�1�C{�OADBANgFWDL_V�ST+ѯ1 1����P4C���[��i/� ����?�1�C��� g�y��������ӏ� *�	��`�?�Q�c��w�2�|Va�up�<ʟ���p3��Ɵ؟Ꟃ�w4��+�=��w5 Z�l�~����w6����ѯ㯂w7 ��$�6���w8S�e�w����wM�Amp������O�VLD  ���yo߄rPARNUM  �{+þ�?�n�qSCH�� ��
��X���{s��UP�DX�)ź��Ϧ�_C�MP_@`���p|P'�yu�ER_CHK���yqbb3֌�.�RSpp?Q_�MOm��_}ߥ�__RES_G�p쩻
�e�����0�#�T� G�x�k�}�������@�������׳����� ����:�Y�^���Y� y������Ӭ������� ��������R�6 UZ�ӥ�u���ҏV 1�FvpVa�@k�p��THR_INRp��(byu�dMASS �Z)MNGMO�N_QUEUE C�uyvup\!��N�UZ�NW���END��߶EX1E����BE��>�OPTIO�����PROGRAM7 %z%���~ϘTASK_I���.OCFG ��z+�n/� DAT�ACc�+@ ��KP@2 �??/?A?S?]51 s?�?�?�?�?�6 p1�?�?�?O"O,F�!�INFOCc��-� �bdlO~O�O�O�O�O �O�O�O_ _2_D_V_ h_z_�_�_�_�_�_�/4A@FD��, 	��!6��K_�!�)fN!fENB��0m��Pfi2YokhG�!2�0k X,		d�o=��·o���e�a$�pd��i�i�g�_EDIT ��/%7����*S�YSTEM*upV�9.40107 �cr7/23/2021 A���Pw��PRGAD�J_p  h �$X[�p $Y�xZ�xW�xқt�ZқtSPEED_��p�p$NEXT�_CYCLE�p����q�FG�p� ��pALGO�_V �pNYQ�_FREQ�WI_N_TYP�q)��SIZ1�O�LA!P�r!�[��M+�����qCREATED��r�IFY�r@!N�AM�p%h�_G>J�STATU��J��DEBUG�rMA�ILTI����E�VEU��LASTx�����tELEM�� � $EN�AB�rN�EASI�򁼁AXIS�p�$P߄�����qR�OT_RA" �rM�AX ��qE��L�C�AB
���C D�_LVՁ`�BAS ��`�1�{���_� ��g$x���RM� 9RB�;�DIS�����X_SPo�΁�� ��u�P� | �	� 2 6\�AN�� �;������Ӓ�� |�0�PAYLO��<3�V�_DOU�qS�x��p�tPREF�� ( $GR�ID�E
���R����Y��rOTO|ƀ�q  �p℄!�p��k�OXY�� � $L��_PO|�נVa.�SRV��)����DIRECT_1T� �2(�3(�4(�U5(�6(�7(�8���qF��A�� �$VALu�GR�OUP������/� !��@!⾣�����RAN�泲���R��/���T�OTA��F��P�W�I=!%�REGEN#�8�������/���ڶnTzЉ����#�_S����8�(�V�[�'���4���GRE��w���H��D�����wV_H��DAY3�V��S_Y�Œ;��SUMMAR��2� $CONFIG_SEȃ���Nʅ_RUN�m�C�о��$CMPR���P�DEV���_�I��ZP�*��q��E�NHANCE�	��
���1���INT��qM)b�q�r2K����OVRo�PGu�IX��;����OVCT�����v�
 4 ����a˟���PSLG"�� \ �;��?��1���SƁϕc��U�����Ò�4�U�  [�Tp�� (`�-��rJ<�Oz� CK�IL_MJ�b��VN�+��TQn�{�N5���C�UL�ȀD�V(�C6�P_h�຀@�MW�V1V��V1d�2s�2d�3*s�3d�4s�4d���'�	�������p	�I=N	VIB1qp1�B 2!pq/,3 3,4 4,�p?� �;��A���N��������PL��TOR�r3�	��[�SA�V��d�M�C_FOLD 	$SL���Պ�M,�I��L� ��pL�b��KEEP_HNADD	�!Ke�UCCOMc�k��
�lOP���pl��.lREM�k��P΢���U��ek�HPW� KS�BM��ŠCOLL�AB|�Ӱn��n��+�IT�O��${NOL�FCALX� �DON�r����o ,��FL�>��$SYNy,�M�C=����UP�_DLY�qs"DGELA� ����Y(��AD��$TAB�TP_R�#��Q�SKIPj% ����OR� �E�� P_��� �)���p 7��%9��%9A�$:N� $:[�$:h�$:u�$:���$:9�q�RA��� X�����MB>�NFLIC]��0�"�U!�o���NO_�H� �\�< _SW�ITCHk�RA_�PARAMG�� ��p��U��W�J��:Cӣ�NGRLT� OO�U�����8X�<A��T_Ja1F��rAPS�WEIG=H]�J4CH�aDcOR��aD��OO���)�2�_FJװ���sA0�AV��C�HOB.�.�N`�J2�0�q$��EX��T$�'QIT ��'Q�pG'Q-�GA�DC�m" � ��<��
R]��
H�<��RGEA��4��U�FLG`g��H���ER	�SPC�6R�rUM_'P��2�TH2No��@Q 1 ���0�����  D q�وIi�2_P�2�5cS�ᰁ+�L10_CI��pe� �pk����U ՖD��zaxT�p�Q(�;a��c��޲+��i���e��` P>`DESIGRb$�VL1:i1Gf�c�g;10�_DS��D�|Qw�POS11�q l�pr��x1C�/#AT�B��U
WusIND��}�mq�Cp�mq`B	�HOMME�r 	aBq2Gr�M_q��� )@Ar3Gr��@� ��$�`!@s4GrG�Y�k�}�������
?t5Grď֏���(����6GrA�S��e�w������w7Gr���П�������8Gr;�M�_�q������6�S �q    �@sM��P�!�K@��! T`M��&M�IO��m�I��2�OK _OPy��� �ػQ�2�pWE"� 7�x EQWQE� � #s%Ȳ$D;SBo�GNA�b� C�P2�<rS23�2S�$ �iP���xc�ICE<@%�P1E`2� @IT��P��OPB7 1�FLO�W�TRa@2��U�$�CUN��`�AUX�T��2Ѷ�ERFA�C3İUU����K�SCH��% �t<_9�EЎA�$FREEFRO	MЦ�A�PX q��UPD"YbA�PT�.�pEEX0����!��FA%bҸp�R�V�aG� & � ��E�" 1�AEL�  �+�jc'���D�  2& ��S\PcP(
  �	$7P�%�R�2� ���T�`AXU���DSP���@�W���:`$���RNP�%�@����K��_MIR�����3MT��AP��0�P"�qD�QSYz������QPG7�BRKqH���ƅ AXI�  ^��i���1x ����BSOC����N��DUMMY{16�1$SV��DE��I�FSPD/_OVR79� �D����OR��֠N�"`��F_����@OVv��SF�RUN�b�"F0�����UF"@vG�TOd�LCH�">�%RECOV��9@�@W�`&�ӂH��r:`_0��  @�R�TINVE��8AO�FS��CK�KbFWD������1B���TR�a�B �FD�� ��1= B1pB�L� �6� A1L�V ��Kb����#��@+<�AM:��0��j���_M@ ~�@h����T$X`x ��T$HBK���F��A�q����PPA�
���	������DVC_DB�3@pA �A"��X1`�X3`��S�@�`�0���Uꣳ�h�CAB PP
R�S #��c�B��@���GUBCPU�"��S�P�`R���11)ARŲ�!$HW_CGpl�11� �F&A1Ԡ@8p�$/UNITr�l e ATTRIr@y"��gCYC5B�CA���FLTR_2_�FI������2bP���CHK_��SCmT��F_e'F_o,��"�*FS�Jj"CHA�Q�'91Is�82RSD����1���_Tg�`� i�SEM�NPMf�T&2� 8p&2- �6DI�AGpERAILAiCNTBMw�LO@4�Q��7��PS��梱 � ��PRBS�Z`�`BC4&�	���FUN5s��RIN�PZaߠ�07Dh�#RAH@���`� `C�@�`C�Q�CBL'CURuH�DA�K�!�H�HDAp�aA�H�C�ELD������C��2jA�1�CTIBU�u�8p$CE_R�IA�QJ�AF Pb��>S�`DUT2�01C��};OI0DF_LC�H���k��LMLF�aHRD�YO���RG�@H�Z0��ߠ�@�UMUL�SE�P�'3iB�$J��J����F?AN_ALM�db�WRNeHARDH��ƽ�P��k@2a�N�r�J�_}�AU�J R+4�TO_SBR��~b�Іje 6|?A�cMPINF���{!�d�A�cREGF�NV��ɣZ�D���NFLW%6r$�M�@� ��f� �0l h'uCM4NF�!�ON	 e!e#�(b8*r3F�3 �	 ����q)5�$�$Y�r���u�_��p�*$ �/�EG0@����qAR��i�«�2�3�u�@<�AX�E��ROB��REMD��WR��c�_����SY`��q� ?�S�I�WRI���vE SATհ�ӭ d���Eg!���t8��^a��Bȉ���9�3� OT�O�a���ARY���ǂ�1����FI�E���$LINK��QGTH��Ti_������30���XYZ���!*�'OFF�����%ˀB��,Bl���e���m�FI� ��C@hIû�,B��_J$��F�����S`����3-!$1�w0���R���C��,�DU���3\�P�3TUR`XS�.�Ձ�bXX�� ݗFL�d���pL�0����34���� 1)J�K��M�5�5p%B'��ORQ�6@��fC㘴��0B�O;��D�,������a�OVE��rM�����s 2��s2��r1���0���0�g /�AN=!�2� DQ�q���q�}R�*���6����s��V���E)R��jA	�2E��.�$C��A���0��XE`�2Ӈ�A��AAX�� F��A�N!�SŴ1_� �Q_Ɇ�^ʬ�^ʴ�^�@�0^ʙ�^ʷ�^�1&� ^ƒP[ɒPkɒP{ɒP �ɒP�ɒP�ɒP�ɒP �ɒP�����ɪ �R>�oDEBU=#$8A`Dc�2����
�AB�7�����V� <" 
��i�q��-!��%� �׆��׬��״����1 �י��׷�JT��DR�.m�LAB��ݥ9 �FGRO� ݒ=l� B_�1�u���}���`����ޥ��qa��AND�����qa� �Eq��1��A@�� �NT$`��c�VEL�1��m��1u�0��QP��m�NA[w�(�CN1� ��3줙��e �SERVEc�p+ $@@d@��7!��PO
�� u_�0T ! ������p,  ]$TRQ�b
d(� -DR2,+�"P�0_ . l8"@!�&ERR��"�I� q���~TOQ����L�p]�e���0�G��%��� R}E�@ / ,��/I -��RA� �2. d�&��"  0�p$`&��2tPM��OC�A�8 1  pC�OUNT�� ���SFZN_C;FG2 4B �f�"T�:#��Ӝ�� t$ `�s3 ���M:0�R�q`C@��/�:0�FA1P��?V�X����H�r���� �P:bΣpHELpe4� 5��B_B;AS�cRSR�f @E�S�!QY 1��Y 2|*3|*4|*5*|*6|*7|*8�L!�RO�����NL��q �AB���0Z A�CK��INT_�uUS`�Pta9_P�U�>b%ROU��P�H@�h9#�u`w�9�T�PFWD_KAR���ar RE���PP8��A]@QUE�i&� �	�f�>`QaI`���9#�j3r��f�SE�ME��6��PA�S�TY4SO�0�D�I'1�`���18�rQ_�TM�cMANRQ�XF�END�$�KEYSWITCaHj31:A�4HE	��BEATM�3PE��pLE��1��HU�~3F�42S?DDO/_HOMBPO:a0EF��PRr��*�v�uC�@O�Qo �OOV_Mϒ��Eq�GOCM���7���v:#HK�q5 D�$�g�Uj�2M�p�4�R��FORC�cW;AR���]:#�OM�p 6 @��Ԣ�v`U|�P�p1��V'p�T3�V4��T�Q#O�0L�R7���hUNLOE0h�dEDVa  �9S�@d8 <pAQ�9�l1MSUPG��UaCALC_P�LANcc1��AY�S1�@�9 � 	X`��P �q;a@�թ�w��2��j�M$P��㣒�fyt$��rSC�M�pm�q ���aq���0�tYzZzE!U�Q�b�� T!�Hr��pPvNPX_A�Sf: 0g AD�D��$SIZ�%a$VA��M_ULTIP�"ns��PA�Q; � �$T9op�B���rS��j!C~ �vFRI	F�2S�0�YT�p{NF[DODBUX�`B��u&�!���CMtA�Е����������\Z ��< � ��p�TEg�����$�SGL��T��X�&�{���㰀��STMyTe�ЃPSEG�2���BW���SHO�W؅�1BAN�`TPO���gᣥ�����ѵ7 V�_G�= Y�$PC����O�FB�QP\�SPb�0A&0^�9`VDG�~�>� �cA00�����P���P����P���P��5��6���7��8��9��A ��b`���P��w᧖S`B��F����h���1���v�h�י1�1�1���1�1�1%�1�2�1?�1L�1Y�1�f�2��2��2��2�ʙ2י2�2�2���2�2�2%�2�2�2?�2L�2Y�2�f�3��3��3��3*ʙ3י3�3���T��3�3%�32�U3߹3L�3Y�3f�U4��4��4��4ʙU4י4�4�4��U4�4�4%�42�U4߹4L�4Y�4f�U5��5��5��5ʙU5י5�5�5��U5�5�5%�52�U5߹5L�5Y�5f�U6��6��6��6ʙU6י6��6�6��U6�6(�6%�62�U6߹6L�6Y�6f�U7��7��7��7ʙU7י7��7�7��U7�7(�7%�72�U7߹7L�7Y�7f�zORV�`_UPD���? �c 
�B����@ x �$TOR�1T� � �cOP �, ZQ_7RE^��� J�J�SsC�A���_U�p�YSL}OA"A � �u $�v��w�@���@��bVALUv10�6��F�ID_L�[C:HI5I�R$FILE_X3eu4s$�C�SAV���B hM �E_B�LCK�3�ȁ�D_CPU��p��p�5hz�pY��R3R� C � PaW��� 	�!LAށ�SR�#.!'$RUN�`G@%$D!'$@�@G%e!$e!'%HR0�3$� '$��T2Pa_�LI�RD  �� G_O�2�0P�_EDI�R@�T27SPD�#E�"i�0ȁ�p�Q�DCS�9@G)F � 
$JPC71q�� �S:C;C9$7MDL7$5P>93TC�`@7UF�@?89S� ?8COBu �@Q�"|�L�G�P;�;� 9:;~8`TABUI_�!"L�HGb�%�0FB3�G$�3A�sR�LLB_AVAI�Bp6`�4�!��I $� 7SEL� NẼ�@RG_D N��Ta<G{SC�PJ �1�/AB�PT�R<D_M]`L�K \M f/Q�L_��FMj��PG�i�U9R�6��PS�_�P\� �p�EE�7B�TBC2�eL� ���``�`b$�!FT�P'T�`TDCg�� BPLp�sLNU;WTH��qhT�gtWR�2$�pERVE.S�T;S�Tw��R_ACkP MX -$�Q�`.S �T;S�PU@�`IC�`7LOW�GF1�QR�2g�`��p�S�ERTIA�d^0iP��PEkDEUe�LA7CEMzCC#c��V�BrpTf�edg�aT�CV�l�adgTRQ �l�e�j|�Scu��edcBu�J7_ 4J!���Se@qde�Q2��0���1�PRcuPJKlvVK<�~qcQ~qw�bspJ0��q�sJJ�s;JJ�sAAL�s�p �s�p�v���r5sS�`N1�l�p�k�`5dXAa_́0QCF�B�N `M GROUP ��bh�NPC0s~D�REQUIR�R�� EBU�C�Q�6g0 2Mz��Pd�VQSGUO�@�)/APPR0C7@� �
$� N��CLOD� ǉS^U܉Se
Q��@A�"P �$PM�]P�`�`sR�_MGa!�C���+��0�@�,�BRK*�NOL�D*�SHORTM!O�!m�Z��JWA�SP�tp`�sp`�sp`�s�p`�sp`�A��7��8�sQ!�QTQ� m��R.Q�cQ�PATH�*� �*���X&���P�NT�|@A�"p��� �INF�RUC4`a��C�`KUM��Y
`�)p ��>�Q��cP���p���PAYLOAh�J;2L& R_Am@ꥁL �����+�R_F2LSHR�T/�LO���0���>���ACRL0z�p�y��ޤsRH5b$H�+���FLEX��:#�JVR P��_�._�_�_QJ�US :�_�Vd`0ǀG��_tQd`�_�_lF1G��ũ�o0oBoTofoxo��E�o�o�o�o �o�o�o ����w z3lt����3EWF�^zT!��X�'qju ��uu~�W؁�� �p�u�u�u�u����� 	��(�T ��P5�G�Y�' AT��l�pEL0�_B��js�J�Sz�JEW�'CTR7B`NA���d�HAND_VB�����TUO@h`+�`TSW��=A�A�V� $$M��e G�A@V�Qs�De�oAA ��@�	$�A5�
G�AU�Ad�� 6���G�DU�Dd�PD�G/ -STI�5V�5Ng�DYF ��+�x ����P&�G�&�A�� lw�o�Q�k�P�������ʕӕܕ��"�J�UW 7 �� ���3%�?!ASYIMT��m�T�V�8o�A�t�_SH�~� �����$����Ưد�J񬢐�#39"�.��_VI��`8�>q0V_UNIrS�4��.�Jmu�2��2A� �4X��4�6a�pt��������&E_����������TE��CH~( X ̱l���TOc�PPСVsSvD�US�RU�P������z@�D�A}@_�5�U��P�EyAa��RP�ROG_NA��}$�$LAST����CANs�ISz@XYZ_SPu�DW]R@Ͱ,VSV@�E1QsENc��DCUR�H�����HR_T��YtQ9S�d���O�TNAuP?�Z) ��I�!A�D�� �Q���#�S����3��vP [ � ME�O��R#B�!T�PPT0F@1�a��̰� h1a�%iT0� $�DUMMY1��o$PS_��RF���  1�lfװFL�A*�YP�bc?$GLB_TI �Up�e`ձ��LIF(!�\����g`OW��P��eVOL#qLb �a_2��[d2[`����b�P�cZ`T�C��$BAUD,v��cST��B�2g`�ARITY0sD_[WAItAIyCJ�2�OU6�ZqyyT�LANS�`�{S�SyZc��BUF_�r��fиx�PyyCHK]_�@CES��� +JO`E�aA�x�bUBYT���� �r�.�.� ��aA���M�������Q] �Xʰ����ST����SBR@M21�_@��T$SV_cER�b����CL�`ʐ�A1�O�BpPGL�h0EW(!^ 4 �$a$Uq$�q$W�9�A��@R����ӃU�م_ "��D$�GI��}$ف ���Ӄ�(!` L��.��"}$F�"E�6�NEAR��B�$F}��TQL���& J�@R� a�7�$JOINTxa�)�хMSET(!b  +�Ec�2�^��Se�
H�_�(!c��  ��U�?����LOCK_FOx@� �PBGLV���GL'�TE�@XM����EMP��:�8K��b�$U�؂Fa�2_���q�`<�h �q�^��CE/�|?��� $KARb�}M�STPDRA܀����VECX�����kIUq�av�HE�OTOOL���V��;REǠIS3���6��ACH̐m b&^QONe[d3����IdB�`@$RAI�L_BOXEa�ι�ROB�@D�?�~��HOWWAR0Axa�i`-�ROLMtb ��$�*���T��`����O_FU�!��HTML58QS��  e�MBՀ�(!d��nP�@�(!e����������}p(!f 	t��m�^a��t��VB�PO��AIPE�N���O����q�|�AORDED��m �z�XT`��A)�t`pPP�O�P go D �`OB� ����ǯ�Uc�`��� ��SYS��ADR���pP`U@^  hs ,"��f$A���E��E�VW�VA�Qi � 1�@ق�UPR�B��$EDI�Ad�V/SHWRU�z���cIS�Uq�pND�Px7���G�HEAD�!h @���!i�KEUq�O`CP)P��JMP���L�UoPRACEV�Tj���IL�5S��C��NE���TICK!M�KQс��HNr�Gk @���HWC��qPHVF��`STYeB+�LO�a����[��C�l3�
�@�F%$�A��D=��S�!�$�1�p a�e�q�eP�v HVSQU��#LyO�b_1TERC`�!�PS?�m  5���R�m@3���ܡ�1O`	c IZ�d�A�eha�qtb}�hA}p9P~r��_DO�B��X�pSSQ�SAXI��q��v�bS�U�@TxL���REQ_ܠ���ET���`�CY%���FY'��Af\!e\d9x�P Ђ{SR$$nl-� w �����c
�u!V
Qh(�A���dC`�A��	�Y��D��p�E"�	CC�C��/�/��/	4��SSC�` oo h5�DSm�̟Q[`SP�@�AT�� 
R��L��XbA7DDR�s$Hp� �IF�Ch�_2CH����pO����- �TuUk�Ir p£CUCpсV��I��Rq�4���c��
�K�
�RV*���Pr \z�D����|,K� P�"CN��*C�����!�TXSCR�EE��s�Pp@�ICNA˃<�4�D"�8����`t Tᫀ �b����O Y6���º�U4h�RR��������R1�T��UE��u ��j �qz`Ś��RSML��U����V�1tPS_��6\��1�9G\���C��2@4� 2��0Ov�R��&F�AMTN_FL*�`Q��W���/BBL_/�WB`�P�w ����BO ��BLE"�Cg�R"�DoRIGHtRD���!CKGRB`�ET����G�AWIDTH�s���RB��a�r��UI��EYհRx� d�ʰ�����`y�BACK��tb>U����PFO��QWL[AB�?(�PI��$URm�~Pр�P�PHy1 y o8 $�PT_��,"�R�PRUp�s5��da�1hq%!t�zV�$ȇ�pU�@�SR ����LUM�S�� ER�VJ��SP��T{ 7� " GE�Rh�� �¯�LPAeE��)^g�lh�lhT�ki5ik6ik7ik pP`�Z�x����$u�1��p�Q z�QUSRل| �<z��PU2�a#2�F�OO 2�PRI*mx9�[�@pTRIPK�m�UNDO��})���Yp��y���Pi����p ~��Rp�qG ��T0���-!�rOS2��vAR��2�s�CA�@����r`�1i�UIaCA����3Ib_�s�OFFA�D@���Ob�r�5�L�t��GU��Ps���������+QSUB`� }��E_EXE���VeуsWO� e�#��w��WAl��p΁fP
 V_CDB���!pT�p�O�V░���3OR�/�5�RAU@6�T�K���__����s |j �OWNj�>34$SRC�0`����DA���_MPFqI����ESP��T�$0��c��g��8n�z�E!� `%�ۂr34J���COP��$`��p_���/�+�6���CT�Cہ铸ہ���DCS��P�4�COMp�@�;��O`�=���K�^�/��VT�q'���Y٤Z��2���@p�w#SB����2�\0˰�_��M��%!]�DI�C#��AY�3G�P�EE�@T�QS�VR�1���eQL�� a� �P�D ��f�z��f� > ���6����A�t��b# �L2SHA�DOW��#ʱ_U�NSCAd�׳OW�D�˰DGDE#L�EGAC)�q'��VC\ C���� v����だm�R F07���7d`C2`7�/DRIVo���Ϡ�C�A]�(�` ���MY_UBY�d?Ĳ� �s��1��$0���𣢌�_ఆ���L��B�M�A$�DEY�	�EXp@C�/�MUb��X��,��0US����;p_R"1�0p#�2�GPACIN*���RG��c�y��:�y��sy�C/�RE�R"!�qsB�y�D@�� L !�G�P��"��y@�R�pD@� &P�Px1Q��	.����RE��SWq�_A$r�u@+�{�Oq�AQA/�3�hEZ�U��Ώ� n��HK
���PJ��_/�Q0{�EAN��ۀ2�x2�Tp�MRCVCAw� �:`ORG���Q�dR	��L�����REFoG�����!�+` 	�p��������<���q�_����r���� S�`C��Ú��q�@D� ��0�!��#q�š�OU����?�� ��Վ2�`J@0� 1�*p�����0 UL�@͋�CO�0)��� NT�[i�Z �Qf�af% L飏���Q��a�V�IAچ� �ÀHyD7 6P$JO�`�oB�$Z_U�Po��2Z_LOW���$�QiBn��1$EP�s�y�� 1!f �� 1¦4ߏ 5�PA��A �CACH&�LO�w�В��1B���Cn�I#F�^��Tm����$H	O2�32{��Uÿ2O�@���Ro��=a���ƐVP��X@A"_'SIZ&�K$Z$�F(��G'���CMPk*F�AIo�G��A9D�)/�MRE���"�P'GP�0е�9�A�SYNBUFǧR�TD�%�$P!�COL�E_2D_4�5WH�sw�~�UӍQO���%ECCU��VE�M��v]2�VIRAC�!5�#�2�!_>��*&�pWp��AG	9R��XYZ@�3�W@���8��4+Qz0T"��IM�16�2P�GRABB�q��;��LERD�C ;�Fc_D��F�f50MHH�PE�R[����JRLAS�@��[w_GEb� �H���~23�ET����"���b��I�D�ҙ6m�?BG_LEVnQ{��PK|Л6\q��GI�@N\P4���P�$�!g�dr�S� �INRT\�Lʁc�Ų���#a��c"!D�qDE����Xа�X��E ��2��d��pAzZ���d�c����D4qȾ�2pT��Un&�� $�ITPr�9p[Q��ՓV�VS9F$�d�  fp/�Lf�UR��QaMZus�dr��ADJ`�C�� ZDVf� D�XAL� � 4 �PERIKB$MoSG_Q3$Q!�o%z���p'���dr:g�qQ� �X�VR\t��B�pT_�\��Rm�ZABCB"����Sr���
��aACTVS' � � $|u<�0�cCTIV�Q!�IOu¥s&D�ITl�x�DVϐ
xѤP���!���pP	S���� �#��!���q!LSTD�!� l �_ST�1��wrq�CHx�� L -�@��u�Ɛ*���P GNA#�C�!q�_FUN�� m�7ZIPu��HR�S$L���XZ��F"��`bƀ�rX�فn��LNK��
Ł��0#�� $x !��ބCMCMk�EC8�C"����P{q? $J8�2�D6!>�O�H�i�T�i�`2�����M���UX�1݅UXE1Ѡ��1C� ��Y���������˗7��FTFG>������{�Z��� �k���l��YD'@ �� 8n�R� U�ӱ$HEIGH�d�:h?(! 'v�|6���� � Gd��qp$B% � E���SHIF��hRVBn�F�`�HpC�  3�(�8H`O�ѡ�Cd��+%D	�"�CE�p�V�1vp��PHER>s� � ,! M��c�u��$POW�ERFL �P|�����|�p�RG�` � �������A�  ���?�p���pd��N�Sb ����?�  B�z|� l�  <@1�|�Z�|�%����˃����ŵ�� 2yӷ�� 	H���l&���>�着A |��t$���*��/�� **:���p�ϥ���2��������������|�����5��� ����%ߟ�I�[߉� ߑ����������� w�!�3�a�W�i���� ��������O����9� /�A���e�w������� '�����= O}s����� ��k'UK] ������C/� �-/#/5/�/Y/k/�/ �/�/?�/�/?�/? �?1?C?q?g?y?�?�? �?�?�?�?_O	OOIOx?OQO�� 	 �O �O�O_�E��3_���O�`_�O�_�_÷PREOF Ӻ�p�p�
��IORITY! 4�|����p����p�SPL`z����WUT8�VqÈ�ODU~������_?�OG�Gx��R��,fHI�BqOy�|kTOE�NT 1��yP(!AF_b�`�o~�g!tcp�o>}!ud�o)~?!icm��0bXY̳�k �|�)� �����p����u�� ����N�5�r�Y��������̏�����*/c̳ӹ���E�W�^|�>���F��!/��4���|��,�7��A��,  ��P����%�|�'���Z��h�z������|��ENHAN�CE 	#�7�A�9�d�����  ��,f�T
�_�S�����PORTe�rb�@�U��_CARTREP�Pr|br�SKSTAg�kS�LGS�`�k�����@Unothing����π�Ϳ>�P�b�To��T?EMP ?is���E/�_a_seibanm_��i_�� ���0��T�?�x�c� �߇ߙ��߽������ �>�)�N�t�_��� �����������:� %�^�I���m������� ���� ��$H3 lWi����� ��D/hS��w���uϪ�VOERSI�P=g � disab�le��SAVE� ?j	26�70H705��k/!�m//*�/C 	�(%b�O�+�/�Se?6?H?Z?l?z:A%<�/�?4�*'_j`W 1�kX �0�ubuE�?OqG�PUR�GE��Bp`�ncqWAF<@�a�TӒ*fW�`�]Daa�WRUP_�DELAY �z�f�B_HOT �%?e'b��OnER_NORMAL�H�Gb�O%_�GSEMI�_*_i_�QQSKI%P�3.��3x��_ ��_�_�_�]?eo+g oKo]ooo5o�o�o�o �o�o�o�o�o5G Yi�}��� ����1�C�U�� y�g���������я�����-�?�7%�$RACFG �[�ќ�3�]�_PA�RAM�Q3y��S; @И@`�G�4W2C۠��2���CbFB�B]�BT�IF���J]�CVT�MOU������]�DCR�3�Y� ��UBh��B�@���4>V�h9�X;�]�>�>�v��_|����;e�m����KZ;�=g;�4�<<���pf@����� � 5�G�Y�k�}��������ſ׿���xURDI�O_TYPE  ��V�5��EDPR�OT_a�&Y>��4BHbCEސ�SǆQ2c� ��B�ꐪϸ���� �����&�ݹ�W�V_ ~�o����߱����� ����A�O�m�r��� 9����������� ���=�_�d����� ������������' I�Nm���� �����#EJ i+k���� ��//4/F//g/ /�/y/�/�/�/�/�/ 	?+/0?O/?c?Q?�? u?�?�?�?�?�??;?�,O��S�INT 2��I���l�G;�� jO|K��鯤O�f�0 �O�K�?�O�? ___N_<_r_X_�_ �_�_�_�_�_�_�_&o oJo8ono�ofo�o�o �o�o�o�o�o"F 4j|b����������B�O�E�FPOS1 1~"�  xO ��o×O����ݏ鈃� ��Ϗ0��T��x�� ��7���ҟm������ ��>�P����7����� ��W��{�����:� կ^����������S� e��� ��$Ͽ�H�� l��iϢ�=���a��� ��� ߻����h�S� ��'߰�K���o���
� ��.���R���v��#� 5�o���������� <���9�r����1��� U�����������8# \����?�� u��"�FX� ?���_�� /�	/B/�f//�/ %/�/�/[/m/�/?�/ ,?�/P?�/t??q?�? E?�?i?�?�?O(O�? �?OpO[O�O/O�OSO �OwO�O_�O6_�OZ_ �O~_�_+_=_w_�_�_ �_�_ o�_Do�_Aozo<cf�2 1r�o .oho�o�o
o.�o R�oO�#�G� k�����N�9� r����1���U����� �����8�ӏ\���	� �U�����ڟu����� "����X��|���� ;�į_�q������	� B�ݯf����%����� [���ϣ�,�ǿٿ �%φ�qϪ�E���i� �ύ���(���L���p� ߔ�/�A�Sߍ����� ��6���Z���W�� +��O���s����� ����V�A�z����9� ��]���������@ ��d��#]�� �}�*�'` ���C�gy ��&//J/�n/	/ �/-/�/�/c/�/�/? �/4?�/�/�/-?�?y? �?M?�?q?�?�?�?0O �?TO�?xOO�O�o�d3 1�oIO[O�O _�O7_=O[_�O__ |_�_P_�_t_�_�_!o �_�_�_o{ofo�o:o �o^o�o�o�o�oA �oe �$6H� ����+��O�� L��� ���D�͏h�� �������K�6�o�
� ��.���R���퟈�� ��5�ПY�����R� ����ׯr�������� �U��y����8��� \�n�������?�ڿ c�����"τϽ�X��� |�ߠ�)�������"� ��nߧ�B���f��ߊ� ��%���I���m��� ,�>�P��������� 3���W���T���(��� L���p����������� S>w�6�Z ����=�a � Z���z /�'/�$/]/��/�/�/@/�/�O�D4 1�Ov/�/�/@?+? d?j/�?#?�?G?�?�? }?O�?*O�?NO�?�? OGO�O�O�OgO�O�O _�O_J_�On_	_�_ -_�_Q_c_u_�_o�_ 4o�_Xo�_|ooyo�o Mo�oqo�o�o�o�o �oxc�7�[ ����>��b� ���!�3�E����ˏ ���(�ÏL��I��� ���A�ʟe���� ���H�3�l����+� ��O���ꯅ����2� ͯV����O����� Կo�����Ϸ��R� �v�Ϛ�5Ͼ�Y�k� }Ϸ���<���`��� ��߁ߺ�U���y�� ��&���������k� ��?���c������"� ��F���j����)�;� M���������0�� T��Q�%�I��m��/�$5 1 �/���mX�� �P�t�/�3/ �W/�{//(/:/t/ �/�/�/�/?�/A?�/ >?w??�?6?�?Z?�? ~?�?�?�?=O(OaO�? �O O�ODO�O�OzO_ �O'_�OK_�O�O
_D_ �_�_�_d_�_�_o�_ oGo�_koo�o*o�o No`oro�o�o1�o U�oyv�J� n������� u�`���4���X��|� ޏ���;�֏_����� �0�B�|�ݟȟ��� %���I��F����� >�ǯb�믆������ E�0�i����(���L� ��翂�Ϧ�/�ʿS� � ��LϭϘ���l� �ϐ�ߴ��O���s� ߗ�2߻�V�h�zߴ� � �9���]��߁�� ~��R���v����#�<	6 1&�� �������������}� ��<��`��� �CUg�� &�J�n	k� ?�c��/�� �	/j/U/�/)/�/M/ �/q/�/?�/0?�/T? �/x??%?7?q?�?�? �?�?O�?>O�?;OtO O�O3O�OWO�O{O�O �O�O:_%_^_�O�__ �_A_�_�_w_ o�_$o �_Ho�_�_oAo�o�o �oao�o�o�oD �oh�'�K] o�
��.��R�� v��s���G�Џk�� �����ŏ׏�r�]� ��1���U�ޟy�۟� ��8�ӟ\������-� ?�y�گů����"��� F��C�|����;�Ŀ _�迃������B�-� f�ϊ�%Ϯ�Iϫ��� �ߣ�,���P�6�H�7 1S����I� �߲�������3��� 0�i���(��L��� p�����/��S��� w����6�����l��� ����=������6 ���V�z�  9�]��� @Rd���#/� G/�k//h/�/</�/ `/�/�/?�/�/�/? g?R?�?&?�?J?�?n? �?	O�?-O�?QO�?uO O"O4OnO�O�O�O�O _�O;_�O8_q__�_ 0_�_T_�_x_�_�_�_ 7o"o[o�_oo�o>o �o�oto�o�o!�oE �o�o>���^ �����A��e�  ���$���H�Z�l��� ��+�ƏO��s�� p���D�͟h�񟌟� ��ԟ�o�Z���.� ��R�ۯv�د���5��ЯY���}�c�u�8 1��*�<�v���߿ ��<�׿`���]ϖ� 1Ϻ�U���y�ߝϯ� ����\�G߀�ߤ�?� ��c����ߙ�"��F� ��j���)�c���� ������0���-�f� ���%���I���m�� ����,P��t �3��i�� �:���3� �S�w /��6/ �Z/�~//�/=/O/ a/�/�/�/ ?�/D?�/ h??e?�?9?�?]?�? �?
O�?�?�?OdOOO �O#O�OGO�OkO�O_ �O*_�ON_�Or___ 1_k_�_�_�_�_o�_ 8o�_5ono	o�o-o�o Qo�ouo�o�o�o4 X�o|�;�� q����B��� �;�������[��� ����>�ُb������!�������MASKW 1 ��������ΗXNO  �ݟ���MOTE � ���S�_CFG' !Z���N������PL_RANG�V�N������OWE/R "��Ϡ���SM_DRYPRoG %���%W���եTART �#Ǯ�UME_P�RO���q���_E�XEC_ENB � ����GSPD�J�������TD�B����RMп��I�A_OPTION��������N�GVERS���`�řI_AIoRPUR�� R��+���ÛMT_֐T� X���ΐOBOT_ISOLC�����������NA�ME8��H�ĚOB?_CATEG�ϣ�,��S�[�.�OR�D_NUM ?�Ǩ��H705  N��ߨ����ΐPC_TIMoEOUT�� xΐoS232s�1$���� LTE�ACH PEND�AN��o���)���V�T�Mai�ntenance_ ConsN�&��M�"B�P�No Use6�r�8���������̒��NPO�$��Ҏ�"���C�H_LM�Q���	�a�,�!UD1�:��.�RՐVAI�Lw��粥*�S�R  t� ����5�R_INTVAL���� ����V_DATA_?GRP 2'���_� D��P�� �����	���� ��B0RT f������/ �/>/,/b/P/�/t/ �/�/�/�/�/?�/(? ?L?:?p?^?�?�?�? �?�?�?�?O O"O$O 6OlOZO�O~O�O�O�O �O�O_�O2_ _V_D_ z_h_�_�_�_�_�_�_ �_o
o@o.oPovodo��o��$SAF_DO_PULSW��[�S���i�SCANd�������SCà�(6�7}���S�S�
������q�q�
qN� �L^p ���5��� �X�$��+��r2M�qqdY�P�`�rJ�	t/� @��@������ʋ|��� r �ք��_ @N�T ��'�9�K�X�?T D��X��� ������ɟ۟���� #�5�G�Y�k�}�����x��䅎������Ǧ  "�;G�oR� ���p�"�
�u��D�i���q$q�  � ���uq%�\� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z����珈������ ������g�;�D�V� h�z���������������(�Ӣ0�r�i�y� ��$�7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/?r�+?=?O?a? s?�?�?�?�?�?8��? OO'O9OKO]OoO�O ��$�r�O�O�O�O 	__-_?_Q_c_u_�_ �Y�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4@FXj|�c�路 g�������0� B�T�f�x���������ҏ������:�.Ҧ��y�3�	��	123456�78��h!B!�� \��p0����Ο�� ���(�:�@��c� u���������ϯ�� ��)�;�M�_�q��� ��R���ɿۿ���� #�5�G�Y�k�}Ϗϡ� �����ϖ�����1� C�U�g�yߋߝ߯��� ������	��-���Q� c�u��������� ����)�;�M�_�q� ��B���������� %7I[m� �������! 3EWi{��� ����////� S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?D/�?�?�?�?�? OO'O9OKO]OoO�O@�O�O�O�O�O*��� �O	_�E�?5_G_Y_�yCz  A��z_   ��x2�r� }��)�
�W�  	�*�2�O�_�_ o$o"l�#\��_ho zo�o�o�o�o�o�o�o 
.@Rdv� ���Mo���� *�<�N�`�r������� ��̏ޏ����&�8��J��X #P$P�Q�R<�u� k��Q  ������S�P����Q�Qt  ЌPÙ۟�P(� `�,b����]�PFl��$SCR_GRP� 1*7+�74� � ��,a �U	 v��~������d���%����ɯ���h]���P�D1� D�7n��3��Fl
C�RX-10iA/�L 234567W890�Pd� r���Pd�L ��,aC
1o��������[ ¶~�+fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@�R�d�t�?��H�~����m��ϴ����������,a��1���U��[�G�imXhuP,[���뾥B�  CBƠߞҷԚ�A�P���  @1`�՚�@9����� ?����H����ښ�F@ F�`A�I�@�m� X��|��������� ��������:�%�7�I�[�B�i������ ����������-Q <u`��En�ٯ���W�P�"+f�@_�5��1`b���x����ͣ�O��,dA������$�Fa�,a �# !"/4/E-!Z(f/�x/G/ (�P�!( � �/�/�/��/�/?�#9b����S7س��M�ECLVL  �,a��ݲ�Q�@f1L_DEFA�ULTn4b1��1`�3HOT�STR�=��2MI�POWERFm0�pU�5�4WFDO�6 �5L�ERV?ENT 1+u1u1��3 L!DU�M_EIP#?5H��j!AF_IN�E�0SO,d!FT$)O�NIO�O!���O� ��O�O!RPC_MAIN�O��H��O>_SVIS�_�I�-_�_!O�PCUf�_�W�y_�_!TP�PP�U�_<Id�_"o!
�PMON_PROXY#o?Feono�R�<o8Mf]o�o!R?DM_SRV�o<I9g�o!R��"�=Hh�oR!
PM�o9LiA�!R�LSYNC��y�8��!ROS�(O��4�6�!
�CE�PMTCOMd7�?Fk%���!	K�OCONS��>Glq��Ώ!K�WASR�C�o?Fm���!NK�USB�=Hn	�>f�!STM�0��;JoU����O֟�c�����CICE_KL� ?%K (%�SVCPRG1���G�1�2G�L�6�3�o�t�6�4����6�5���į6�6��6�7@��6���W�R�9_�d�3���6�9��� 6�a�ܿ6����6��� ,�6�ٯT�6��|�6� )���6�Q���6�y��� ^����^�ʿD�^�� l�^�ϔ�^�Bϼ�^� j���^����^���4� ^���\�^�
߄2� ��6��/����V� �<�'�`�K���o��� ����������& J5nY���� ����4F1 jU�y���� �/�0//T/?/x/ c/�/�/�/�/�/�/�/ ??>?)?P?t?_?�?�
�_DEV ~I�MC:�8�4���4GRP� 2/E�0+�b�x 	� 
 ,@�0�?OD!OKODdOvO]O�O �O�O�O�O�O�O_�O _N_5_r_Y_�_�_/C
E�0�_�_�_o �_'ooKo]oDo�oho �o�o�o�o�o�o�o�o�5Y�_D	�0 i@������ � �=�$�a�s�Z��� ~��������؏�lD6OS�D�~�1O������ן
���� ���U�<�y�`��� ����ӯ*��V ��	A �_:�ů^�E�����{� ����ܿÿտ���6� �Z�l�Sϐ��	A�q ����%��Ϲ����υ� �'߅�v�]ߚ߁߾� �߷������*�5�N� ��r��������� �����&�8��\�C� ��g�y����������� g�4-jQ� u����� B)fx_�� ��)��/,// P/7/t/[/m/�/�/�/ �/�/?�/(??L?^?�E?�?�7d �[~�
�6 s�p�A;*=� 6�?�=���D��>����g��:�0��ī����|@�-�@��5_�eA5��-�=BG+h��&���6)AB��m�����`x��=�?7O%?TELEOP8OcN�[~y��5�o��ʾTF������������|��ҝ�����E�1�E�@�*�A`�~��n�!��$��A���M�Y<�T�������C=�J����Gc��McO��IJO/_�[~���6r _�1<��׻��y;�?�	A`�ʛ1bP���N	V�A��&@в@����@)E�]�1������0ד�� x���Q��U?�Q��O`�__ _oDU�NU�9��6>���E�bQ�2]��j_ ��r�AS�AT��@��@G$���_ ��yC�� �Pr}��Q� ?2i?�R�_�o��_�_�oDU�K�5���l�������S���`
�� 3>v�ĚM�@�@�V��@�%@������q���]V��N��N�!C(�uµ��� �®����ow�o�o�DU�b��5?��T��@O�P�%��*�-��Ƒ��N�PA�����
Q@���q�A��M��{�B&�b�r'C9rt��1��^Ѻ@fK�������p�m�5>���@�����͙~�E��A������c�N'pA(��AC8AD�����A�y��Nd�A��R���ֺ�����s��`_�^`��\�n�S�BW�c�v�"��?/����H?��4@�� �+79���$ΏA8	A�Alܾc`�fߩ@�c+�Ne?�6A�z2��L�Q� f��t���`�D��2��D�)�DT�m��6M��W�1�������F0�<?
u���8�NW`�@�^}A1Nu�@X�ƿP��A%��N�j!���g(�E�u�B��y�!F�`G�/������:�p��6
������\��w�������kuf@��In_�PI3��@K�@�"����P��섆��NuN�A��Q�¸!C=������º��`��ٯ�п;�t2�0��Bq̾���?P�������lG-���~�u�AR���@&G Az����:�AX����NzQBA������V�����uC����׿�����ϒ����6 *���f��?#� ;����>b8�34��=+F':�V��?��r@��/�>�@?[����n�MA��q�����
]�@����3�xA?8m^�C߂ϔ�y߆<���5�1*a�:�����2��  ����?�!����OLp��A���� ���!�`����`�V�h�M�Ż��5����]�_�?��A������+@�t���M?�<n@���@�o���[��A�
ޭ��@�C��/����=ؕ�{Ӎ�S�(� :��BU�I�IN�<�r�``���������%�'� ��ho��(L:p ^��������� �$H6l�� �\����� / /D/�k/�4/�/�/ �/�/�/�/�/?^/C? �/?v?d?�?�?�?�? �?$?	OO�?�?�?<O rO`O�O�O�O�?�O O �O__$_&_8_n_\_ �_�O�_�O�_�_�_o �_ o"o4ojo�_�o�_ Zo�o�o�o�o�o ro�oi�oB��� ����J/�n� b��r����������� "��F�Џ:�(�^�L� n���������ߟ��� � �6�$�Z�H�j��� ҟ�������د��� 2� �V���}���F�h� B����Կ
���.�p� Uϔ�ψ�vϘϚϬ� �����H�-�l���`� N߄�rߔߖߨ��� � �D���8�&�\�J�� n���������� ��4�"�X�F�|���� ��l���h�����0 T��{��D�� ����,nS ��t���� �/F+/j�^/L/ �/p/�/�/�//�/? �/�/�/$?Z?H?~?l? �?�/�??�?�?�?O O OVODOzO�?�O�? jO�O�O�O�O_
__ R_�Oy_�OB_�_�_�_ �_�_�_oZ_�_Qo�_ *o�oro�o�o�o�o�o 2oVo�oJ�oZ� n���
�.� "��F�4�V�|�j��� �Ǐ�������� B�0�R�x�����ޏh� ҟ�������>��� e�w�.�P�*���ί�� ���X�=�|��p� ^�������ʿ���0� �T�޿H�6�l�Z�|� ~ϐ������,϶� � �D�2�h�V�x����� ��ߞ������
�@� .�d�ߋ���T��P� ��������<�~�c� ��,������������� ��V�;z�n\ ������. R�F4jX�| �������/ B/0/f/T/�/��/� z/�/�/�/�/?>?,? b?�/�?�/R?�?�?�? �?�?�?O:O|?aO�? *O�O�O�O�O�O�O�O BOhO9_xO_l_Z_�_ ~_�_�_�__�_>_�_ 2o�_BohoVo�ozo�o �_�oo�o
�o. >dR��o��ox ����*��:�`� ����P�����ޏ̏ ���&�h�M�_��8� �������ڟȟ��@� %�d��X�F�h�j�|� ����֯���<�Ư0� �T�B�d�f�x���� տ������,��P� >�`϶�ܿ��쿆��� �����(��Lߎ�s� ��<ߦ�8߶����� � ��$�f�K���~�l� ����������>�#� b���V�D�z�h����� �������:���. R@vd����� ����*N< r���b��� ��&//J/�q/� :/�/�/�/�/�/�/�/ "?d/I?�/?|?j?�? �?�?�?�?*?P?!O`? �?TOBOxOfO�O�O�O O�O&O�O_�O*_P_ >_t_b_�_�O�_�O�_ �_�_oo&oLo:opo �_�o�_`o�o�o�o�o  "H�oo�o8 �������P 5�G�� ��h����� ���(��L�֏@� .�P�R�d������� � �$�����<�*�L� N�`���؟������� ޯ��8�&�H���į ��ԯn�ȿ���ڿ� ��4�v�[Ϛ�$ώ� � ���ϲ������N�3� r���f�Tߊ�xߚ��� ����&��J���>�,� b�P��t������� "����:�(�^�L� �������r���n���  6$Z����� J������ 2tY�"�z� ����
/L1/p �d/R/�/v/�/�/�/ /8/	?H/�/<?*?`? N?�?r?�?�/�??�? O�?O8O&O\OJO�O �?�O�?pO�O�O�O�O _4_"_X_�O_�OH_ �_�_�_�_�_�_
o0o�r_Wo�U�P�$S�ERV_MAILW  �U�`��Q~vdOUTPUT�h_�P@vd�RV 20f  �` (a\o�ovd�SAVE�l�iTO�P10 21�i� d 6 s��P
6r _�Pz:p�a6 *�a 2ohz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ���0&�8�iuYP�c�FZN_CFG ;2e�c�T��a�e|�GRP 2�3��q ,B �  AƠ�QD;�� BǠ�  B�4�SRB21��fHELL�4ev�`�o��/�>�%RSR>�?�Q� ��u�����ҿ����� �,��P�;�t�_Ϙ�������  ��¼����Ϸͻ�b�P�&�'�ސW
��2�Pd��g���HK 15�� ,ߡ߫ߥ������� ��@�;�M�_�������������OMM 6��?���FTOV_ENB��d�au�OW_R�EG_UI_��bIMIOFWDL*��7.�ɥ��WAIT�\�`ٞ����`����d��TIM�������VA�`����_�UNIT[�*yL]Cy�TRY��u-v`ME�8���a�w֑d ��9� ������<���X�Pڠ6p`?�  ��o+=�`VL��l�fMON_AL�IAS ?e.��`heGo���� ��/)/;/M/�q/ �/�/�/�/d/�/�/? ?%?�/I?[?m??�? <?�?�?�?�?�?�?!O 3OEOWOO{O�O�O�O �OnO�O�O__/_�O S_e_w_�_�_F_�_�_ �_�_�_o+o=oOoao o�o�o�o�o�oxo�o '9�o]o� �>������ #�5�G�Y�k������ ��ŏ׏������1� C��g�y�����H��� ӟ���	���-�?�Q� c�u� �������ϯ� ����)�;��L�q� ������R�˿ݿ�� Ͼ�7�I�[�m��*� �ϵ������ϖ��!� 3�E���i�{ߍߟ߱� \�����������A� S�e�w��4����� ������+�=�O��� s���������f����� '��K]o� �>����� #5GY}�����l�$SMO�N_DEFPRO�G &����� &�*SYSTEM*����RECAL�L ?}� (� �}8copy� frs:ord�erfil.da�t virt:\�tmpback\�=>192.16�8.56.1:15400/�/�/�-�}/K"mdb:*.*`/r/{/??0?6�$3xK$:\�/U0��/0�/�?�?�?� 4K5aS?e?�%�?O#O5O I/[/�/?�O�O �O�/bO�/}O_ _2_ E?�?�?{?�_�_�_�? T_f_�?
oo.oAOSO �OwO�o�o�o�O�Olo �O*=_O_�_s_ ����_�_^�_� �&�9oKo]o���� �����od��o��"� 4�G��}������ �V�h����0�C� U�ޏy���������ӏ n�����,�?�Q�� u���������ϟ`�����(ϻ�tpdisc 0�������ϝϯ�B�conn 1k�e�w��� ,�?�Q�گu��ߘߪ� ��ϯj����(�;� M��q�7��ﹿ˿ \��ρ��$�6�I�[� ����������b��� }� 2E�����{� �����Tf��
 .A�S���w��� �����l��//*/ =O�s�/�/�/� �^/��/?&?9K ]�/?�?�?�?�d? �?O"O4OG/�/�? }/�O�O�O�/VOhO�/ __0_C?U?�?y?�_ �_�_�?�?n_�?oo�,o>W�$SNPX�_ASG 2:����Vao�  b%�7o�~o  ?�GfPA�RAM ;Ve�`a �	lkP�>TDP>X�d�� ��I`OFT�_KB_CFG � CS\eFcOPI�N_SIM  
Vk�b+=OYs�I`RVNORDY?_DO  �eu�krQSTP_D�SB~�b�>kS�R <Vi �� & TELE�O�e�{v>TW`I`T�OP_ON_ER�RxGb�PTN �VeP���D:�RING_P�RM'��rVCNT?_GP 2=Ve�ac`x 	���DP`��я����BgVD��RP 1>�i�` �Vq؏0�B�T�f�x� ��������ҟ���� �,�>�e�b�t����� ����ί���+�(� :�L�^�p��������� ʿ�� ��$�6�H� Z�l�~ϐϷϴ����� ����� �2�D�V�}� zߌߞ߰��������� 
��C�@�R�d�v�� ��������	��� *�<�N�`�r������� ��������&8 J\n����� ���"4[X j|������ �!//0/B/T/f/x/ �/�/�/�/�/�/�/? ?,?>?P?b?t?�?�?��?�?�?�?�?O�P�RG_COUNT��f�P�)IENB�e�+EMUC�dbO_U�PD 1?�{T  
ODR�O�O�O �O�O__A_<_N_`_ �_�_�_�_�_�_�_�_ oo&o8oao\ono�o �o�o�o�o�o�o�o 94FX�|�� �������0� Y�T�f�x��������� �����1�,�>�P� y�t���������Ο�� 	���(�Q�L�^�p� ���������ܯ� � )�$�6�H�q�l�~��� ����ƿؿ���� ��I�D�V�"L_INF�O 1@�E9�@��	 yϽ��������>�~?�zN>G�q<����� A��Y���[��2�#�@"�?Nl,������` ?@ <�@��o� C���B���C��_��0C+�r�|�2��p����-@YSDEBU)G:@�@�o�d�I��SP_PASS:E�B?��LOG �A���A  ro�i�v�  �A�o�UD1:\x��}���_MPC�ݐ�Ek�}�A&�� ��AK�SAV B���IA���*�i��1�SVB�TEM_TIME 1C����@ 0  m�n�.i�ԝ��*���MEMBK  �EA��������X|�@� Z�i��������ȼ�h�9
�� ��@�`r���〮���� �@Rdv�����
Le�// (/:/L/^/p/�/�/�/ �/�/�/�/ ??$?6?H?Z?��SKV�[�EA`j��?�?�?���@�x]2���?i�  0Po�^
:O. @R�O�O�O}N���ǘ ��OBDp��O_'_9_-L2�Y_�_�_�_�_�_o�U�_�_�o'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk�_?T1SVGUNwSPD�� '�����p2MODE_?LIM D���2�t2�p�qE�݉u�ABUI_DCS' H}5���0�G �0��D��|-�X�>�ލ�*���� 
��e��i���r�i������uEDI�T I��xSC_RN J���rS�G K�.�(���0߅SK_OPT�ION��^����_�DI��ENB  �/����BC2_�GRP 2L��0�MPC�ʓ�|/BCCF/�N����c ����`� >�W�B�g���x����� կ��������S� >�w�b���������Ͽ �����=�(�a�L� �ϗ�Ň�϶������� v��
�/�U�@�yߧ� ��`�iМ��߰����� 
���.��>�@�R�� v����������� *��N�<�r�`����� ����������̀ 4FX��|j�� �����B 0fTvx��� ��/�,//</b/ P/�/t/�/�/�/�/�/ �/�/(??L?d?v? �?�?�?6?�?�?�?O  O6OHOZO(O~OlO�O �O�O�O�O�O�O __ D_2_h_V_�_z_�_�_ �_�_�_
o�_.oo>o @oRo�ovo�ob?�o�o �o�o<*Lr `������� �&��6�8�J���n� ����ȏ���ڏ��"� �F�4�j�X���|��� �����֟��o$�6� T�f�x���������ү �������>�,�b� P���t��������ο ��(��L�:�\ς� pϦϔ��ϸ�������  ��H�6�l�"��ߖ� ������V������2�  �V�h�z�H����� ����������
�@�.� d�R���v��������� ����*N<^ `r������� &8�\Jl� �������"/ /F/4/V/X/j/�/�/ �/�/�/�/?�/?B? 0?f?T?�?x?�?�?�? �?�?O�?,O�DOVO tO�O�OO�O�O�O�O��O_ V4P�$TB�CSG_GRP �2O U��  �4Q 
 ?�  __q_[_ �__�_�_�_�_�_o�%k8R?SQF\dאHTa?4Q	 �HA���#e>�w��>$a�\#e?AT��A WR�o��hdjma�G�?L�fg�bp�o�n�ff�hf��ͼb4P|j���o*}@��Rhf�?ff>�33pa#eB<qB�o+=xrRp�qUy�rt~��H`�y rIpTv�pBȺ t~	xf	x(�;��� f���N�`���ˏڋ�����	V3.0�0WR	crxlڃ	*��3R~td��HH��� \��.�]�  cC�.�����8QJ2?SR�F]����CFG [T UPQ SPVܚ��r�ܟ1��1�W�e�	P e���v�����ӯ���� ����Q�<�u�`� ��������Ϳ�޿� �;�&�_�Jσ�nπ� �Ϥ�������WRq@ �0�B���u�`߅߫� ���ߺ������)�;� M��q�\������ 4Q _���O ���J� 8�n�\����������� ������4"XF hj|����� �.TBxf ��nO����/ />/,/b/P/�/t/�/ �/�/�/�/�/�/?:? (?^?p?�?�?N?�?�? �?�?�?�? O6O$OZO HO~OlO�O�O�O�O�O �O�O __D_2_T_V_ h_�_�_�_�_�_�_
o �_o@o�Xojo|o&o �o�o�o�o�o�o* N`r�B�� �����&��6� \�J���n�����ȏ�� ؏ڏ�"��F�4�j� X���|���ğ���֟ ���0��@�B�T��� x�����ү䯎o��� ̯ʯP�>�t�b����� ���������Կ&� L�:�p�^ϔϦϸ��� ������� �"�H�6� l�Zߐ�~ߴߢ����� �����2� �V�D�z� h������������ �
�,�.�@�v��� ����\������� <*`N���� x���8J \(����� ���/4/"/X/F/ |/j/�/�/�/�/�/�/ �/??B?0?f?T?v? �?�?�?�?�?�?OO ��2ODO�� O�OtO�O �O�O�O�O_�O(_:_ L_
__�_p_�_�_�_ �_�_ o�_$oo4o6o Ho~olo�o�o�o�o�o �o�o D2hV �z�����
� �.��R�@�b���v� ��&OXO֏菒���� �N�<�r�`������� ̟ޟ🮟��$�&� 8�n�������^�ȯ�� �گ��� �"�4�j� X���|�����ֿĿ� ���0��T�B�x�f� �ϊϜ���������� �>�P���h�zߌ�6� �ߪ����������:� (�^�p���R���p���� ���  &��*� *�>�*���$TBJOP_G�RP 2U����  ?_���C*�	V��]�Wd������X  �*��� �,? � ���*� @&�?��	� �A�����C�  DD������>v�>\?� ��aG�:��o��;ߴAT3������A�<���MX����>��\�)?���8Q������L��>̼0 &�;iG.���Ap< � F�A�ff�v��� �):VM�.��� S>o*�@��R�Cр	����p�����ff��:�6/�?�3=3�B   �� /������>)/:�S���� <�/�/@��H�%&/и/��=� <#��
*��v�;/��ڪ!?���4B� 3?'?2	��2?hZ? D?R?�?�?�?F?�?�? �?�?OAOO�?`OzO`dOrO�O�O*�C�*����A��	V3.�00{�crxl��*P��%�%c�5Z F� �JZH F6� �F^ F�� �F�f F� �G� G5 �G<
 G^] �G� G����G�*�G�S G�; G��ER�Du�\E[� �E� F( �F-� FU` �F}  F�N �F� F�� �Fͺ F� �F�V G� �Gz Ga O9ѷ�Q�LHe�fJ4�o,b*��0c1���OH�ED_?TCH Xd�+X�2S�&�&�dA$'X�o�o*�1F��TESTPARS�  ��cV�HR�pABLE 1Yd� N`*����R�g$j�g�h�h�)�1��g	�h
�h��hHu*��h�h:�h%vRDI0n�GYk}��u	�O�#�-�?�Q�c�u�)rS�l� �z6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z���I���m�Fwͩ ��ȏڏ쏘������x)r��NUM [ ��n����2� Ep�)r_CFG Z��I����@V�IMEBF_�TTqD��e޶V�ER�����޳R� 1[8{ 8$�o*�%�Q� ��د  9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}��ߡ߳� ����������1��� E�W�i�{������ ��������/�A�S� e�w����������������+=O�_Ԗ��@��`LIoF \��D`B����DR�(FP�
�!p�!p� �d� ��MI_CH�AN� � D_BGLVL��f�ETHERAD� ?u��0`�1�_}�ROUmT�!�j!���SNMASK�Y�j255.�%S///A/S�`O�OLOFS_DI�p�CORQC?TRL ]8{��1o�-T�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OL�/6O�%OZOcPE_DE�TAI7�*PGL�_CONFIG �c������/�cell/$CID$/grp1^O@�O�O�O
__|��� G_Y_k_}_�_�_0_�_ �_�_�_oo�_CoUo goyo�o�o,o>o�o�o �o	-�oQcu ���:���� �)���_�q���������׮}N�����%�7�I�a�KOq�P�� M�����ʟܟ� �G� $�6�H�Z�l�~���� ��Ưد������2� D�V�h�z������¿ Կ���
ϙ�.�@�R� d�vψϚ�)Ͼ����� ���ߧ�<�N�`�r� �ߖ�%ߺ�������� �&��J�\�n��� ��3����������"� ��F�X�j�|���������@�User� View �I}�}1234567890����+`=Ex �e����2��B������`r��3�Oa�s����x4 >//'/9/K/]/�~/x5��/�/�/�/ �/?p/2?x6�/k? }?�?�?�?�?$?�?x7Z?O1OCOUOgOyO�?�Ox8O�O�O�O�	__-_�ON_TR �lCamera���O�_�_�_�_�_�_˂E�_o)o;n ��Uogoyo�o�o�o�)  mV�	�_�o# 5GY o}���o�������F_� mV=�k�}������� ŏl����X�1�C� U�g�y���2�D��"� ן�����1�؏U� g�y�ğ������ӯ� ����D��k��E�W�i� {�����F�ÿտ�2� ��/�A�S�e��nU Y9������������	� ��-�?�Qߜ�u߇ߙ� �߽���v�D�If�� -�?�Q�c�u�ߙ�� ���������)�;� ��D��I��������� ������)t�M�_q���N�`�9 3��0B�� Sx�1����P�//�J	oU0� U/g/y/�/�/�/V�/ �/�/�?-???Q?c? u?/./tPv[?�?�? �?OO(O�/LO^OpO �?�O�O�O�O�O�O�? oU�k�O:_L_^_p_�_ �_;O�_�_�_'_ oo $o6oHoZo_;%N��_ �o�o�o�o�o �_$ 6H�ol~��� �moe��]�$�6� H�Z�l�������� ؏���� �2��e &�ɏ~�������Ɵ؟ ���� �k�D�V�h� z�����E�e��5�� ��� �2�D��h�z� ��ׯ��¿Կ���
���  ��9�K� ]�oρϓϥϷ�����<����   �� 5�G�Y�k�}ߏߡ߳� ����������1�C� U�g�y�������� ����	��-�?�Q�c� u��������������� );M_q��  
��(  }�-�( 	 � ������# 35G}k���:�
� �Y�
/ /./��R/d/v/�/�/ �/����/�/�/A/? 0?B?T?f?x?�/�?�? �??�?�?OO,O>O �?bOtO�O�?�O�O�O �O�O_KO]O:_L_^_ �O�_�_�_�_�_�_#_  oo$ok_HoZolo~o �o�o�_�o�o�o1o  2DVh�o�o� ��	��
��.� @��d�v�������� Џ���M�*�<�N� ��r���������̟� %���&�m�J�\�n� �������ȯگ�3� �"�4�F�X�j����� ������ֿ����� 0�w���f�xϊ�ѿ�� ���������O�,�>� Pߗ�t߆ߘߪ߼��� �����]�:�L�^��p����߻@  ����������� ���"frh:\�tpgl\robots\crx!��10ia_l.xml��D�V�h�z������������������ ��0BTfx� �������� ,>Pbt��� �����/(/:/ L/^/p/�/�/�/�/�/ �/��/?$?6?H?Z? l?~?�?�?�?�?�?�/ �?O O2ODOVOhOzO �O�O�O�O�O�?�O
_ _._@_R_d_v_�_�_ �_�_�_�O�_oo*o <oNo`oro�o�o�o�o��o�n �6� |���<< 	� ?��k!�o; iOq����� ����%�S�9�k�@��o�����я�����(�$TPGL_�OUTPUT �f������ �&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��������į�p�ր2�345678901�����1�C�K� ���r���������̿ d�п��&�8�J��}T�|ώϠϲ���\� n�����0�B�T��� bߊߜ߮�����j��� ��,�>�P����߆� ��������x���� (�:�L�^���l����� ������t���$6 HZlz��� ���� 2DV h ����� ��/./@/R/d/v/ /�/�/�/�/�/�/�/~ۂ $$�� ί<7*?\?N?�?r?�? �?�?�?�?�?OO4O &OXOJO|OnO�O�O�O �O�O�O_�O0_"_T_}�an_�_�_�_�_�_��]@�_o	z ( 	 V_Do2o hoVo�ozo�o�o�o�o �o
�o.R@v d������� ��(�*�<�r�`����ܦ�  <<I_ˏݏ����� ��:�L�֪��}���)� ��ş�������k�� C�ݟ/�y���e����� ��������-�?�� c�u�ӯ]�����W�� �Ϳ��)χ���_�q� �yϧρϓ�����M� �%߿��[�5�Gߑ� ��߫���s����!� ��E�W��?���9� ��������i���A� S���w���c�u���� /�����=) s�����U�� �'9�!o	 [�����K� #/5/�Y/k/E/w/�/ �/�/�/�/�/?�/ ?U?g?�/�?�?7?�?��?�?�?	OO��)�WGL1.XML��_PM�$TPOF?F_LIM ���P����^FNw_SVf@  �T�xJP_MON �g��zD�P��P2ZISTRTC�HK h��xF�k_aBVTCOMP�AT�HQ|FVWV_AR i�M:X.�D �O R_�P��BbA_DEFPROG %�I�%TELEO�Pi_�O_DISP�LAYm@�N�RIN�ST_MSK  ��\ �ZINU�SER_�TLCK�l�[QUICKM�EN:o�TSCRE�Y`��Rtpsc�Tat`yixB��`_�iSTZxIR�ACE_CFG �j�I:T�@	�[T
?��hHNL� 2k�Z���aA[  gR-?Qcu�����z�eITEM �2l{ �%$�12345678�90 ��  =<�
�0�B�J�  !P�X�dP���[S� ��"���X�
�|��� W���r�֏����.�� 0�B�\�f�����6�\� n�ҟ��������>� ��"���.�����ί R����Ŀֿ:��^� p�9ϔ�Tϸ�xϊ�� ���d���H��l�� >�Pߴ�\�������v�  ������h�(�ߞ� ��4�L��ߦ����� @�R��v�6���Z�l� ��������*���N� �� ������������ X���J
n ���b��� �"4F�/|</ N/�Z/���//�/ 0/�/?f/?�/�/e? �/�?�/�?�?�?,?�? P?b?t?�?�?DOjO|O �?�OOO(O�O�O^O _0_�O<_�O�O�_�O �__�_�_H_�_l_~_�Go�dS�bm�oLjψ  �rLj 8�a�o�Y
 �o�o��o�o{jUD1:�\|��^aR_G�RP 1n�{?� 	 @�PR d{N�r����~��p���q+��<O�:�?�  j�|� f����������ҏ� ���>�,�b�P���t�0��������	e����\cSCB 2ohk U�R�d�v����������Я�RlU�TORIAL �phk�o-�WgV_C�ONFIG q�hm�a�o�o��<�OUTPUT rhi}�����ܿ�  ��$�6�H�Z�l�~� �Ϣϴ�z�ɿ���� � �$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ����*<N` r�������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/��/�/??0? B?T?f?x?�?�?�?�? �/�?�?OO,O>OPO bOtO�O�O�O�O�?�O �O__(_:_L_^_p_ �_�_�_�_�_f�x�ǿ oo,o>oPoboto�o �o�o�o�o�o�O (:L^p��� ����o ��$�6� H�Z�l�~�������Ə ؏��� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я��� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t�����������������X���#�� N�_r����� ��&8J�� n������� �/"/4/F/X/i|/ �/�/�/�/�/�/�/? ?0?B?T?e/x?�?�? �?�?�?�?�?OO,O >OPOa?tO�O�O�O�O �O�O�O__(_:_L_ ^_oO�_�_�_�_�_�_ �_ oo$o6oHoZok_ ~o�o�o�o�o�o�o�o  2DVgoz� ������
�� .�@�R�d�u������ ��Џ����*�<� N�`�q���������̟ ޟ���&�8�J�\��k��$TX_SCREEN 1s%� �}�k�����ӯ���	���Z��I�[�m�� �����,�ٿ���� !�3Ϫ�W�ο{ύϟ� ������L���p��/� A�S�e�w��� ߭߿� �������~�+��O� a�s���� ���D� ����'�9�K����� ������������R��� v�#5GYk}�����$UALRM_MSG ?����� �n��� 	:-^Qc������� /�S�EV  ��2&�ECFG �u����  �n�@�  Ab! �  B�n�
  /u����/�/�/�/�/ �/??%?7?I?W7>!�GRP 2vH+; 0n�	 /�?�� I_BBL_N�OTE wH*T��lu�䐠w�T �2DEF�PRO� %� (%�Ow�	OBO-BTELEOPGO #O�O�O�O�O�O�O�O�_�O&_�?�0FKE�YDATA 1x<���0p W'n��?�_�_z_�_�_�Z�,(�_on�(POOINTo>o �_�coJo�ono�o�o d?TOUCHU`O�o �o�o7[mT �x�������!��E��Z��/�frh/gui/�whitehome.pngQ�����س�ŏ׏�h�pointz���/�A� S��\���������ȟ ڟi����"�4�F�X� �|�������į֯e��h�touchup���/�A�S�e��}h�arwrg�� ����ÿտ�n��� /�A�S�e����ϛϭ� �������τ��+�=� O�a�s�ߗߩ߻��� ���߀��'�9�K�]� o����������� ���#�5�G�Y�k�}� T������������ �1CUgy� �����	� ?Qcu��(� ���//�;/M/ _/q/�/�/�/6/�/�/ �/??%?�/I?[?m? ?�?�?2?�?�?�?�? O!O3O�?WOiO{O�O �O�O@O�O�O�O__ /_�OS_e_w_�_�_�_ �_N_�_�_oo+o=o �_aoso�o�o�o�oV���k�b�����o}�o8J$v,6�{.���� �����/��S� :�w���p�����я� ʏ��+��O�a�H� ��l�������ߟ�� �'�9�Ho]�o����� ����ɯX�����#� 5�G�֯k�}������� ſT������1�C� U��yϋϝϯ����� b���	��-�?�Q��� u߇ߙ߽߫�����p� ��)�;�M�_��߃� ��������l��� %�7�I�[�m������ ��������z�!3 EWi������ ���П/AS ew~����� �/�+/=/O/a/s/ �//�/�/�/�/�/? �/'?9?K?]?o?�?�? "?�?�?�?�?�?O�? 5OGOYOkO}O�OO�O �O�O�O�O__�OC_ U_g_y_�_�_,_�_�_ �_�_	oo�_?oQoco uo�o�o�o:o�o�o�o )�oM_q� ��6�����h%�7�9�����b�t���^�������,��돞� ���3�E�,�i�P��� ����ß�������� �A�S�:�w�^����� ��ѯ����ܯ�+�
 O�a�s��������Ϳ ߿���'�9�ȿ]� oρϓϥϷ�F����� ���#�5���Y�k�}� �ߡ߳���T������ �1�C���g�y��� ����P�����	��-� ?�Q���u��������� ��^���);M ��q������ l%7I[� �����h� /!/3/E/W/i/@��/ �/�/�/�/�/�?? /?A?S?e?w??�?�? �?�?�?�?�?O+O=O OOaOsOO�O�O�O�O �O�O_�O'_9_K_]_ o_�__�_�_�_�_�_ �_�_#o5oGoYoko}o �oo�o�o�o�o�o �o1CUgy� �����	��� ?�Q�c�u�����(��� Ϗ������;�M�@_�q�������~ ����~ ����ҟ���Ο�*��, �[���f������� ٯ�������3��W� i�P���t���ÿ��� ο��/�A�(�e�L� �ϛ�z/��������� �(�=�O�a�s߅ߗ� ��8���������'� ��K�]�o����4� ���������#�5��� Y�k�}�������B��� ����1��Ug y����P�� 	-?�cu� ���L��// )/;/M/�q/�/�/�/ �/�/Z/�/??%?7? I?�/m??�?�?�?�? �?���?O!O3OEOWO ^?{O�O�O�O�O�O�O vO__/_A_S_e_�O �_�_�_�_�_�_r_o o+o=oOoaosoo�o �o�o�o�o�o�o' 9K]o�o��� �����#�5�G� Y�k�}������ŏ׏ ������1�C�U�g� y��������ӟ��� 	���-�?�Q�c�u��� �����ϯ������0���0���B�T�f�>�����t�,��˿~��ֿ �%��I�0�m��f� �ϊ�����������!� 3��W�>�{�bߟ߱� ���߼�����?/�A� S�e�w������ ��������=�O�a� s�����&��������� ��9K]o� ��4���� #�GYk}�� 0����//1/ �U/g/y/�/�/�/>/ �/�/�/	??-?�/Q? c?u?�?�?�?�?L?�? �?OO)O;O�?_OqO �O�O�O�OHO�O�O_ _%_7_I_ �m__�_ �_�_�_�O�_�_o!o 3oEoWo�_{o�o�o�o �o�odo�o/A S�ow����� �r��+�=�O�a� ���������͏ߏn� ��'�9�K�]�o��� ������ɟ۟�|�� #�5�G�Y�k������� ��ůׯ������1� C�U�g�y�������� ӿ������-�?�Q��c�uχ�^P���>^P������� �ͮ���
���,��;� ��_�F߃ߕ�|߹ߠ� ���������7�I�0� m�T��������� ���!��E�,�i�{� Z_������������� /ASew� ������+ =Oas��� ���//�9/K/ ]/o/�/�/"/�/�/�/ �/�/?�/5?G?Y?k? }?�?�?0?�?�?�?�? OO�?COUOgOyO�O �O,O�O�O�O�O	__ -_�OQ_c_u_�_�_�_ :_�_�_�_oo)o�_ Mo_oqo�o�o�o�o�� �o�o%7>o[ m����V� ��!�3�E��i�{� ������ÏR����� �/�A�S��w����� ����џ`�����+� =�O�ޟs��������� ͯ߯n���'�9�K� ]�쯁�������ɿۿ j����#�5�G�Y�k� ���ϡϳ�������x� ��1�C�U�g��ϋ߀�߯����������`�����`���"�4�F��h�z�T�,f���^������� ��)��M�_�F���j� ������������ 7[B�x� ����o!3E Wixߍ���� ���///A/S/e/ w//�/�/�/�/�/�/ �/?+?=?O?a?s?�? ?�?�?�?�?�?O�? 'O9OKO]OoO�OO�O �O�O�O�O�O_�O5_ G_Y_k_}_�__�_�_ �_�_�_o�_1oCoUo goyo�o�o,o�o�o�o �o	�o?Qcu ��(����� �)� M�_�q����� ���ˏݏ���%� 7�Ə[�m�������� D�ٟ����!�3� W�i�{�������ïR� �����/�A�Яe� w���������N���� ��+�=�O�޿sυ� �ϩϻ���\����� '�9�K���o߁ߓߥ� ������j����#�5� G�Y���}������ ��f�����1�C�U��g�>�i��>������������������,��? &cu\���� ���)M4 q�j����� /�%//I/[/:�/ �/�/�/�/�/���/? !?3?E?W?i?�/�?�? �?�?�?�?v?OO/O AOSOeO�?�O�O�O�O �O�O�O�O_+_=_O_ a_s__�_�_�_�_�_ �_�_o'o9oKo]ooo �oo�o�o�o�o�o�o �o#5GYk} �������� 1�C�U�g�y������ ��ӏ���	���-�?� Q�c�u�����p/��ϟ �����;�M�_� q�������6�˯ݯ� ��%���I�[�m�� ����2�ǿٿ���� !�3�¿W�i�{ύϟ� ��@���������/� ��S�e�w߉ߛ߭߿� N�������+�=��� a�s�����J��� ����'�9�K���o� ����������X����� #5G��k}���������}������@&�HZ4,F/ �>/�����	/ �-/?/&/c/J/�/�/ �/�/�/�/�/�/?�/ ;?"?_?q?X?�?|?�? �?���?OO%O7OIO XmOO�O�O�O�O�O hO�O_!_3_E_W_�O {_�_�_�_�_�_d_�_ oo/oAoSoeo�_�o �o�o�o�o�oro +=Oa�o��� ������'�9� K�]�o��������ɏ ۏ�|��#�5�G�Y� k�}������şן� �����1�C�U�g�y� �������ӯ���	� �?-�?�Q�c�u����� ����Ͽ���Ϧ� ;�M�_�qσϕ�$Ϲ� �������ߢ�7�I� [�m�ߑߣ�2����� �����!��E�W�i� {���.��������� ��/���S�e�w��� ����<������� +��Oas��� �J��'9 �]o����F����/#/5/G/��$UI_INUS�ER  ����h!� � H/L/_ME�NHIST 1y�h%  �( u ��+�/SOFTPAR�T/GENLIN�K?curren�t=editpa�ge,TELEOP,1�/�/?!?�y)�/�%menu�"1133�/}?�?�?γ? �'E?W>71@l?�?O#O5O�(�?W?54�?�O�O�O�O IO[OmBk?__+_=_�?�O�!2�O�_�_�_��_�Oa_c348,2`�_o$o6oHo��Io�no�o�o�o�o�o�� \a�!\o�o/A SVow����� `���+�=�O�� ���������͏ߏn� ��'�9�K�]�쏁� ������ɟ۟j�|�� #�5�G�Y�k������� ��ůׯ��o�o�1� C�U�g�y�|������� ӿ������-�?�Q� c�uχ�ϫϽ����� ��ߔ�)�;�M�_�q� ��ߧ߹�������� ��7�I�[�m���  ������������� �E�W�i�{������� ����������A Sew���<� ��+�Oa s���8��� //'/9/�]/o/�/ �/�/�/F/�/�/�/? #?5? �2�k?}?�?�? �?�?�/�?�?OO1O CO�?�?yO�O�O�O�O �ObO�O	__-_?_Q_ �Ou_�_�_�_�_�_^_ p_oo)o;oMo_o�_ �o�o�o�o�o�olo�%7I[F?���$UI_PANE�DATA 1{�����q�  	�}  �frh/cgtp�/flexdev�.stm?_wi�dth=0&_h�eight=10��p�pice=TP�&_lines=�15&_colu�mns=4�pfo�nt=24&_p�age=whol�e�pmI6)  r3im�9�  �pP� b�t������������ Ǐ��(�:�!�^�E� ����{�����ܟ�՟��I6� � � [0 � J�O�a�s��������� ͯ@����'�9�K� ��o���h�����ɿۿ ¿���#�5��Y�@� }Ϗ�vϳ�&��Ɠs �����)�;�Mߠ� q�䯕ߧ߹������� V��%��I�0�m�� f������������ !��E�W����ύ��� ��������:�~�/ ASew��� ��� =$ asZ�~��� �d�v�'/9/K/]/o/ �/��/�/*�/�/�/ ?#?5?�/Y?@?}?�? v?�?�?�?�?�?O�? 1OCO*OgONO�O�/ �/�O�O�O	__-_�O Q_�/u_�_�_�_�_�_ 6_�_o�_)ooMo_o Fo�ojo�o�o�o�o�o �o%7�O�Om �����^_� !�3�E�W�i�{���� ��Ï��������� A�S�:�w�^������� џDV��+�=�O� a�������
���ͯ߯ ���|�9� �]�o� V���z���ɿ���Կ �#�
�G�.�k�ޟ�}�|ϵ����������)��4ߧ�#�`�r� �ߖߨߺ�!������ ����8��\�C��� y������������������$UI_P�OSTYPE  ���� �	 �s�B�QU�ICKMEN  �Q�`�v�D�RE�STORE 1|���  '������������mASew �,������ +=Oan� ����//� 9/K/]/o/�/�/6/�/ �/�/�/�/�??0? �/k?}?�?�?�?V?�? �?�?OO�?COUOgO yO�O6?@O�O�O.O�O 	__-_?_Q_�Ou_�_ �_�_�_`_�_�_oo )o�O6oHoZo�_�o�o �o�o�o�o%7 I[�o����ށ�SCRE��?���u1sc���u2�3�4��5�6�7�8���sTATM�� �����:�USER��p��rT�p�ksT���4��5��6���7��8��B�NDO_CFG }Q�X����B�PDE����None���v�_INFO �2~��)���0%�D���2�s�V��� ����͟ߟ��'� 9��]�o�R���z���OFFSET 	�Q�-���hs��p �����G�>�P�}� t���Я��׿ο�� ��C�:�L�^Ϩ����͘���
����av���WORK �!�����.�@ߢ�u��UFRAME  ����RTOL_ABRT������ENB�ߣ�GRP� 1�����Cz  A����� �*�<�N�`�r�����U�����MSKG  �)���N��%!��%z����O_EVN������+�ׂ3�«
 h��UEV��!�td:\eve�nt_user\��u�C7z���jpF���n�SPs�x�spotweld��!C6��������!���G|'�� 5kY���� �>���1� Ug���/�� 	/^/M/�/-/?/�/c/ �/�/�/�/$?�/H?�/4:J�W�3�����#8C?�?�? �?�? �?�?O+OOOOaO<O �O�OrO�O�O�O�O_ �O'_9__]_o_J_�_��_�_�$VALD_CPC 2�«� �_�_� w��qd�R�*o_o(qo��hsNbd�j�` ��i�da{�oav�_�o oo3BoWi{�o �o�o�o��o� PA�0�e�w���� ������(�=� L�a�s�
�������ʏ �����$�ޟH�:� o���������ڟ؟� ���� �2�G�V�k�}� ������¯ԯ���� �.��R�S�yϋϚ� ���������	��*� <�Q�`�u߇ߖϨϺ� ��������&�8�M� \�q���߶���n� �����"�4�F�[�j� �������������� �!0�B�Wf�{� ���������� ,>teT��� ����/+/: La/p�/�/./�� ���//'?6/H/? l/^?�?�?�/�/�/�/ �/?#O�?D?V?kOz? �O�O�?�?�?�?�?_ O1_@ORO9_vOw_�_ �_�O�O�O_�__-o <_N_`_uo�_�o�o�_ �_�_�_o&o;Jo \oq�o����o�o �o� �"7�FXj ���������� �!�0�E�T�f�{��� ����ßҏ����
� ,�A�P�b�����x��� ��Ο�����(�*� O�^�p���������R� ܯ� ��Ϳ6�K�Z� l�&ϐ��Ϸ���ؿ� ��"� �2�G���h�z� �ߞϳ���������
� �1�@�U�d�v�]�� �����������,�� <�Q�`�r������ ��������&�;J� _n��������� �����$F[j |������� 0E/Ti/x� �/��/�/�/�// ,/.?P/e?t/�/�/�? �?�?�?�/??(?:? L?NOsO�?�?�O�?�O �OvO OO$O6O�OZO o_~O�OJ_�O�_�_�_��O_ _F_D_V[�$�VARS_CONFIG ��P�xa  �FP]S�\lCM�R_GRP 2�Nxk ha	`��`  %1: �SC130EF2# *�o�`]T�VU�PY�h`�5_Pa�?�  A@%pp:*`�Vn No9xCVXdv��a���<uA�%p�q��_R��_R B���#�_Q'�� H��l�;���{����� ؏ÏՏ�e��D�/��A�z�-�����ddIA�_WORK ��xeܐ�Pf,�		�Qxe���G��P ���YǑRT�SYNCSET � xi�xa-�WINURL ?=�`������������ȯگSIONT�MOU9�]Sd� ���_CFG ��S۳�S��P�` F�R:\��\DAT�A\� �� wMC3�LOG@�   UD13��EXd�_Q' ?B@ ����x��e_ſx�ɿ�VW �� n6  ���VV��l�q  =���?��]T<�y�Y�TRAcIN���N� 
gCp?�CȞ��TK�t��b�xk (g� ����_��������� U�C�y�g߁ߋߝ߯߸�����_GE��nxk�`_P�
�PX�RꋰRE��xe\*�`hLEX�xl�`1-e�VMPHASE  xe�c�ecRTD_�FILTER 2]�xk �u�0 ����0�B�T�f�x� ����VW�������� �$6HZl_iS�HIFTMENU� 1�xk
 <b�\%������� ���=&s J\��������'/�	LIV�E/SNA�c%?vsfliv��9/W��� 7�U�`\"menur/w// �/�/�����]��+MO��y��5`h`KZD4�V�_Q<���0��$WAITDINEND��a2>p6OK  �i�<����?S�?�9TIM.�����<Gw?M �?*K�?
J�?
J�?�8RELE��:G6p3x���r1_ACTO �9Hܑ�8_<� ��ԙ�%�/:_af�BR�DIS�`�N�$�XVR��y���$ZABC�b1�NS; ,��j�I��2B_ZmI1�@VSP�T �y��eG�
�*�/o�*!o�7o�WDCSCHG� �ԛ(��P\g�@�PIPL2��S?i��o�o�o�ZM�PCF_G 1��ii�0'¯S;MsҖS��i��p'���g��e2��  �?5���3|Y�=�y�2�/��6�B��65�=���6
*��~�`C���B���C�_��I�1�q>�����F��=�5�[�����c��������Z�~���Ï��>��0C+�r?�|�2��ڏ�ӈ�����*�@�N� x��$�6�H�0N�`�ȌTp���o�_C_YLIND�� {� Х� ,(  *=�N�G�:�w�^����� ��ѯ� ��7����<�#�5�r� ����������޿y�_� ���8�ύ�nπ��r�ã wQ �5 �����S�����(��h��X�זr�A���SPHERE 2���ҿ��"ϧ��� ���P�c�>�P�̿t� ��ߪ�����'�� �]�o�L���p�W�i�������������PZZ�F �6