��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1CES0�2eG �� QA> �1
 � $SOFT��T_ID�2TOT_AL_EQ 0�1�@N" �@U SPI�
 �0^�EX�3CR�E -DdBSIG�J@dOvK�@PK�_FI90	$�THKY"WPAN�E�D � DUMMY1dIT1TU�4QQ!Rx1R�� � $TIT91� ��� �Td�TP0�ThP�T5�V6�VU7�V8�V9�W0�W��WOQ�U�WgQ�U�W1��W1�W1�W1�W2��R �@SBN_CmF�!@$<!�J� ; ;2�1_CM�NT�$FLAsGS]�CHEK"{$�b_OPTJB��@� ELLSETUP  `@�HO8@9 PR�1%x�c#�aREPR�hu0D+�@��b{u[HM9 MN�B;1^ UTOBJ U��0 49DoEVIC�STI/@��� �@b3�4pBܢd�"VAL�#IS�P_UNI�tp_�DOcv7�yFR_F�@|%u13��A0s�C_WA�t,q�z�OFF_T@N�DEL�Lw0dq�1��Vr?^q�#S?�o`Q"U�t#*�Q�TB��%�MO<� �E � [�M�����REV��BIL��]aXI�� v�R  �!D�`��$NOc`M�|�� ��ɂ/#ǆ� ԅ����X�@Ded �p E RD_E���h�$FSSB�6�`KBD_SEV�uAG� G�2Q"!_��2b�� V!�k5�p`(��C�0q_ED|� � � t2d�$!S�p-D%$� ��#�B�ʀ_�OK1��0] P_C�� ʑ0t��U �`LACI�!�a�Y�� ��qCOMM� # $D
� ��@���J_�\R�0BIGALL;OW� (Ku2:-B�@VAR���!|�AB ���BL�@� � ,K�q��r�`S�p�@M_O]�˥��CCFS'_UT��0 "�A�Cp'��+pXG��b�0� 4� IMCM ��#S�p�9���i �_�"t\b���M�1 h$�IMPEE_F�s���s��� t����D_(�����D��F��� �_����0 aT@L��L�DI�xs@G�� �P�$I�'�ƺذFed X@G�RU@��Mb�NF�LI�\Ì@UIR�E�i42� SWIYTn$`0_N�`S 2�CF�0M� 	�#u�D��!��v`(����`J�tV��[ �E��.p�`�ʗELBOF� �շ �p`0���3����� F�2T��A`�rq1�J1��z _To!@��p��g���G�� �r0WARNM�p#tC�v`�ç` �� COR-UrF�LTR��TRAT�9 T%p� $AC�CVq��� ��r$�ORI�_&�RTr��S<�]`CHG�0I���TW��A��I'�T��HK�� �202�a�1��HDR�2��2B�2J; S���3��U4��5��6��7��8��9��׀
 �2w @� TRQ��$vf��'�1�<�_�U<�G��0COec  <� P�b�t�53�>B_�LLEC��!>~�MULTI�4�"�u�Q;2�CHILID��;1_��@T�w "'�STY92	r��=��)2���x����ec# |r0 56$J ђ��`�L��uTO���E^	EXTt����2���22"]����$`@D	�`&��ղ���� %�"��`%�a�k�����s=����& '�E�Au��Mw�9 n�% ��TR�� ' L@U#�9 ���At�$JO�B����PM�}IG��( dp���� ��^'#j�~ǝ�p{OR�) t$�3FL�
RNG%Q@�TBAΰ �v&r�* `1t(��0 �x!�0�+aP�p�%4��*�Ё͐U��q�!�;2J��_R��>�C<J��8&<J D`5C�F9���x"�@J�P_�p�7p+ \@RaO"pF�0��IT�s�0NOM��>Ҹ4s(�2�� @U<PPgў�P8,|Pn��0�1P�9�͗ RA���pl�?C�� �
$TͰ.tMD3�0T��pQU�`�΀+AHlr>�T1�JE�1\�J����PQ��\Q��hQCY�NT�P��PDBG�D̰�0-���PU�6$$Po�|�u�AX�����TAI�sB�UF,�]��A�1. �����F�`PI|�U-@PvWMuXM�Y��@�VFvWSIMQ�STO�q$KEE�SPA��  ?B�BP>C�B�2��/�`�ˏMARG�u2�F�ACq�>�SLEW�*1!0����
ۅ2M�CW$0'���pJqB�Ї�qDECj��exs�V%1 �Ħ�CHNR�MP�s�$G_@�gD�_x�@s��1_FP�5�@TC�fFӓC�Й���qC��+�VK�*��"�*�JRx���SEG�FR$`IOh!�0S�TN�LIN>�csP!VZ҅2�A�D2����r 2��hr�r�1��3` +^?���� �q�`��q|`�����t8��|aSIZ#�!� �T�_@%�I��qRS�*s��2y{�Ip{�pTpLF�@�`ΰ�CRC����CC TѲ�Ipڈ�a���bL�MIN��a1순�*��D<iC �C/����!uc�OP4�n j�EVTj���F��_!uF���N����|a��=h?K�NLA�C2�AV'SCA�@A�s�1�4�  cSaF�$�;�Ir �4(�@�05��	D-O o%g��,,m�����ޟ��BRC�6� n���sυ�U���R�0HANC��$cLG��ɑDQ$t��NDɖ��AR۰N���aqg��ѫ�X�ME`��^�Y�[PS�RAg�X�AZ�П���rEOB�FCT��A��`�2rt!Sh`0ADI��O��y�s"y�n!�������~#C�G3t!��'BMPmt@�Y�3�a�fAES$�����W�_;�BAS#XYOZWPR��*�m!��	�1U�87 � ƀI@d���8\�p_C:T���#���_L
 � 9 ���C�/�(zJ�L%B�$�3�D��5��FORC�b�_;AV;�MOM*�q�	SaԫBP`Ր�y�HB�P�ɀE�F����AY�LOAD&$ER �t&3�2�Xrp�!�*zR_FD�� /: T`I�Y3���E�&��Ct��M-S�PU
$(kpLD��9 �b�;�Bn�	EVId�
�޸!_IDX��$ ���B@X�X<&��SY5�  �H�OPe�<��ALAR�M��2W�r���0=C h�@Pnq�`M\q�J@$PL`A&�M#�$�`��� 8�	����V�]�0��U�PM�{�U��>�TITu�
%�![q�BsZ_;���? �B� pQk��6NO_HEADE^az��}ѯ ��`􂳃���dF�ق�t���@�@��uCIRTR�`��ڈ�L��D�CB@4�RJƱ��[Q���A��2>���OR�r��Ox����T`UN_OO�Ҁ$����T���J��I�VaC|q
� OPXWOY���B��$SKADR��D�BT�TRL��C��րfpbDs��~ГDJj4 _�DQX}��PL�qwb#WA���WcD�A���A=�2�UMM3Y9��10����DB����D;[QP�R��*M�Z���E� O�Y1$�a�$8��L)FL!/��9����0GG/�_cPC�1Hf/x$E+NEA@Tf�I�/_c��RECOR`"J�H @ �E$L�#F$#PR��`�+jp��nq�_D$�qPROSS]�
����R�r�` u�$TRIyG96PAUS73>ltETURN72�+MR:�U 0Ł0�EW$��`SIGNsALA�QR$LA�м�5�1G$PD�'H$Pİ�AI�0�Ab�C�4�C��DO��D�2�!�6GO_oAWAY2MOZq��Z�W DCS��CwSCBg�K Իa\#���ERI�0Nn�!T�`$�����FCBxPL�@QBGAGE�� �P��ED|BD�wA[CD�OF�q[F0�FoC��MPMAB0XoC�?$FRCIN��2Dxk��@��$NE�@��FDL8�� L� ����=��Rw��_��P� OVR1�0���lҠ�$E�SC_�`uDSB�IO����pTe�E�VIB�� `s��Z�8�V��pSSW��$�&VL��:�Lk��X����ѣ�bQ����US�C�P��A=�	Q��MP1%e&S*`�(bt`:'c5۳ESUd�� -cWg&SWg?cWd�����Wd��Wd.���AUT�O$�Ya҃�ac�SB ����-d��&SwB[���GB�f$VOLTr�g ��  � GAOD!�q���@:ЗORQҀKra�$DH_THE&0��Rgp� qtnwALPAHnt��o��w0 Vp]�$�.�Ra�[��s�5 �`r�CQ#BUD�S� %F1M��sV
���;��Lb�tk����BRTHR��L��T(`�Z��VɖL��DE  �1��2�⋅�������� kѯ�aәTt0V�ꆸ� �����̈Я�-�"��N~��sS2����IwNHB��ILTG0 ɡ�T?��3$�w��E���PqQxQ�TqPe��0Y�AF}�O�ນ�� ڗ��qPڳē��`��bPܙ���PL?�x��3���TMOU�� ēS���� ��s�/�S1H8���O�Aܙ��I�����CDIƑ˩o�S#TI��գ�O:ҋ�,0���AN��Qg`�S��+r�#x$�Ј���w�_����PR	A�P`vC����GMCNeQe�����VERS��r�oPIw�FPåǲШ۷-G.�DN��G>���B��F�2�Ƿ�Mʪ7�F��_�MN�D ̠,����d�{ƭa����OB���U˱z���DI���#���3� ����A���w�Fx���3�ON�5��Q��VAL�CR[�_�SIZ��b�;Qn�REQ�Rb��]2b���CHq�΂�ڃ��`������:�n�S_U���X��wWFLG����wU$CV�iM8GP�QδFLXP�92`3R�u���EAL�P�-�C	��+rT��W���� �R�c���NGDMS7� ��K>S��P_M'0h�STW`v������AL�P ���Q���U���U�IAG,�o��d�U�J-�T"A-`� �� �A�����H`��Q`��6��Pq_D&��1s ��.�P�F�>2�=T�� ?7 @1A>��#�#L��?_=i @@>�LD�c���0�FRI�0 `Ѐ��1}ѲIV\1�*�^1�UP`��a��C�LW��
`�L=S&-c&&S�C .w�� L���!����d�Q$w�҇��$w�����
�P�5R�SM���V0h b� r��d^2AW�a�_TRp}�8@NS_PEA����< ��$�SAVG�8�6G]%8���CAR �`0�!�$���"CRa����$ d�#E�@��"STD���!Fpo��'�QOF��%��"RC���&RC۠�(F��2A�R#7���%, gMEA�Q_�a��
QQ�(�al2��u4Ib�r7�I�R�9wQ�7�8M�/��!CpR�  ��p�2F<�SDNX�a0 
 W2QM P $Mi� �s$cA�$C�cm�9����4�AT�0CY_ N LS!IG1x'yB��y@@H2Y�NO�����SDEVI�@ �O@$�RBT�:VSP�3�CuT�DB�Y|�A	W`3CHNwDGDAP H@�GRP�HE iXL��U��VS�Fx2��DL1p Q6ROp��sFB�\]�FEN�@���S��ChAR �d�@DOd�PMCSb�P薇P�R��HOTSWz42�D�MpELE�1/e��8C8`�RS T�@��`�r� hf��`OL�GCHA�Fk�Fs����C�A@T � �$MDLUb 2S@�E���q�6�q	0P�i�c�e�cJ��	u�ݢ�#~5t+w�PTOb��� �b�5_C�SLAVS� U;  ��INP �	V��ЊyA_;�ENU�AV $R�PC_T�q�2 1bL�w���tSHO+� WA ���A�a�q�2�rh�v�u�v�sCF� X` ,f��r�OG gE��%D�,h�J`C�Iߣi�cMA��D�x AY?�9W� p�NTV	�D�sVE�0@�SKI��!T�`g?Ň2�� JZs�! Cꆻ��f��_SV/ �`XC�LU��H���ON�L��'�Y�T��OT�:eHI_V,11 AoPPLY��HI4`�;�U�_ML�� ?$VRFY8�	�zU�M{IOC_I�D��J 1/��߃O�@�X�LSw"`@$DUMMY4���ڑz�Cd L_TP��p��kC��^1CNFf����E��@T�y� D�_#UQ_��ݥ�YPCP��=�� ������aD���� Y 9+�
0RT_;P��~T��CCb Z�r�TE���=�פr�DG�@[ D��P_BAe`Lkc�!��_���H�Md��E �\�pAb=cAR�GI�!$���`[ܶ��tSGNA] q��`U��IGN��X���� ��V��|����ANNUN���&�˳�EU�J'�ATCH��J��y��t^ <@g�����&:c$Va����X��qqEF] I��_ _ @@FͲ�ITb�	$TOT�i �C�O�c� @EmM�@NI�a`tB���c���A>���D{AY@CLOAD�D`\�n������EF7�+XI�Ra��K����O%��a�ADJS_R�!@b��>�H2�"[�
 c�%��`	a͠MPI�J��DH�8��?�Ac 0��ѐ��� ��Z�ϡ�U|i ��CTRL� �Yp d��TRA�8 ?3IDLE_PAW  �Ѡ��Q��V�G�V_���`c ��o�;Q@e� 1q$��6`<cTAC-3@��P�LQ�Z�Rz�\ A-u:ɰSW;�A\���/J��`�b�K�OH�(OP9P; �#IRO� �"gBRK��#AB � �O������� _ ���F���`d͠, j@S�oRQDW��MS��P6X�'z��IFEgCAL�� 10^tN��V��豊�V�(0L��CP
��N� 9Yb�0FLA_#�3OVL ��HE���"SUPPO��ޑ\B�L�p��&2X�*$Y-
Z-
W-
��`/��0GR�XZ�q6�$Y2�CO�PJ�SA�X2R��*r�!��:��"&pr0��0)��f `�@CACHE��c��0�s0�LAZ SUFFI, C��Ja\��r�6��NaMSW��g 8�KEYI�MAG#TM�@S���n
2j�r��bO�CVIE��~�h �aBGL����`�C?�@� @���i��m!`STπ!� �����n����/EMAI�`N��`A�rpZ�FAU� �jH�"Jaa��U�3��a� }�k< �$I#�US�� �IT'�BUF`�r�DNB���SUBu$��DC_���J"��"SAV�%�"k�������';��P�$�UOR	D��UP_u �%��8OTT��_B`��8@�LMl�F4��C7AX�@Cv���Xu 	��#_9G���1YN_����l6���D�E��M�����T��F���caC�DI`BEDT�)@C��~�m�rI�GD�!c�&��l`������P��FZP n (�pSV� )d\�ρ�ɚ�B��o�� ����>"$3C_R�IK��kB��hD�{pRfgE.(ADS�P~KBP�`�IIM@�#�C�Aa�A��U�Gh���iCM! IP��0KC��� �DTH� �Sd�B*�T��CHS�3��CBSC��� ��V`�dYVSP�#[T_Drc/CONV�Grc[TH� �Fu F�ቐd�C�0j1��SC5�e]C�MER;dAFBC�MP;c@ETBc �p\FU DU�i ��+�~�CD�I%P702#R�EO����qWӏ�SQ��QǀSU��MSS�1ju�D4`�TB�Aa��A�1r� "�Й��4$ZO@s���l��U6�&��eP���eC�Nc�l��l�l�iGR#OU�W)��S c�MN�kNu�eNu�eNpR|b|�i�cH�pi��z
 �0CYC���s�w��c��zDEL�_D��RO�a���qVf���v{�O�2��� 1��t��:R�ua�.#�7 ���AL� �1�sˢI1¡�J0�PBX���z�ER^�T�Gbt ,!@��5���aGI1LcR1s 
L�0ԠNO��1u����������P����C�ڠ	�����ge�,��J0�0vH *	�LU�1#J�Q��V 
�[�7Az���z��z�@n�z��z�Fz�7w��8w�9w���y���1���1��1��1��1�Ě1њ1ޚ1�2R��2����2��2��U2��2Ě2њ2ޚU2�3��3��3�����3��3��3Ě3*њ3ޚ3�4���2XTF��1w6�.(�0@�f�0�U�0ŷ�e�P�FDR5�xTU VE��?1���SR���RE�F���O�VM~C)�A2�TR�OV2�DT� R�MXa�IN2���Q�2�'INDp�r�
���0�0�0Gu1��[�G`��r{�D_�[�RIV�P��b�GEAR~AI%Or�K"N�0��y�p�5`@�a�Z_�MCM� �� �F��UR�Ryǀ��!�? ��p?\nЋ�?n�ER� v�K�!�P��zI:�5PXqB�RI0%���#ETUP2_ g{ ���#TDPR�%TBp�����Ղ��"BAC�2| T(��"�4)�:%	`^B���p�IFI��b� Mc���.�PT��ޔFLUI�}c � ��K UR�c!���B�1SPx E�ESMP�p�2$��S^�?x��Jق0
3�VRT���0x$S�HO��Lq�6 AS�ScP=1��PӴBG_���-���<�FORC��g㶙d~)"FUY�1�2\�2�1I�h� p�w |��NAV�aS�������S!"~�c$VISI��6#�SCM4SE�����:0E�V�O��$����G@��$��I���@�FMR}2��� � 5`�r�@�� ߠ2�I�9 F�"�_�~��LIMIT_1�dC_LM�����͟DGCLF����DMY�LD����5�Ɣ������M�Fc��D u	 T�F9S0Ed� P��Q|C�0$EX_Q�hQ1i0�P�aQ3��5��GoQ���� ����RSW�%OyN�PX�EBUG�L�'�GRBp�@U�S�BK)qO1L� ��POY 
)��P���M��OXta`S�M��E�"�a���`_?E � o�F�^��TERMZ%�c%Nd�ORI�1_ �|)KSMepO��_ �|&ȃ��`�(�c%I�UP�>� �� -����b���q#� ����G�*� ELTO0Q�p�0�PFIrc�1�Y��P�$�$�$U;FR�$��1�L0e� OTY7�PT�4q�k3NST�pP�AT�q4PTH	J�a`EG`*C�p1ART� !5� y2�$2REL�:)ASHCFTR1�1�8_��QR�Pc�& � $�'@�� ��s�1 @�I�0�U�R��$P�AYLO�@�qDYN_k�����1|��'PERV��RA��H ��g7�p�2�J�E-��J�RC���ASY�MFLTR�1WJ*7����E�ӱ1�I��aUT�pbA�5��F�5P�PlC�Q1FO5R�pM�I!���W��/&�0F0�cs�H��Ed� �m2XN���5`OC1!>?�$OP�����c�����bRE�PR.3�1a�F��3e��R�5e�X�1>(�e$PWR��_���@R_�S�4��et�$3UD��e��Q72 ����$H'�!^�`ADDR�fHL!�G�2�a�a�a���R���U�� H��SSC����e-��e���eƪ�SEE��aSC=D��� $���PE_�_ ��!rP������.HTTPu_��HU�� (��OBJ��b(�$��fLEx3�PWq��� � ���ะ_��T?#�rS�P��z�sKRN�LgHIT܇ 5��P���P�r������PL��PSS<�ҴJ�QUERY_FL�A 1�qB_WEBwSOC���HW��1U���`6PIN'CPU���Oh��q�����d���d���� ��IHMI_ED^� T �RH�;?$��FAV� d�~Ł�IOLN
◓ 8��R���$SLiR$INoPUT_($
`���P�� ـS�LA� �����5�1��C��Bd�I�O6pF_AS7��$L%�}w%�A��\b.1�����T@HYķ����Rqh�wUOP4� `y� ґ�f�¤�������`PCC
`����#��>�QIP_ME��7� Xy�IP�`�U�_NET�9����Rĳs�)��DSaP(�Op=��BG`�����M�A��� lLp:CTAjB�pAF TI�-U��Y ޥ�0�PSݦBUY ID I�rF ��P��a��L �y0�,�����Ҥ�NQ�Y R��I�RCA�i� �k ěy0�CY�`EA�����񘼀�CC�����R�0�A�7QD�AY_���NTVA����$��5 ���gSCAd@��CL����� ���𵁛`8�Y��2e�o�N_�PACP�q��ⱶ��,� N����
�xr���:p<�N� 2��Ы��(ᵁ����xr۠L�ABy1��Y ��UN�IR��Ë ITY�듭��ed�R#�5�|��R_URL��o�$AL0 EN�Шҭ� ;�T��T_}U��ABKY_z���2DISԐ�kSJ4g����P�$���ED��g�R��З A�d/���J����FLs��7 Ȁ���
�U�JR� ��pF�{0G��E7��J�7 O R$J8BI�7��R�d�7���E�8{�H�APHI�QS��DeJ�7J8�B��L_K�E*�  �K���LM[� � �<X�XRl�u���WATCH_VA��xo@D�tvFIELc�ΘcyE ��4� �o1Vx@��-�CTh[�9�m��`LGHӿ�� $��LG_SIZ�t�z��2y�p�y�FD��I x���+!��w�\ ���� v��S���2��p��������\ ���A�0_gCM]3NzU
RAFQ\vv�d(u�"B��2�p����I��+ `�\ ��v�RS����0  �ZIPD�Uƣp�LN=��ސ�p�z6���f��>sD�PLMCDAUiEAFp���T�uGH�R.OGB�OO�a�� C��I�IT+���`揖RE���SCRX� �s��DI��SF0n�`RGIO"$D�@����T("�t|�S�s�{�W$|�X��JG=M^'MNCH;�|�FN��a&K�'uЅ)�UF�(1@�(FWDv�(HL�)STP�*�V�(%Г(��(RS"9HIP�+��C[T�#  R��&p:'^9U=q�$@9'�H%C𜓚"Gw)�0PO�7�*��#W�}$���)EX��TUI�%I���Ï���r�CO#C� *�$S���	)��B@�NOFANA|��Q
��AI|�t:��EDCAS��c�C�c�BO�HEO�GS���B�HS�H(IGN�����!�O���DDEV<7LAL�ѩ�|�­Ц(�;�T�$��2�p�������#A���(��`�{�Y��POS1
�U2�U3�Q	��2�@��Ш ��{�PtD ����&q)��0��d��VSTӐR�Y�r�B@ ` �$E.fC.k�p<p=fPf8���4�ѩ LRТ�  ��x�c�p��<�Fp�dY�@!�_ ������Kq&���c��MC7� ���CLDPӐ��TRQLI#ѽ�yt�FL��,r�5s8�D�5wS�LD5ut5u�ORG��91HrCRESERV���t���t�� �c�� � 	u95t5u��PTp��	xq�t>�vRCLMC�� �����qq�M��k�������$DEBUGMAS��ް��J?U8$T@��Ee�g��pFRQՔ߮ � j�HR/S_RU7��a��yA��k5FREQ� �$/@x�OVEAR��n��V#�P�!7EFI�%�a��pg��t���t� \RМԁd�$U�P��3?A��PS�P��	߃C��͢a��9U\�l�?(P����MISC� d�@�QRQ��	��TB � Ȗ0A՘�AX����ؗ�EXGCESj�	᫒M���\�������� �T��SC�P � H��̔_��ƘǰP]�����KHԳK��J� m�B_K�FL�IC�dB�QUI[REG3MO��O˫�3�&�ML�`MGմ �`��T����aNDU�]���>��k�G�Df��I�NAUT���RSM>�a��@N�r]3x-��p5�PSTL\�w� 4X�LOC�V�RI%��UEXɶA�NGuBu�R�ODA��������YBMFO����Y�b@p�e4�2k�SUP�ev��FX��IGG� � �A��c ���cQ6�dD�%�b|� !`��!`��|��3w�ZW�a�TI��p�q M���[�� t��MD
��I�)֟@����HݰM��DIA�����W,!�wQ�1*�D�)��O���n]�� 0�CU��VP��p��O!_V��ѻ ���S�LX�5������P��h0N���P��KES2���-$B� �����ND2����2_{TX�dXTRA�C�?�/��M�|q�`�Pv��XҰ�Pt �SBq`�USWCS��T��	���PULYS��A�NSޔ��<R��JOIN��H��~`j�=��b��b�����P=��$��b$���TA����S���hS�HS�E��SCF�baPJ��R��PLQ������LO��н�.���^����8�p������0�RR2���� 1��eA^�q d$��Iΐ�+�G�A2+/� w�PRIN��<$R SW0�"�a/�ABC�D�_J%�¡u��_Ju3�
�1SPܠ$e�u�P��3����`u��J/���r��qO8QIF��CS�KP"z{�{�J���QL2LB�Ұ_AZ�r�~E�LQ��OCMP0ೕ�T���RT������1�+���P1���>@�Z�SMG�0��=�JG�`SCyL�͵SPH_�@���%V�u� R�TER`  �< A)_�@G1"�A�@c̔�\$DI�
"23=UDF  �~ �LW�(VELqIqN�b)@� _BL�@ u��$G�q�$�'�'�%8`<�� ECHZR/��TSA_`� ���E}`<����5�B��1}`_�� �@)5D2d%��A4I��N9�t&pPDH�A�����P$V `�#>A�$��Ͳ�$�Q�R}ӆ��H �$BELv�|��<!_ACCE�!�c��7/��0IRC_4] ��pNTT��SO$PS�rL�  d�/Es��F{�@F 
��9gGCgG36B���_�Q�2�@�A��n�1_MGăDD�A]"ͲFW�`���3�E�C�2�HDE�KPP�ABN>G��SPEE�B�Q%_pB�QY��Y��11$USE_t��,`Pk�CTReT�YP�0�q P�YN���Ae�V)хQM���ѷ��@O� YA�TINCo�ڱ�B�DՒ8�WG֑ENC�����u�.A�2Ӕ+@INP�OQ�I6Be��$N�T�#�%NT23_�"�2IcLO� �2_`��I�_�if� _�k��? �` ej�C400fMOSI�A���ОA����PERCH  �c��B" �g��c�� lb=�����oU�@�@	A6B(uLeT	~��1eT�ljgv�fTRK@%�AY��"sY� �q6B�u�s۰�]��R�U�MOMq�ՒY�M!P�^��C�s�C�JR��DUF �BS_�BCKLSH_C 6B)����f���St�H���RR��QDCLAL�M-d���pm0��CH�K���GLRTY���d��Y��)�N�d_UM]�ԉC�p�A!�=PLMT� �_L�0��9��E �.� ��#E)�#H� `=��Q3po�xPC�a�xHW�頿EׅCMqCE��@�GCN_,1ND�Ζ�SF�1�iVoR��g<!��6B�n��CATގSH)� ,�DfY��f��7A����܀PAބ�R_	P݅�s_ �v���s����JG�T�]���Y�����TOR�QUaP��c�yPO�U��b��P%�_W �u�t��1D��3C��3�C�IK�IY�I�3F��6�����@VC"�00RQ�t��1���@8ӿ��ȳJRK���,��UpDB M��Up�MC� DL�1BrGRVJ�Cĭ3Cĳ3$��H_��"�j@q�CO1S~˱~�LN��� µ�ĭ0�����u��ʈ�̓��Z���f$�M�Y��؊���>�T�HET0reNK2a3�3hҧ3��CBm�kCB�3C! AS� ���u��ѭ3��m�SB8�3��x�GTS$=QC�����������$DU��Kw�B(�%(��%Qq_��a��x�{�K���b(��\�A`Չ��p�{�{��LPH~�g�Aeg�S µ��������g����(��֚�V��V��0���V��V��V��V���V	�V�V%�H���������G�����H���H��H	�H�H*%�O��O��OV	��UO��O��O��O��UO	�O�O�Fg�����	�����SPBALANCE_-ѶLE��H_`�S�P!1��A��A��PFULCElTl���.:1��UTOy_����T1T2��22N���29`�!@�qnL�=B�3�qTXp�Ov 
A4�INSE9G�2�aREV��`�aDIF�uS91�l8't"1�`OB.!t�M��w2�9`��,�?LCHWARRCBAB�� ��#�`-�(�Q 5�X�qPR��&8��2�� 
�""���1eROB͠CR�6B5�����C�1_���T � x $WEIGH�PF`$��?3àI�Q�g`IFYQ�@LAGĒRq�S�R �RBI�Lx5OD�p�`V2S�T�0V2P!t�W0P�01�&1/0�30
�Px�2�QA  2řd^[6DEBUg3L_@z�2�MMY9&E� Nz�D`$D�_A�a$�0��O� �
�DO_:@A.1� <B0�6��m�Q�B�2�0N�-cdH_p`�P�2O��� �� %"��T`"a��T/!�4�)@TICKh3| TE11@%�C ��@N͠�XC͠R?��Q�"�E��"�E8@PROMP��SE~� $I�R��Q��R;pZRMCAI)��Q�R4U_r0C2S; �q�PR8�7COD�3FU�Pd6ID_[�vU R!�G_SUFFu� �l3�Q;Q�BD�O�G �E�0�FGR r3�"�T�C�T�"�U�"��Uׁ�T8D�0�B0Hnb _FI�19*c7ORD�1 50�2�36V�+b�Q1@$�ZDT}Us0�1;E��4 *:!L_N�AmA�@�b�EDEF_I�h�b�F�d�E�2��F�4�F�c�E�e�FISP��PAKp�Ds�C�d��44בi��2�D�"�It�3D�O|#OBLOCKEz���S�O�O�Gq�R�PUM�U�b�T�c�T�e�T !r�R�s�U�c�T�d�R �6�q�S� ���U�b��U�c�S�Z��X�@P@` t�@qe�)@W�xt���s���TE��<D�( l1LOOMB_��ɇ0V2wVIS;�ITYV2�A��O�3A_FR1I��a SIq�BQR�@��@�3�3
V2W��W�4����9_e��QEAS^3�R@ϡ��_�[p:R�4��5�6_3ORMU�LA_Iz���T�HR^2 �Gtg��30f��<8�5COEFF_O�A	 ��A���GR�^3Sg0BC�AnO/C$��]3����1GRP� ?� � $�p�YBX�@TM~w���u��B�s��bCER, T�ttsd�0�  �L�L�TSpS~�_SV Nt�ߐ���0�@����0� ��SETUsMEA*P�P���W0�1+b/0� � h��  @ڐo� l�o�cqz��b�@cqq`tP�G��R�� Q\p*q[p��>�c �NPREC>at��5@MSK_$|��� PB11_USER�e"�{ ���VEL���{ 0��$Ō!I]`��MT�ACFG��� � �@@ O�"NO�RE-0l@o�V�SIb.1�d��6�"UXK��fP!��DE�� �$KEY_�3>�$JOG��0SV������!��}��SW�"�a\aS�ՐT�|�GI�!0| ^�� 4 h��'d2�!XYZc���3z� ��_ERR#�C� 8Ԡ�AfPV��d��1����$BU�F��X�����MO�R|�� HB0CU d�lA�!��GQ\aB�,"�!a$� ����a��u��?�G~�� � $SIՐ����VO��T�0O�BJE_��ADJyU)B��ELAY��4�%�DR�OU.`=ո�ВQ0b=��T����0���;BDIR����; I�"0DY�NW�#���T��"R����@�0�"�OPWwORK���,%@�SYSBUy�SCOP��ޑ�U�b; P�pN�<�PA��t�>�"��OP�PU�d!0�`!��l�IMAGw�B0y�23IM�Õ�INe�d�~��RGOVRD��-��o�Pq��0��PJ�Os���"L�pBa�|��o�PMC_Ee`���1Ny M A�211�2v���SL_���� � $OV�SL�ǫ�?q�`��2�" -�_��k�P���k�Pu���2�C�� �`�Ź���_Z�ER�D��$G�� 2=���G� @*���%O~PRI��� 
JP�8+ 1=!/�L�����T� �0ATUS>��TRC_T���sB��}fs�9s�18Re`��� DFAm�����L���"��0a� ޱ��XEw{���Ī�C0vUP��+p	qPXP�j��43 ��PG�\���$SUB�e�%�qe9JMP�WAIT z}%L�O��F�A�RCV!FBQ�@x"�!R�� �.x"ACC� R&�B��'IGNR_PL^9DBTB�0PqFy!BWbP�$w�Uy@��%IGT�PI��T'NLN�&2R��r�L�NP��PEED| \HADOW�06�w��E[q4jO!�`SPDV!� L�bAz�`�07�3UCNIr��0"!R���LYZ`� o��P�H_PK��e�RETRIE9{�q����0'PFI"��� �G`�0D 2}�g�DBGLV�#?LOGSIZ��EqKKT�!U��VDD�#�$0_T�G�MՐCݱ��|@eMRvC}�3֟CHECK0���)PO�V!�k�I��LE(!��PArpT(�2K�W��@P2V!�� h $AR@IBiR� c�a/�O�P8�ӐATT��2��IF|@z�Aq4S�3UX8����PLI2V!�� $g���ITCiHx"[�W �AS9�N2 vTLLB�V!�� $B�A�DYs��BAM�!���Y9�PJ5Ƚ�Q��R6�V�Q_KGNOW�Cb��U��#AD�XV��0D�+i?PAYLOAt��BIc_��Rg�RgZOc�L�q��PLCL_�� !7��b�Q�B��d���fF�iC�֠�js��d�I�hR�ؠ�g�ҢdB����JL��q_J�a#���AND��Ĳ.t�b�a����q�PL0AL_ �P�0���QTրC��DNcE����J3CpWv� TPPDCK������>��_ALPHgs�s�BE��gy|��K�1�� � �\��HoD_1Oj2ydD��AR�*��;��&���TIA4U�5:U�6��MOM��a����n���{�Y�B� A�Da���n���{�PUB��R��҅n�҅{�¡��2�Wp��W � � PMsbT�� BxQ���� e$PI��81�@�TgJ��niJ�IV�Id�Ir��[��3!��>!��r�Ӫ�U3HIG�SU3�%�4 얎4�%� ���"�����!
��!�%SAMP ���^��_��%�P4s ю���[ 	� ��3 ���0���&�C�@����^��Sp��H&0	�IN�SpB�����뤕"��6��6�V�GAMM�SyI�� #ETْ��;�D�tA�;
$ZpIBR!62]IT�$HIِ_��H��C�˶E��ظAҾ���LWͽ�
���@7���rЖ,0�qC�%�CHK��" �~I_A�����Rr �Rqܥ�Ǚ��ԥ��ɾWs �$�x �1���I7RC�H_D�!� RN{��#�LE��ǒ!�,��x���90MSWsFL�$�SCR((G100��R@��3]B ��ç��a����َ0���PI3A9�MET�HO����%��AX�H�XX0԰62ESRI��^�3��R�0$u	��pF{�_���I?ⲣ1�L�L�_�a�OOP����wᜲ���APP:���F����@{���أRT�V�OBp�0T����;��� 1�I��� ���r���RA�@MG�A1�B&�SV-��;P_@CURg�;��GRO[0S_SaA�Q��Y�#NO�pC!"�tY��Zo lox�������!b����&�DO�1A���A�� ��Х��A���A"�WS�c �2h�*��� � ��YL(H�qܧ��SrZ� ]B�o�@��ĵq�_�C1��M_W����g���c�M@� �`Vq�$pԐx1o�3"�PMJ�,��C �'A� 9�!Wi:�$�LWQ|ai �tg�tg�tg{t� ��N`���S��SpX�0O�sRqZ��P� �*�� ���M�� ������������X���X ��@��PL�q_~R� |�q#(Y����& n��&{�Y�Z��'�&t���Q��D�#0�� �}`�$PQ�PMO�N_QUc� �{ 8�@QCOU��n%PQTH��HO�n^0HYS:PES�RF^0UEI0O��@O|T�  �0PGõz�RUN_TO�q�0ْ.�� PE`�5C��A<�IND}E�ROGRA�nP� 2g�NE_NO�4�5IT��0�0�INFO�1� ��Q�:A�� �PO�IB� (��SLEQݖFAѕF@�6 �OSy�T� 4��@ENAB��0P�TION.S%0ER�VE���G��A0zCG�CF�A� @R0JX$Rq�2���R�H��O�G "�EDI�T�1� �v�K��ޓʱE�NU�0W*XAUTu�-UCOPY�ِN\�����MѱNXP\[q�PR�UT9� _RN�@O;UC�$G�2�T>���$$CL`��O����Qa�a� �P�S�@�X��PXK�QIGRTU��_�PA� _WRK 2 e��@ 0 � �5�QMoYh\Jo|m |l	�`�m�oa�`��o�o�f�e�l}�aI�[ct'`BS�*� �1�Y� <7����� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P��b�t���������srC�C��LMT�P����s  dѴIN�ڿ�дPRE_EXE��)�Ƅ0jP���za'`DV��S��@e)�%s�elect_macro����kϤ�qt�IOCNVVB�� 5��P��USňw����0V 14kP $$p��a�|�`?��Ɛ >�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ ���$�ѰLARMRE?COV ^������LMDG ��Ь�LM_�IF ��d�  YST-32�3 Collab�orative �speed li�mit (TCP) ) e����� �8�J�\�n��?, 
 ����#�8TELEOP� ǘLINE 6�ǑAUTO RU�NNINGǘJO�INT 100 1%�����$���1�@�$�@���ROG-057 �Power Fa�il Recov���memory �is clear�쏹�˯��NGTO�L  @� 	 A   ��Ѱ�PPINFO �� f�L�^�p����  ������ k���ۿſ�����5���Y�C�iϏ�%��� ٯ����������'߀9�K�]�o߁ߓߙ�P�PLICATIO�N ?t���|�Ha�ndlingTo�olǖ 
V9.40P/17����
88340�����F0�	�54�9��������7D�F5�О�ǓNon}e��FRA��� ؒ��,�_A�CTIVE1�  ��� �  ��ސM�OD��������CHGAPONL��� �OUPLE�D 1	��� �>�B�T�f���CUR�EQ 1
��  UTp�p�p�	�� ������l��������������i3l�;p���^�H��A�t
HTTHKY�FXv |��*<N `������� �//&/8/J/\/�/ �/�/�/�/�/�/�/�/ ?"?4?F?X?�?|?�? �?�?�?�?�?�?OO 0OBOTO�OxO�O�O�O �O�O�O�O__,_>_ P_�_t_�_�_�_�_�_ �_�_oo(o:oLo�o po�o�o�o�o�o�o�o  $6H�l~ ��������  �2�D���h�z����� ��ԏ���
��.� @���d�v���������Ƃ�TO�����DO?_CLEAN���E�NM  �� p�������ɯۯ�v�DSPDRYRLL���HI��o�@�� G�Y�k�}�������ſ�׿����ϻ�MA�X��,�����=�X�,�<�9�<���PLU�GG,�-�9���PRUC��Bm�q�6��(ϗ�O����SEGF�K���� �m� �G�Y�k�}ߏ�����LAP$�7ޡ���� ��+�=�O�a�s������ �TOTA�L_ƈ� �USENU$�1� �������RGDISPM+MC�d�C�O��@@�1�O"�D���-�_STRIN�G 1��
��M��S��
~��_ITEM1��  n���������  $6HZl~ ��������I/O SI�GNAL��T�ryout Mo{de��InpN�Simulate�d��Out`�OVERR!� �= 100��I?n cyclT���Prog Ab�orj��JSt�atus��	Heartbeat���MH Faul<��Aler�! /!/3/E/W/i/{/�/�/�/ (���(� ���/??&?8?J?\? n?�?�?�?�?�?�?�?��?O"O4OFO�/WORИ�~A�/XO�O�O �O�O�O __$_6_H_ Z_l_~_�_�_�_�_�_�_�^PO���"` �KoEoWoio{o�o�o �o�o�o�o�o/�ASew��bDEV%n�p9o��� �#�5�G�Y�k�}��� ����ŏ׏�����|1�C�PALT�- j��OD�������ȟڟ ����"�4�F�X�j��|�������į֯X�GRIB�������6� H�Z�l�~�������ƿ ؿ���� �2�D�V�h�z�����R�-��&� ���������"�4�F� X�j�|ߎߠ߲�������������PREGn�W���0�~��� ����������� �2� D�V�h�z���������~$�$ARG_~@�D ?	����� � 	$$	[]�$:	���SBN_CONF�IG�XW�qRCII_SAVE  $zm���TCELLSE�TUP 
%�  OME_IO�$$%MOV_qH� ��REP���#��UTOBAC�K� 	t�FRA:\D� �.D�z '`��D�w� �s � 25/1�1/29 20:_26:16D�;�D���#//h�� C/j/|/�/�/�/�/D��X/�/??(?:?L? �/p?�?�?�?�?�?�? g? OO$O6OHOZO�? ~O�O�O�O�O�O�O��ׁ  c_F_\�ATBCKCTL.TM�)_;_M___\q_8INIm���j~CMESSA�G� �Qz �[ODGE_D� �j�X�O�p�_@PAUS�6` !� , 	�; :oHg,		2oloVo �ozo�o�o�o�o�o�o  
D.Pz}d`?TSK  mw<}_CUPDT�P�W�d�p�VXWZD�_ENB�Tf
�vS�TA�U�u��XI}SX UNT 2�v�wy � 	�p/�� ��L��g��^�? :L�D�R��  �� ������Ut���D�R�.��1o���[ #g ?o� ��y���p���,�/�MET���2@��y PQ�A�##,@���A�{�@��A#�AmbM��>z��>%;�>$�H<�ԡ�?��>}���5�SCRDCFG� 1Y ��w���@�%�7�I�pD�Q�	 ܟ������ϯ��Z� �~�;�M�_�q�����0��6���FGR9��pX�_ԳPNA� s	FѶ_ED�P�1��� 
 ��%-PEDT-`¿ R�v���Es�� -FE�D�;�9/�>���  ����2�����B� ��ˀ�{�����j�����3 ��#� �G�Y���G����6�����4����� �Yި��Z�l������5K������Y�t�@��&�8���\���6 ��d��Y�@����(��7�S0w Y�w��f���!8�W��{�IZ��@C/��2/���9{/��//LZݤ/?V/0h/�/�/��CR�� �?�?Tn?�? ?2?�?�V?԰!�NO_DE�L�ҲGE_UN�USE޿дIGALLOW 1��   (*SYSTEM*
��	$SERV_�GR[�@`REGƜE$�C
��@NU�M�J�C�MPMU|?@
�LAYK��
�PMPA�L�PUCYC10� N3^P!^YSUL�SU_�M5Ra�C�Lo_�TBOXOR=I�ECUR_�P�M�PMCNVV��P10I^�PT4�DLI�p�_�I	*�PROGRA�D?PG_MI!^KoF]`AL+ejoTe]`�B�o�N$FLU?I_RESU9W�o�O�o�dMR�N�@�<�?�;M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3��E�W�2BLAL_OUT �K���WD_ABOR:P�cO��ITR_RT/N  �$�빸�?NONSTO��� lHCCFS_UTIL ��̷CC_AUXA�XIS 3$� h}�j�|�����ƽ�CE_RIA_IL`@�נ��FCFG $��/�#��_LIMv�B2+� �8p7� 	��B\���$�8p
Ԡ��)�Z��%�/�����[����� ���!�����L��(
5������PA�`GP 1H�����A�SϨe�w�6�CC� CU7��J��]��p��}����� C���U������������Ué�̩�ձ�ߩ�U�������;����PCk���������������������Ա��������� D� D!��!�!�!� ���&?��HE@O�NFIpC�G_�P�P1H�  +EH��ߟ߱�����������C�KPAUSf�Q1H�ף IR �S�H�A��e��� ������������E��+�i�{�a���A�?Iץ�MؐNFO� 1���� �3��$4��Q�*sB|Ӷ¬�|,A�V/���A��~��'����ײ�&���úמ�3��@����|�hPb�O� �� ��LLECT_��!�����EN�+`�ʒ���NDEַ#�/��1234567890�"�A��/ҵHw��#)j��< i{��;��/� �/`/+/=/O/�/s/ �/�/�/�/�/�/8?? ?'?�?K?]?o?�?�?@�?�?O�?��$�� ��IO #&��"S▒O��O�O�O`GTR�2'DM(��^�?�NN��(oM Z��_M[OR)q3)H��7� �U3��Y�_�_�_�_�_P�[bR�kQ*H�,S�I?<�<Ѡ<c8pKFd����P,�� ;ϒo�o�o˿�o�oœh�UY@E�oS� �sja.�PDB.���4�cpmidbg03��Рs:��>uq�pz��v  E��>x��}.���}�`��|�<�m!gP���t��~f��������@ud1:��?��XqDEF �-��zC)*�c�O�buf.txt�J��|K�[`�/DM��>���R�A���MCiR20_{RCdX���hS21������CzA�d4�EI��jA��]A����F]� B��e;t�H�j��C1�aCN/��I؂�DH�����LڒYE��E�>�MS?o�F��&ġ���>��&N��f2�3DLD�	>	P!�� 2��}��yc
f�@x9� C�ğ�  D4G�E����  E%q��F�� E�p��u�F�P E���fF3H ��GM�����?5�>�33H��?�xn9�q@�QG5����RpA?a���=L��<#�QU�@,�Cϒ����RSMOFST �+i�����P_Tu1Ɠ4DMA =����MODE 5�dm�@��	Q�M;��%��?����<�M>�̽Ͷ�TESTc�2i�`�R�6�O�K�ECN�AB���n� 8���\�n�CdB�f��Cpp�����	P:d�QS ���� ������4�IJ7>���>B8m�5$�RT_c�P�ROG %j%�d�1�h@NUSE�R��x�KEY_T�BL  e������	
��� !"#$%&'�()*+,-./�(:;<=>?@�ABCc�GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������>��͓���������������������������������耇���������������������9�4A8�LCK��F�<y��STAT��2�=X�_ALM������_AUTO_D�O�E�FDRw 3:i�2hi�AUS�x��i�$g ��A����� �T*g�2�  bf��/�/9/ ;�*pm�P/z/�~/h/ �/�/�/�/�/?"=� G?Y?k?/|?�?L/�? �?�/�?�?OO�?*O @OvO�O6?�O�O�O~? �O	_�?*_$_BOD_6_ p_~_T_�_�_�_�_�O o)o;o�OLoqo_�o �o�_�o�o�o�o�o�o FXo��No ���o���� @�N�$�b�x�����n ������A��b� \�z�|�n�������ʟ ���(�֏O�a�s�� ����T�ʯį��֯ ����2�H�~���>� ��ɿۿ���ϼ�2� ,�J�L�>�xφ�\Ϛ� �����Ϧ��1�C�� T�y�$Ϛߔ߲ϴߦ� ��������N�`�� ����V߼����� �����H�V�,�j� ������v����� $I��jd���v �����0�� Wi{&��\� ����/&/�:/ P/�/�/F�/�/�/� �/?�:?4?R/T?F? �?�?d?�?�?�? O�/ 'O9OKO�/\O�O,?�O �O�?�O�O�O�O�O
_  _V_h_O�_�_�_^O �_�_�O
oo"_$oo Po^o4oro�o�o�o~_ �o	�_,Q�_r l�o�~���� �&�8��o_�q���. ����dڏԏ���  �.��B�X�����N� ǟٟ럖���!�̏B� <�Z�\�N�����l��� �������/�A�S��� d���4�����¯Ŀ�� ���Կ�(�^�p�� �ϩϻ�f����Ϝ�� �*�,��X�f�<�z� �����߆����#��� 4�Y��z�t�ߔ�� ���������.�@��� g�y���6����l��� ��������(6J `��V������ )��JDbdV ��t���/� 7/I/[/l/�/<�/ �/��/�/�/?�/? 0?f?x?&/�?�?�?n/ �?�?�/OO2?4O&O `OnODO�O�O�O�O�? __+_�?<_a_O�_ |_�O�_�_�_�_�_�_  o6oHo�Ooo�o�o>_ �o�ot_�o�oo�o 0>Rh��^o ����o�1��oR� L�jl�^�����|��� Џ���?�Q�c�� t���D�����ҏԟƟ  ���"�8�n���.� ����˯v�ܯ���"� �:�<�.�h�v�L��� ��ֿ迖��!�3�ޯ D�i���τϢ��ϖ� ���ϴ����>�P��� w߉ߛ�FϬ���|��� ��
����8�F��Z� p���f�������� �9���Z�T�r�t�f� ���������� �� GYk�|�L�� ������* @v�6���~ �	/�*/$/BD/6/ p/~/T/�/�/�/�/� ?)?;?�L?q?/�? �?�/�?�?�?�?�?�? OFOXO?O�O�ON? �O�O�?�O�OO__ @_N_$_b_x_�_�_nO �_�_o�OoAo�Obo \oz_|ono�o�o�o�o �o(�_Oaso ��To���o�� ���2�H�~���> ��ɏۏ����2� ,�J�L�>�x���\��� ��������1�C�� T�y�$����������� ��į��N�`�� ������V���ῌ�� �����H�V�,�j� �϶���v����߾� $�I���j�d߂τ�v� �߾ߔ������0��� W�i�{�&ߌ��\��� ���������&���:� P�����F�������� ����:4R�TF ��d��� �� '9K��\�,� �������
/  /V/h/�/�/�/^ �/�/�
??"/$?? P?^?4?r?�?�?�?~/ �?	OO�/,OQO�/rO lO�?�O~O�O�O�O�O �O&_8_�?__q_�_.O �_�_dO�_�_�O�_�_� o.ooBoXo�otc��$CR_FDR_�CFG ;re��Q
U�D1:�W�TJ�d � �`�\�bHISoT 3<rf  �`  ?�RW@tAtBtUC�PpDtEt�Itg�Pqotw��_��bINDT_�EN6p�T��q�bT1_DO  �U�u�s�T2��wVAR �2=�gp h�q  y�������R��TF4��T�m[��RZ�`�STOP��rTRL_DELETNp��t ��_SCR?EEN re�r�kcsc�rU�w�MMENU 1�>��Ap<�\% �_��T��R��S/� U���e�w�ğ������ џ�	�B��+�x�O� a�����������ͯ߯ ,���b�9�K�q��� ����࿷�ɿ���� %�^�5�Gϔ�k�}��� �ϳ��������H�� 1�~�U�gߍ��ߝ߯� ������2�	��A�z� Q�c��������� ��.���d�;�M��� q������������Y�Ӄ_MANUAL�{��rZCD�a?x�y�rG ���R��f"
�"
?|�(��PdTGRP� 2@�y�B1� � s��� ��$DBCO�pR�IG���v�G_E�RRLOG A���Q�I[m ��NUMLIM��s��u
�PXWORK 1B�8���//�}�DBTB_�� !C%���S"� ��aDB_AWAYz��QGCP �r�=�ןm"_AL(�F�_�Yz���p�p�vk  1D� , 
��/"�/%?/(_M�pqw,�@�=5ONTIM6����t�_6�)�
�0�'MOTN�ENFpF�;REC�ORD 2J�� �-?�SG�O� �1�?"x"!O3OEOWO �8_O�O�?�OO�O�O �O�O�O(_�OL_�Op_ �_�_�_A_�_9_�_]_ o$o6oHo�_lo�_�o �_�o�o�o�oYo}o 2�oVhz��o� �C�
��.�� R��K��������Џ ?��ߏ�*�����+� b�t�㏘�����Ο=� O�����:�%���p� ߟ񟦯��O�ǯ�]� �����H�Z����� ����#�5����ϩ��i"TOLEREN�Cv$Bȿ"� L���� CSS_CC�SCB 2K�\0"?"{ϰϟ� ��7��
����@�R� d�3߈ߚ�"�x��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy���� �������R�LL]�La��m1T#2 C��C��F�^ +A�C�pC���#�0�� 	 A����B���?�  �$�����\0袰�0��B� �`#s�K/]/o/�ϓ/�/�/s/�/�/��LڮL��|C�++@I���ǒ1Ȧ���.?��/`?;
�@��O?�?�?�?�Ȏ0AF��?{F�A OO�7�1���9M	AB
AZOdBAE�9�$O�O�O�Oi:P��`^�@0�DJCA�� @��
�X-._] M?�> O�ڴ�q_�_�_�_:W�A<o:[<��/o�/�_+oPobo�to�eACHC�V�ZWB$�Dz�cD�` �a=/�o�oo�oW�a.+!��2=t,y�D�p�Yrm�U I?�-t�s�js�w�y j�������Q���@`��$��� ��A����Bމ�o� �'�9��_]�o�N��� r���ɟ۟&_�B�ʄ���YZ>`�?��B�BX@�{�>�ZR��Y9�D��Z�l�~����`_м¯� ��
���̯9�,�]�o� �� �H�����ٿ뿊� �ƿ3�E�W�iϬ��� $ϱ����� Ϟ���� /�A�S߶�w�V�h߭�`���S���ߐ�_ �f	��H�?�Q�~�u� ����������� �D��-�g�q����� ��������
@ 7Icm��߾�  �����) M@qdv�� �����//I/ P�m/�v/�/�/�/�/ �/�/�/?3?*?<?i? `?r?�?^/�?�?�?�? �?O/O&O8OJO\O�O��O�O�O�O�O�O�g	o  Q�PՄs �PC4p*p�p6U6P�\C9p/p��� ]V^PM]�6P�b:P�>P�VJ_�^P��bP�fP�Vr]v�	�Tp Q
k���_o�o�id1Q&oNo �;o_co�oˏUUA �  �o�k1Q@� � �o�k�b�����Up �� 1���6��1C���C��cPfL��?#�c>_�{���`�cP��@@�d��r�`Be�cP>�s�qC��p癙��b�t<��o?�PH�)S�B�tq�q�p�r��`B���eIC��&�Q�4( �oz�UU��mO���@F@��yl>�X���9��Q��-R�� �f���#��C%��c��`ځ`  �?�p���U�[?����}t��$���$�DCSS_CLL�B2 2M���p�P�^?�NS�TCY 2N����   �������ʟ؟��� � �2�D�Z�h�z��������¯ԯ��SA�D�EVICE 2O��!�$��4&V� h�������˿¿Կ� ��
�7�.�[�R�ϑ���ϵ�����4(A�HN?DGD P��*��Cz�A�LS 2Q��_�Q�c�u߇���߽߫���?�PARAM RP��1��`�&�RBT 2T��� 8�P<C�'p �qi�l��s@"�R��(qI�ʹX��0�pB CW  ��B\x�N��`�Z����%��)� ��X�j��p����zq��I���B �(s,�F� �p�V��q���b��B ��4&c �S�e� l�4+����H1~ޡ���D�C��$Z��b���A�,� 4�u@�X�@��^@w����]B���B��cP%��C4��C3:^C4��nЬ ��p8�-�B{B���A���� l���C�C3��JC4jC3���yn+�3 Dff 2�A PB W4+@:�]o�W �����/�/ P/'/9/K/]/o/�/�/ �/�/?�/�/�/?#? 5?�?Y?k?�?�?�o�? �?O�?6O!OZOlOWO �O�Es�?�?�?�O�O _�O�OL_#_5_G_Y_ k_}_�_�_�_ o�_�_ �_oo1o~oUogo�o �o�o�o�owO D /Aze����O �o�o
��o��R�)� ;���_�q��������� �ݏ�<��%�r�I� [�m��������ǟٟ &�8��\�G���k��� ����گů����� F��/�A�S�e�w�Ŀ ������ѿ����� +�x�O�aϮυϗϩ� ������,���b�t� ﯘ߃߼ߧ������ ���:��C�U߂�Y� k����������� 6���l�C�U�g�y� ���������� ��	 -?Q���� ���@+d vQ������ ��*///%/r/I/ [/�//�/�/�/�/�/ &?�/?\?3?E?�?i? {?�?�?U�?�?"O4O OXOCO|OgO�O{� �?�O�?�O�O0___ f_=_O_a_s_�_�_�_ �_�_o�_oo'o9o Ko�ooo�o�o�o�o�o �O:%^I�������H�$D�CSS_SLAV�E U����	���z_�4D  	��A�R_MENU V	� �j�|�������ď�BY�� ��~�?�SHOW 2W>	� � �b�a G�Q�X�v��������� П֏���� @�:� d�a�s���������� ߯��*�$�N�K�]� o�������̯ɿۿ� ��8�5�G�Y�k�}� �϶�����������"� �1�C�U�g�yߠϝ� ���������	��-� ?�Q�c��s����� ��������)�;�M� t�������������� ��%7Ip�m ���������� !3ZWi�� �J����// DA/S/e/��/��/ �/�/�/�/?./+?=? O?v/p?�/�?�?�?�? �?�??O'O9O`?ZO �?�O�O�O�O�O�OO �O_#_JOD_nOk_}_ �_�_�_�_�O�_�_o 4_.oX_Uogoyo�o�o �o�_�o�o�ooBo ?Qcu���o:����CFG MX)�3�3q5p��FRA:\�!�L+�%04d.WCSV|	p}�� �qA g�CHo�zv�	����3q�����́܏� �|��4��JP�����qp1� �R�C_OUT Y���C��_�C_FSI ?~i� .� ������͟����� >�9�K�]��������� ίɯۯ���#�5� ^�Y�k�}�������ſ �����6�1�C�U� ~�yϋϝ��������� �	��-�V�Q�c�u� �ߙ߽߫�������� .�)�;�M�v�q��� ����������%� N�I�[�m��������� ��������&!3E ni{����� ��FASe �������� //+/=/f/a/s/�/ �/�/�/�/�/�/?? >?9?K?]?�?�?�?�? �?�?�?�?OO#O5O ^OYOkO}O�O�O�O�O �O�O�O_6_1_C_U_ ~_y_�_�_�_�_�_�_ o	oo-oVoQocouo �o�o�o�o�o�o�o .);Mvq�� �������%� N�I�[�m��������� ޏُ���&�!�3�E� n�i�{�������ß՟ ������F�A�S�e� ��������֯ѯ��� ��+�=�f�a�s��� ������Ϳ����� >�9�K�]φρϓϥ� ����������#�5� ^�Y�k�}ߦߡ߳��� �������6�1�C�U� ~�y����������� �	��-�V�Q�c�u� �������������� .);Mvq�� ����% NI[m���� ����&/!/3/E/ n/i/{/�/�/�/�/�/��/�/3�$DCS�_C_FSO ?����71 P ? ?T?}?x?�?�?�?�? �?�?OOO,OUOPO bOtO�O�O�O�O�O�O �O_-_(_:_L_u_p_ �_�_�_�_�_�_o o o$oMoHoZolo�o�o �o�o�o�o�o�o%  2Dmhz��� ����
��E�@� R�d���������ՏЏ ����*�<�e�`� r���������̟��� ��=�8�J�\�����|��?C_RPI4>F?�������3?��&�o����� >SLү@d������%� 7�`�[�m�Ϩϣϵ� ���������8�3�E� W߀�{ߍߟ������� �����/�X�S�e� w����������� �0�+�=�O�x�s��� ���������� 'PK]o��� �����(#5 Gpk}����� Q���/6/1/C/U/ ~/y/�/�/�/�/�/�/ ?	??-?V?Q?c?u? �?�?�?�?�?�?�?O .O)O;OMOvOqO�O�O �O�O�O�O___%_ N_I_[_m_�_�_�_�_ �_�_�_�_&o!o3oEo noio{o�o�o�o�o�o �o�oFASe�������>�N�OCODE Z�U��?�P�RE_CHK �\U��pA �p?�< ��pU�x]�o�U� 	 <Q� �������ۏ�Ǐ� #����Y�k�E����� {�şן��ß���� C�U�/�y�����s��� ӯm���	���?�� +�u���a�������ɿ �Ϳ߿)�;��_�q� K�}ϧϝ������ω� ��%����[�m�Gߑ� ��}߯��߳����!� ��E�W�1�c��g�y� ������������A� S�-�w���c������� ������+=a sM_����� �'�]o	 ������/ #/�G/Y/3/e/�/i/ {/�/�/�/�/?�/? C?9Ky?�?%?�?�? �?�?�?	O�?-O?OO KOuOOOaO�O�O�O�O �O�O�O)_____q_ K_�_�_a?�_�_�_�_ o%o�_Io[o5oGo�o �o}o�o�o�o�o�o �oEW1{�g� ��_����/�A� �M�w�Q�c������� ���Ϗ�+���a� s�M���������ߟ� ��'���3�]�7�I� �����ɯۯ���� ���G�Y�3�}���i� ��ſ��������1� C���+�yϋ�eϯ��� ����������-�?�� c�u�Oߙ߫߅ߗ��� �����)��M�_�U� G���A�������� �����I�[�5���� k������������� 3EQ{q�� �]����/A ewQ���� ���/+//7/a/ ;/M/�/�/�/�/�/� �/?'??K?]?7?�? �?m??�?�?�?�?O �?5OGO!O3O}O�OiO �O�O�O�O�O�/�O1_ C_�Og_y_S_�_�_�_ �_�_�_�_o-oo9o co=oOo�o�o�o�o�o �o�o__M_�o k�o����� ���I�#�5���� k���Ǐ��ӏ��׏� 3�E��i�{�5c��� ß�����ӟ�/�	� �e�w�Q�������ѯ 㯽�ϯ�+��O�a� ;��������Ϳ߿y� ���!�K�%�7ρ� ��mϷ��ϣ������� ��5�G�!�k�}�W߉� �ߩ������ߕ��1� ��g�y�S���� ��������-��Q� c�=�o���s������� ������M_9 ��o���� �7I#mY k������!/ 3/)/i/{//�/�/ �/�/�/�/�/?/?	? S?e???q?�?u?�?�? �?�?OO�?%OOOE/ W/�O�O1O�O�O�O�O __�O9_K_%_W_�_ [_m_�_�_�_�_�_�_ o5oo!oko}oWo�o �omO�o�o�o�o1 UgAS��� ���	����Q� c�=�����s���Ϗ�o ������;�M�'�Y� ��]�o���˟���� ۟�7��#�m��Y� �����������!� 3�ͯ?�i�C�U����� ��տ�������	� S�e�?ωϛ�uϧ����Ͻ������$�DCS_SGN �]	�E��-����30-N�OV-25 16�:44 ��2}9R�20:27_��x�x� [}�t��q�т�xҚ����JѨ�EƼÿ�� ��ǖ� � 1�HOW ^�	� �x�/�VERSIO�N =�V�4.5.2��EF�LOGIC 1_~���  	������C��R�%�PR�OG_ENB  ���:�{�s�UL�SE  X���%�_ACCLIM^�����d��WRSTJNT��vE��-�EMO|��zя�$���INIT� `2����O�PT_SL ?	�	�	�
 	Rg575��]�74b��6c�7c�50��1����C���@�TO�  L��� �V.�DEX��dE�x��PATH A=�A\k}���HCP_CLN�TID ?�:�� D�ռ��I�AG_GRP 2�e	�����z�	 @�  �
ff?aG�x��B�  2Ě�/�8[I@c��ς!�7@��z�@^�@
��!��mp2�m15 8901?234567�����  ?����?�=q?���
?޸R?��Q�?��?������(�?��z���x�@�  A_�Ap !7�A�88_�B4��� ��L�x�
��@�@���\@~�R@xQ��@q�@j��H@c�
@\���@U�@Mp��//'$�; ��O)H��@Ct >�d 9��@4�/�\)@)� #t ?{@��/�/�/�/�/P'?����?���_ ?}�p�?u?n�{?s ?\�Q�? ?2?D?V?h8_�
=?����0�w5�z�H?p��h��?^�R��?�?�?�?�?h8��*t0���@�?��0�;@&O8O JO\OnOP'�$_�_ Y_k_�O?_�_�_�_�_ �_s_�_�_1oCo!ogo yoo�o��Bj"� �2x{1�@"?���f�t0�d"5!�
u4V��u"�BP3t�A>u��?@[q���@`,=q��=b��=�E1�>�J�>�n��>��H"<�o� �z�s�q��� �x�C�@<(�]Uz� 4�� Z����A@x�?* �o��m*�P�b���t n���2���Ώ����ޮi>J��&�byN2�"��G�N�R�o@�@v���0��^��@ffr!l Ο�33���(���"C�� ƒI��CH�)C.?dBت"8"����'���"~�A�?�&"K����pf�B��@�p�������p���?A��g����4���ٽ����	`Ơ	�9�WS�A�C�ײ�&��úםxО������3��N�T������3�@�����| �<E�q"����ǿ����ֿ���ú_���x�:���9�σǺG��!�o��C�T_CONFIG� f��|��egY��ST�BF_TTS��
@����О�}���1��MAU������MS�W_CF��g� � # ��OCVIE�W��h!�-�� �s߅ߗߩ߻��ߟ� a�����,�>�P��� t�������]��� ��(�:�L�^���� ����������k�  $6HZ��~�� ����y 2 DVh�����X��v�RC�i���!�0./S/B/w/�f/�/�/�/��SBL�_FAULT �j*6��!GPMS�K���'��TDIAOG k��-�������UD1�: 6789012345I2��=1���%P\υ?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�Od696�I�r�
t?�O|�TREC	P"?4:
B44_[7M[ s?p_�_�_�_�_�_�_ �_ oo$o6oHoZolo�~o�o�O�O�O�o7�U�MP_OPTIO2=��.�aTR���:�)uPME���Y_TEMP  �È�3BC�rgp�B�QtUNI�����gq�YN_BR�K lL�7�EDITOR�a�a@�r�_
PENT 1m�)  ,&?TELEOP^P �z��pPSNA��:�&MTPG��p+�=��/����� z�����ۏ���� 5��Y�k�R���v��� ş���П����C� *�g�N�v�������������ޯ��?�Q����EMGDI_S�TAzuV�gq�uNC�_INFO 1n<!��b���X����������n�1o!� C��o����
�d�oU�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫���  u����
��*�B�*� P�b�t������� ������(�:�L�^� p���������2����� ��9�CUgy �������	 -?Qcu�� ������//1 ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?��? �?�?O)/OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�?�?�_�_o�_ 3O=oOoaoso�o�o�o �o�o�o�o'9 K]o����_�_ ����+o5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� �������ӟ���	� #�-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ����7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߹��������� �%�/�A�S�e�w�� ������������ +�=�O�a�s������� ���������'9 K]o����� ���#5GY k}�	����� �/1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? ��?�?�?�?/O)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�?�_�_�_ �_O�_!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �_�_����o� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o�������ɟ ۟���#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߝ��߹� ���������%�7�I� [�m��������� �����!�3�E�W�i� {��߇���������� /ASew� ������ +=Oas����� �����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?���?�?�?�?� �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�?�_ �_�_�_�?�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m�_u����_ ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�� ������u������ +�=�O�a�s������� ��ͯ߯���'�9� K�]�w���������ɿ �����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g߁� �ߝ߯���ۿ����	� �-�?�Q�c�u��� �����������)� ;�M�_�y߃������� ������%7I [m����� ��!3EWq� c��������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?i{�?�?�? �?��?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_�? s?}_�_�_�_�?�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qk_u�� ��_�����)� ;�M�_�q��������� ˏݏ���%�7�I� cQ���������ٟ ����!�3�E�W�i� {�������ïկ������/�A�[� �$�ENETMODE� 1p��_�  k�k��f�����j�OAT�CFG q�����Ѵ��C����DATA 1�rw�Ӱ���*	�*��'�9�K�]�"l�dlύ�e��� ����������'ߡ� ��]�o߁ߓߥ߷�1� ��U����#�5�G�Y� ���ߏ��������� ��u��1�C�U�g�y� �����)�������	 -����cu�����j�RPOS/T_LO��t�[�
׶#5Gi�R�ROR_PR� �%w�%L�XTA�BLE  w��ȟ����RSE�V_NUM ��?  ���  ��_AUTO_ENB  ���Xw_NO5! uw����"  *�*x �x �x �x + �+w �/�/�/Q$FLsTR=/O&HIS#�]�J+_ALM �1vw� �[x,e�+�/Q?c?u?��?�?�?�/_"W   w�v!���:j��TCP_VER �!w�!x�?$E{XT� _REQ�&s�H)BCSIZKO�=DSTKhIf%��?BTOL  �]Dz�"�A =D_BWD�0�@�&��A���CDI�A �wķ���]�KST�EP�O�Oj�POP�_DO�Oh�FDR_GRP 1xw��!d 	�?�_��yP�s�Y�Q'��M"���l���T� �����VyS�_�]yPA��41B�o�A��҃A��AH?��A�d��]]�B
�A8��o@���]A=
o �_Uo@oyodo�o�o�o��o  @�7>��Ơ?�ք<��>@R\�j
 M,� a�a,bfF��o(2�o �oZE~�]@.`�tO@S33�u�]@�q��g��yPF@� ��|yPG�  �@�Fg�fC�8yRL��]?�  h���6�X����8�75t��5��ߛ5`+��]�����o������� }���㿴n�ũh�F�EATURE �y���@���Handling�Tool �]�English� Diction�ary�4D S�t��ard��A�nalog I/�O>�G�gle S�hiftZ�uto� Softwar�e Update��matic B�ackup���g�round Ed�it ��Came�raU�FY�Cnr�RndIm���o�mmon cal�ib UI��n�ˑ�Monito�r$�tr�Rel�iabn��DHC�P �[�ata A�cquis3�\�iagnos��R�v��isplayΑL�icensZ�`�o�cument V�iewe?�^�ua�l Check ?Safety��?hanced����s�Frܐ�xt. DIO /�sfi��@�end�Err>�L��\�4�%s[�rP�K� �@
��FCTN Men�u��vZ���TP ;In��facĵ��GigE־�Đp� Mask Ex�c�g=�HT԰Proxy Sv���igh-Spe�Ski�� Ť�O��mmunic��onsV�ur����q��V�ײconnecwt 2��ncrְ�stru!��ʴ�e�ۡ��J��X�KAR�EL Cmd. �L�ua���Ru�n-Ti<�Env��Ȟ�el +��s��S/W�ƥ����r�Book(Sy�stem)
�MA�CROs,M�/OOffseu�p�HO���o�u�MR8�4����MechStop"+�t����p�im�q����x�R�����od>o�witch���.��4�Optm8F��,�fil䬳��g��p�ulti-�T�Γ�PCM 'fun�Ǽ�o���������Regie�r,q���riݠF����S�Num Sel���/�:� Adju�a�*�W�q�h�tat�u��ߪ�RDM� Robot�s�cove'���ea���<�Freq Awnlyq�Rem���O�n5�����Ser�voO�!��SNPgX b-�v�SN԰�Cliܡ?r�Li#br&�_�� ��q �+oJ�t��ssag��X�@ ����	��@/Iս�MIL�IB��P Fi�rm���P��AcycŐ͛TPTXk��eln���������orquo�i�mula=��|u(�Pa&��ĐX�B�&+�ev.���r�i��TUSB �port �iP�f�aݠ&R EV�NT� nexcept�����%5��VC�rl�c��؁V���"�%q�+S�R SCN�/SGE��/�%UI	�Web Pl��>��A4�3��ۡ��ZDT �Applj�
�{1EOAT����&0?�7Grid�񾡬=.�?iR�".5� F����/גRX-10�iA/L�?Ala�rm Cause�/��ed(�All Smooth5�<��C�scii+�V��Load䠌JUp9l�@w�toS ���rityAvoi+dM(�s7�t�@�ycn������_�CS+���. c��XJo���-T3_�H�.RX��U���Xc?ollabo�����RA�:�.9D��iqn���NRTHI�
�On��e Hel����ֿ�����1�trU�ROS Eth$��A������;�,�G �B�,|HUapV�%�W�t ԰��_iRS�ݐ�64MB DRAM�o�cFRO���L8F� FlD�����2M L�A:�opm�ԕex@�V�
�sh�q��wc�e�u��p��|ty"n�sA�
�%�r����J��^�.v� P)Q/sbS�`���O�N��mai��U����R�q�T1�^FC+Ԍ%̋Fs9�ˌk�̋��Typ߽FC�%�hױV�N Sp�F�orްK��Ԭ�lu�!����cp�PG j��֡�RJ�[L`Sup"}��֐f��3crFP��lu� ��#al�����r��i��
q�4@а�ue�st,IMPLE ׀6*|HZ���c0�BTea(�|����$rtu���V�9H�MI�¤��UIFNc�pono2D�B C�:�L�y�p������� ��ʿܿ	� ��?�6� H�u�l�~ϫϢϴ��� ������;�2�D�q� h�zߧߞ߰������ ��
�7�.�@�m�d�v� ������������ 3�*�<�i�`�r����� ����������/& 8e\n���� ����+"4a Xj������ ��'//0/]/T/f/ �/�/�/�/�/�/�/�/ #??,?Y?P?b?�?�? �?�?�?�?�?�?OO (OUOLO^O�O�O�O�O �O�O�O�O__$_Q_ H_Z_�_~_�_�_�_�_ �_�_oo oMoDoVo �ozo�o�o�o�o�o�o 
I@Rv �������� �E�<�N�{�r����� ��Տ̏ޏ���A� 8�J�w�n�������џ ȟڟ����=�4�F� s�j�|�����ͯį֯ ����9�0�B�o�f� x�����ɿ��ҿ���� �5�,�>�k�b�tφ� ���ϼ��������1� (�:�g�^�p߂ߔ��� �������� �-�$�6� c�Z�l�~������ ������)� �2�_�V� h�z������������� ��%.[Rdv �������! *WN`r�� �����//&/ S/J/\/n/�/�/�/�/ �/�/�/??"?O?F? X?j?|?�?�?�?�?�? �?OOOKOBOTOfO xO�O�O�O�O�O�O_ __G_>_P_b_t_�_ �_�_�_�_�_ooo Co:oLo^opo�o�o�o �o�o�o	 ?6 HZl����� ����;�2�D�V� h�������ˏԏ� ��
�7�.�@�R�d��� ����ǟ��П����� 3�*�<�N�`������� ï��̯����/�&� 8�J�\����������� ȿ�����+�"�4�F� Xυ�|ώϻϲ����� ����'��0�B�T߁� xߊ߷߮��������� #��,�>�P�}�t�� ������������ (�:�L�y�p������� ��������$6 Hul~������  Hg552��21�R7850J�614ATUP�'545'6VwCAMCRIb�UIF'28cN�RE52VR6�3SCHLI�C�DOCV�C�SU869'0^2EIOC�4�R69VESET�?UJ7UR68�MASKPR�XY{7OCOB#(3?+ &3j&[J6%53�H�(�LCHR&OPLGz?0�&MHCRS&]S�'MCS>0.'{552MDSW+7vu'OPu'MPRv&t��(0&PCMz�R0q7+ 2� �'5�1J51�80JP�RS"'69j&FR�DbFREQM�CN93&SN�BA��'SHLB�FM1G�82&H{TC>TMIL��TPA�TPT�XcFELF� �8�J95�T�UTv'95j&UE�V"&UECR&UF]RbVCC
XO�&wVIPnFCSC�F�CSG��IW�EB>HTT>Ra6��H;RVCGiW{IGQWIPGS�V�RCnFDGu'H7.�7R66J5']R�8R51
(6�(%2�(5V�J8�8�6�L=I% �84vg662R64�NVD"&R6�'R[84�g79�(4��S5i'J76j&Du0�gF xRTSF�CR�gCRXv&CsLIZ8ICMS�\Sp>STYnG6)7GCTO>��7�;NNj&ORS�&C �&FCB�FCFv�7CH>FCR"&�FCI�VFC�'JԗPO7GBfM�8OLnaxENDS&LU�&WCPR�7LWS�x�C�STxTE�gS�60FVR�IN�7IHaF�я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{���� ���/AS ew������ �//+/=/O/a/s/ �/�/�/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� �������� %�7�I�[�m�������Ǐُ�  ?H552���21�R78�5�0�J614�AwTUP7�5457��6�VCAM�C�RI��UIF7�2�8��NRE�52�v�R63�SCH��LICƚDOC�V�CSU�86�97�0F�EIOC�Ǜ4�R69v�EgSETW�u�J7u��R68�MASK^�PRXY��7�OCO��3W�����6�3�J65�53�6�H$�LCHƪO�PLGW�0�MH�CRǪS��MCS�V�0��55F�MD�SW���OP��M�PR���6�06�PCM��R0E˓�F�l��6�51f�51���0f�PRS��69��FRD��FRE�Q�MCN�93�6�SNBAכ%�SHLB�ME��ּ�26�HTCV�TMsIL�6�TPAV�oTPTX��EL�ē�6�8%�#��J9�5��TUT��95��UEV��UEC�ƪUFR��VCC�f�O��VIP��C;SC��CSGƚ$��I�WEBV�HTTV�R6՜��S����CG��IG��IP�GS'�RC��DGv��H7��R66f��5�u�R��R51*f�6�2�5v�#�)J׼��6��LU�5��s�v�4��66F�R�64�NVD��R�6��R84�79��4��S5�J7�6�D0uFR�TS&�CR�CR�X��CLI&�e�C�MSV�sV�STY:��6�CTOV�#��V�75�NN�ORqS����6�FCBV��FCF��CHV�F�CR��FCIF�F�C��J#��G
Mv��OL�ENDǪ�LU��CPR��L�u�S�C$�StT�E�S60�FVmRV�IN��IH�� �m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s�������軏͏ߏ�S�TD�LANG���0�B�T�f� x���������ҟ��� ��,�>�P�b�t��� ������ί���� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢϴ��� ������� �2�D�V��h�zߌߞ߰���RB=T
�OPTN���� ��'�9�K�]�o�������������DPN	���)�;�M�_� q��������������� %7I[m �������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu���� �����)�;�M� _�q���������ˏݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+�=� O�a�sυϗϩϻ��� ������'�9�K�]� o߁ߓߥ߷������� ���#�5�G�Y�k�}� ������������� �1�C�U�g�y����� ����������	-?Qc�f�������99���$FEAT_AD�D ?	����  	�#5GYk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ���������DEM�O y   �L�B�T߁� xߊ߷߮��������� ��G�>�P�}�t�� ������������ C�:�L�y�p������� ��������?6 Hul~���� ��;2Dq hz������  /
/7/./@/m/d/v/ �/�/�/�/�/�/�/? 3?*?<?i?`?r?�?�? �?�?�?�?�?O/O&O 8OeO\OnO�O�O�O�O �O�O�O�O+_"_4_a_ X_j_�_�_�_�_�_�_ �_�_'oo0o]oTofo �o�o�o�o�o�o�o�o #,YPb�� �������� (�U�L�^��������� ��ʏ����$�Q� H�Z���~�������Ɵ ����� �M�D�V� ��z�������¯ܯ� �
��I�@�R��v� ��������ؿ��� �E�<�N�{�rτϱ� �Ϻ��������A� 8�J�w�n߀߭ߤ߶� ��������=�4�F� s�j�|�������� ����9�0�B�o�f� x��������������� 5,>kbt� ������1 (:g^p��� ���� /-/$/6/ c/Z/l/�/�/�/�/�/ �/�/�/)? ?2?_?V? h?�?�?�?�?�?�?�? �?%OO.O[OROdO�O �O�O�O�O�O�O�O!_ _*_W_N_`_�_�_�_ �_�_�_�_�_oo&o SoJo\o�o�o�o�o�o �o�o�o"OF X�|����� ����K�B�T��� x�������ۏҏ�� ��G�>�P�}�t��� ����ןΟ����� C�:�L�y�p������� ӯʯܯ	� ��?�6� H�u�l�~�����Ͽƿ ؿ����;�2�D�q� h�zϔϞ�������� ��
�7�.�@�m�d�v� �ߚ��߾�������� 3�*�<�i�`�r��� ����������/�&� 8�e�\�n��������� ��������+"4a Xj������ ��'0]Tf �������� #//,/Y/P/b/|/�/ �/�/�/�/�/�/?? (?U?L?^?x?�?�?�? �?�?�?�?OO$OQO HOZOtO~O�O�O�O�O �O�O__ _M_D_V_ p_z_�_�_�_�_�_�_ o
ooIo@oRolovo �o�o�o�o�o�o E<Nhr�� �������A� 8�J�d�n�������я ȏڏ����=�4�F� `�j�������͟ğ֟ ����9�0�B�\�f� ������ɯ��ү���� �5�,�>�X�b����� ��ſ��ο����1� (�:�T�^ϋςϔ��� �������� �-�$�6� P�Z߇�~ߐ߽ߴ��� ������)� �2�L�V� ��z���������� ��%��.�H�R��v� ��������������! *DN{r�� �����& @Jwn���� ���//"/</F/ s/j/|/�/�/�/�/�/ �/???8?B?o?f? x?�?�?�?�?�?�?O OO4O>OkObOtO�O �O�O�O�O�O__0]  'XF_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX j|������ ���0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ����������
��.�   /�)�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ����� ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�� ������������ &�8�J�\�n������� ����������"4 FXj|���� ���0BT fx������ �//,/>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodo vo�o�o�o�o�o�o�o *<N`r� �������� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$�
4�8�+�N�`�r� �ߖߨߺ�������� �&�8�J�\�n��� ������������"� 4�F�X�j�|������� ��������0B Tfx����� ��,>Pb t������� //(/:/L/^/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�? �?�?�?�?�?O O2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�o�o�o�o�o�o &8J\n�� �������"� 4�F�X�j�|������� ď֏�����0�B� T�f�x���������ҟ �����,�>�P�b� t���������ί�� ��(�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢ� ����������� �2� D�V�h�zߌߞ߰��� ������
��.�@�R� d�v��������� ����*�<�N�`�r� �������������� &8J\n�� ������" 4FXj|��� ����//0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O �O�O�O�O�O�O __�$_6Y�$FEAT�_DEMOIN [ ;T�fP�<P}NTINDEX[[�jQ�NPILEC�OMP z�;���QiRIU��PSETUP2 �{�U�R��  N �Q�S_A�P2BCK 1|~�Y  �)7XDok%�_8o<P�P &oco9U�_�oo�oBo �o�oxo�o1C�o g�o��,�P� ����?��L�u� ���(���Ϗ^�󏂏 �)���M�܏q���� ��6�˟Z�؟���%� ��I�[�������� D�ٯh������3�¯ W��d������@�տ �v�Ϛ�/�A�пe� ���ϛ�*Ͽ�N���r� ��ߨ�=���a�s�� ��&߻���\��߀�� '��K���o���|�� 4���X������#��� G�Y���}������B� ��f�����1�Y�P�P�_ 2�P*�.VR8���*��������l P�C���FR6�:�2�V�T zPz�w�]PG<���*.Fo/"��	�:,�^/�STMi/�/ D/�-M/�/�H�/�?�'?�/�/g?�GIFq?�?�%�?D?V?�?�JPG�?O�%`O�?�?oO�
JSyOĢO��5C�OMO%
�JavaScri3pt�O�?CS�O&_��&_�O %Ca�scading �Style Sh�eetsR_��
A�RGNAME.D)T�_��� \�_S_еA�T�_�_�PDI'SP*�_���To��_�QLaZooCLLB.ZIwo2o$ K:\�a\�o�i�ACollabo�o��o
TPEINS�.XML�_:\�![o�QCusto�m Toolba�rbiPASSW�ORDQo��FR�S:\�dB`Pa�ssword Config���/� �(�e�������� N��r�����=�̏ a������&���J��� 񟀟���9�K�ڟo� ������4�ɯX��|� ��#���G�֯@�}�� ��0�ſ׿f������ 1���U��y��ϯ� >���b���	ߘ�-߼� Q�c��χ�߽߫�L� ��p��ߦ�;���_� ��X��$��H����� ~����7�I���m��� �� �2���V���z��� !��E��i{
� .��d��� �S�wp�< �`�/�+/�O/ a/��//�/8/J/�/ n/?�/�/9?�/]?�/ �?�?"?�?F?�?�?|? O�?5O�?�?kO�?�O O�O�OTO�OxO__ �OC_�Og_y__�_,_ �_P_b_�_�_o�_o Qo�_uoo�o�o:o�o ^o�o�o)�oM�o �o��6��l ��%�7��[��� �� ���D�ُh�z�� ��3�,�i������ ��ßR��v�������$FILE_D�GBCK 1|������� < �)
�SUMMARY.�DG!�͜MD:�U���ِDia�g Summar�y����
CONSLOG��n���ٯ����Consol�e log���	?TPACCN�t��%\�����TP �Accounti�n;���FR6:�IPKDMP.ZIPͿј
�ϥ����Excepti�on"�ӻ��MEMCHECK���������-�Memor?y Data�����(n )��RI�PE�~ϐ�%ߴ��%�� Pack�et L:���L��$�c���STAT���߭� %�A�Status<��^�	FTP�����	��/�mme?nt TBD2�^�� >I)ETHERNEw�
�d�u���﨡Ether�nJ�1�figur�aAϩ��DCSV�RF&���7������ verify� all:����{4��DIFF/���'���;�Q�dif�f��r�d���CHG01������A����,it�2���27@0���fx3�8��I �p��VTRNDIAG.LSu&8����� Ope���L� ��nost�ic����)�VDEV�DAT�������Vi�s�Device�+IMG��,/�>/�/:�i$Ima�gu/+UP E�S/�/FRS:�\?Z=��Upd�ates Lis�tZ?��� FLEXEVEN��/�/��?���1 UIF� EvM�M���-�vZ)CRSEONSPK�/˞�q\!O���CR_TAOR_PEAKbO�ͩPSRBWLD'.CM�O͜E2�O�\?.�PS_ROB�OWELS���:G�IG��@_�?d_���GigE�(O��Nߵ@�)UQHADOW__D_V_�_���Shadow ?Change�����dt�RRCME�RR�_�_�_oo���4`CFG Err{oro tailo� MA�k�CMSGLIBgoNo`o`�o|R�e��z0ic�oޭa�)�`ZD�0_O�os��ZDf�Pad�l �RNOTI�Rd����Notifi�c����,�AG ��P�ӟt��������� Ώ]�����(���L� ^�폂������G�ܟ k� ����6�şZ�� ~������C�د�y� ���2�D�ӯh����� ���¿Q��u�
�� ��@�Ͽd�v�Ϛ�)� ����_��σ�ߧ�%� N���r�ߖߨ�7��� [�����&��J�\� �߀���3����i� ���"�4���X���|� �����A�����w� ��0��=f��� ��O�s� >�bt�'� K���/�:/L/ �p/��/�/5/�/Y/ �/ ?�/$?�/H?�/U? ~??�?1?�?�?g?�? �? O2O�?VO�?zO�O O�O?O�OcO�O
_�O ._�OR_d_�O�__�_ �_M_�_q_oo�_<o �_`o�_mo�o%o�oIo �o�oo�o8J�o n�o��3�W� {�"��F��j�|� ���/�ď֏e�������0��$FILE�_FRSPRT � �������?�MDONLY 1|S��� 
 �)�MD:_VDA�EXTP.ZZZ�1�⏹�ț6%�NO Back? file ���S�6P�����>� �K�t�����'���ί ]�򯁯�(���L�ۯ p������5�ʿY�׿  Ϗ�$ϳ�H�Z��~� Ϣϴ�C���g���� ��2���V���cߌ�� ��?�����u�
��.�@���d��߈��C�VISBCKq�[���*.VD����S��FR:\��ION\DATA\���v�S�Vision VD��� Y�k����y��B��� ��x���1C��g ���,�P�� ��?�Pu �(��^��/ ��M/�q/�/>/�/ 6/�/Z/�/?�/%?�/ I?[?�/??�?2?D?��?9�LUI_CONFIG }S�����; $ 	�3v�{S�;OMO_O`qO�O�O�I#@|x�? �O�O�O__%\�OH_ Z_l_~_�_'_�_�_�_ �_�_o�_2oDoVoho zo�o#o�o�o�o�o�o 
�o.@Rdv� ������� *�<�N�`�r������ ��̏ޏ�����&�8� J�\�n��������ȟ ڟ쟃���"�4�F�X� j��������į֯� ���0�B�T�f��� ��������ҿ�{�� �,�>�P�b����Ϙ� �ϼ�����w���(� :�L�^��ςߔߦ߸� ����s� ��$�6�H� ��Y�~������]� ����� �2�D���h� z���������Y����� 
.@��dv� ���U�� *<�`r��� �Q��//&/8/ �\/n/�/�/�/;/�/ �/�/�/?"?�/F?X? j?|?�?�?7?�?�?�? �?OO�?BOTOfOxO �O�O3O�O�O�O�O_ _�O>_P_b_t_�_�_ /_�_�_�_�_oo�_�:oLo^opo�o�o$h�  x�o�c�$�FLUI_DAT�A ~���>�a(a�d�RESULT 3��ep ��T�/wiza�rd/guide�d/steps/?Expert�o= Oas���������z�Con�tinue wi�th Gpance�:�L�^�p����������ʏ܏� � �b-�a�e�0� �0`��c�a?��ps������� ��ҟ�����,�>� P��0ow��������� ѯ�����+�=�O��a�?�1�C�U�e�cllbs�ֿ���� �0�B�T�f�xϊϜ� [�����������,� >�P�b�t߆ߘߪ�i��{��ߟ�]�e�rip(pſ-�?�Q�c�u� ������������ �)�;�M�_�q����� �����������������`�e�#pTi�meUS/DST 	��������!3E�Enabl(�y��� ����	//-/?/
Q/�b�)�/M_q24|�/�/? ?)?;?M?_?q?�?�? Tf�?�?�?OO%O 7OIO[OmOO�O�Ob/�t/�/�/Z�"qRegion�O5_G_Y_ k_}_�_�_�_�_�_�_��America!�#o5oGoYoko}o �o�o�o�o�o�o��A�y�O�O3�O_qEditor�o�� �������+��=� � Touch Panel rs� (recommenp�)K������� Ə؏���� �2�D�|�%��I[qaccesoܟ�  ��$�6�H�Z�l�~������Conne�ct to Network��֯� ����0�B�T�f�x�(����x��@��}�䏟�,!��s Int?roduct!_4� F�X�j�|ώϠϲ��� �������0�B�T� f�xߊߜ߮��������� ɿ��" �i�{�������� ������/�A� �e� w��������������� +=�H�3��+�O��� �� 2DVh z�K������ 
//./@/R/d/v/�/ �/Yk}�/�?? *?<?N?`?r?�?�?�? �?�?�?��?O&O8O JO\OnO�O�O�O�O�O �O�O�/_�/1_�/X_ j_|_�_�_�_�_�_�_ �_oo0oBoS_foxo �o�o�o�o�o�o�o ,>�O_!_�E_ �������(� :�L�^�p�����So�� ʏ܏� ��$�6�H� Z�l�~���O��s՟ ���� �2�D�V�h� z�������¯ԯ毥� 
��.�@�R�d�v��� ������п⿡��ş '�9���`�rτϖϨ� ����������&�8� ��\�n߀ߒߤ߶��� �������"�4��=� �a��Mϲ������� ����0�B�T�f�x� ��I߮��������� ,>Pbt�E� ��i����( :L^p���� ���� //$/6/H/ Z/l/~/�/�/�/�/�/ ����/?�V?h? z?�?�?�?�?�?�?�? 
OO.O�ROdOvO�O �O�O�O�O�O�O__ *_<_�/??�_C?�_ �_�_�_�_oo&o8o Jo\ono�o?O�o�o�o �o�o�o"4FX j|�M___q_��_ ���0�B�T�f�x� ��������ҏ�o�� �,�>�P�b�t����� ����Ο�����%� �L�^�p��������� ʯܯ� ��$�6�G� Z�l�~�������ƿؿ ���� �2��S�� w�9��ϰ��������� 
��.�@�R�d�v߈� G��߾��������� *�<�N�`�r��Cϥ� g���ύ���&�8� J�\�n����������� ������"4FX j|������� ���-��Tfx �������/ /,/��P/b/t/�/�/ �/�/�/�/�/??(? �1U??A�?�? �?�?�? OO$O6OHO ZOlO~O=/�O�O�O�O �O�O_ _2_D_V_h_ z_9?�?]?�_�_�?�_ 
oo.o@oRodovo�o �o�o�o�o�O�o *<N`r��� ���_�_�_�_#��_ J�\�n���������ȏ ڏ����"��oF�X� j�|�������ğ֟� ����0����u� 7�������ү���� �,�>�P�b�t�3��� ����ο����(� :�L�^�pς�A�S�e� �ω��� ��$�6�H� Z�l�~ߐߢߴ��߅� ����� �2�D�V�h� z����������� �����@�R�d�v��� ������������ *;�N`r��� ����&�� G	�k-����� ���/"/4/F/X/ j/|/;�/�/�/�/�/ �/??0?B?T?f?x? 7�?[�?�?�?O O,O>OPObOtO�O�O �O�O�O�/�O__(_ :_L_^_p_�_�_�_�_ �_�?�_�?o!o�OHo Zolo~o�o�o�o�o�o �o�o �ODVh z������� 
���_%o�_I�s�5o ������Џ���� *�<�N�`�r�1���� ��̟ޟ���&�8� J�\�n�-�w�Q���ů ������"�4�F�X� j�|�������Ŀ��� ����0�B�T�f�x� �ϜϮ���������� �ٯ>�P�b�t߆ߘ� �߼���������տ :�L�^�p����� ������ ��$����� �i�+ߐ��������� ���� 2DVh '������� 
.@Rdv5� G�Y��}���// */</N/`/r/�/�/�/ �/y�/�/??&?8? J?\?n?�?�?�?�?�? ��?�O�4OFOXO jO|O�O�O�O�O�O�O �O__/OB_T_f_x_ �_�_�_�_�_�_�_o o�?;o�?_o!O�o�o �o�o�o�o�o( :L^p/_��� ��� ��$�6�H� Z�l�+o��Oo��sou� ���� �2�D�V�h� z����������� 
��.�@�R�d�v��� ������}�߯���� ٟ<�N�`�r������� ��̿޿���ӟ8� J�\�nπϒϤ϶��� �������ϯ��=� g�)��ߠ߲������� ����0�B�T�f�%� ������������� �,�>�P�b�!�k�E� ����{�����( :L^p���� w��� $6H Zl~���s��� ����/��2/D/V/h/ z/�/�/�/�/�/�/�/ 
?�.?@?R?d?v?�? �?�?�?�?�?�?OO ���]O/�O�O�O �O�O�O�O__&_8_ J_\_?�_�_�_�_�_ �_�_�_o"o4oFoXo jo)O;OMO�oqO�o�o �o0BTfx ���m_���� �,�>�P�b�t����� ����{oݏ�o��o(� :�L�^�p��������� ʟܟ� ��#�6�H� Z�l�~�������Ưد ����͏/��S�� z�������¿Կ��� 
��.�@�R�d�#��� �ϬϾ��������� *�<�N�`����C��� g�i�������&�8� J�\�n�����u� �������"�4�F�X� j�|�������q����� ��	��0BTfx ������� ��,>Pbt�� �����/�� ��1/[/�/�/�/�/ �/�/�/ ??$?6?H? Z?~?�?�?�?�?�? �?�?O O2ODOVO/ _/9/�O�Oo/�O�O�O 
__._@_R_d_v_�_ �_�_k?�_�_�_oo *o<oNo`oro�o�o�o gOyO�O�O�o�O&8 J\n����� ����_"�4�F�X� j�|�������ď֏� ����o�o�oQ�x� ��������ҟ���� �,�>�P��t����� ����ί����(� :�L�^��/�A���e� ʿܿ� ��$�6�H� Z�l�~ϐϢ�a����� ����� �2�D�V�h� zߌߞ߰�o��ߓ��� ���.�@�R�d�v�� ������������ *�<�N�`�r������� ����������#�� G	�n����� ���"4FX �|������ �//0/B/T/u/ 7�/[]/�/�/�/? ?,?>?P?b?t?�?�? �?i�?�?�?OO(O :OLO^OpO�O�O�Oe/ �O�/�O�O�?$_6_H_ Z_l_~_�_�_�_�_�_ �_�_�? o2oDoVoho zo�o�o�o�o�o�o�o �O_�O%O_v� �������� *�<�N�or������� ��̏ޏ����&�8� J�	S-w���cȟ ڟ����"�4�F�X� j�|�����_�į֯� ����0�B�T�f�x� ����[�m����󿵟 �,�>�P�b�tφϘ� �ϼ������ϱ��(� :�L�^�p߂ߔߦ߸� ������ ￿ѿ�E� �l�~�������� ����� �2�D��h� z��������������� 
.@R�#�5� �Y���� *<N`r��U� ����//&/8/ J/\/n/�/�/�/c�/ ��/�?"?4?F?X? j?|?�?�?�?�?�?�? �??O0OBOTOfOxO �O�O�O�O�O�O�O�/ _�/;_�/b_t_�_�_ �_�_�_�_�_oo(o :oLoOpo�o�o�o�o �o�o�o $6H _i+_�O_Q�� ��� �2�D�V�h� z�����]oԏ��� 
��.�@�R�d�v��� ��Y��}ߟ񟵏� *�<�N�`�r������� ��̯ޯ𯯏�&�8� J�\�n���������ȿ ڿ쿫���ϟ�C�� j�|ώϠϲ������� ����0�B��f�x� �ߜ߮���������� �,�>���G�!�k�� Wϼ���������(� :�L�^�p�����S߸� ������ $6H Zl~�O�a�s�� ��� 2DVh z�������� 
//./@/R/d/v/�/ �/�/�/�/�/�/�� �9?�`?r?�?�?�? �?�?�?�?OO&O8O �\OnO�O�O�O�O�O �O�O�O_"_4_F_? ?)?�_M?�_�_�_�_ �_oo0oBoTofoxo �oIO�o�o�o�o�o ,>Pbt�� W_�{_��_��(� :�L�^�p��������� ʏ܏���$�6�H� Z�l�~�������Ɵ؟ ꟩��/��V�h� z�������¯ԯ��� 
��.�@���d�v��� ������п����� *�<���]����C�E� ����������&�8� J�\�n߀ߒ�Q����� �������"�4�F�X� j�|��Mϯ�q����� ����0�B�T�f�x� �������������� ,>Pbt�� ���������� 7��^p���� ��� //$/6/�� Z/l/~/�/�/�/�/�/ �/�/? ?2?�; _?�?K�?�?�?�?�? 
OO.O@OROdOvO�O G/�O�O�O�O�O__ *_<_N_`_r_�_C?U? g?y?�_�?oo&o8o Jo\ono�o�o�o�o�o �o�O�o"4FX j|������ �_�_�_-��_T�f�x� ��������ҏ���� �,��oP�b�t����� ����Ο�����(� :�����A����� ʯܯ� ��$�6�H� Z�l�~�=�����ƿؿ ���� �2�D�V�h� zό�K���o��ϓ��� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� �����������#��� J�\�n����������� ������"4��X j|������ �0��Q�u 7�9�����/ /,/>/P/b/t/�/E �/�/�/�/�/??(? :?L?^?p?�?A�?e �?�?�/ OO$O6OHO ZOlO~O�O�O�O�O�O �/�O_ _2_D_V_h_ z_�_�_�_�_�_�?�? �?o+o�?Rodovo�o �o�o�o�o�o�o *�ON`r��� ������&��_ /o	oS�}�?o����ȏ ڏ����"�4�F�X� j�|�;����ğ֟� ����0�B�T�f�x� 7�I�[�m�ϯ����� �,�>�P�b�t����� ����ο�����(� :�L�^�pςϔϦϸ� ���ϛ�����!��H� Z�l�~ߐߢߴ����� ����� �߿D�V�h� z������������ 
��.������s�5� ������������ *<N`r1�� ����&8 J\n�?��c�� ����/"/4/F/X/ j/|/�/�/�/�/�/� �/??0?B?T?f?x? �?�?�?�?�?��?� O�>OPObOtO�O�O �O�O�O�O�O__(_ �/L_^_p_�_�_�_�_ �_�_�_ oo$o�?Eo Oio+O-o�o�o�o�o �o�o 2DVh z9_������ 
��.�@�R�d�v�5o ��Yo��͏���� *�<�N�`�r������� ��̟����&�8� J�\�n���������ȯ ��я������F�X� j�|�������Ŀֿ� ����ݟB�T�f�x� �ϜϮ���������� �ٯ#���G�q�3��� �߼���������(� :�L�^�p�/ϔ��� ������ ��$�6�H� Z�l�+�=�O�a����� ���� 2DVh z�������� 
.@Rdv� ����������/ ��</N/`/r/�/�/�/ �/�/�/�/??�8? J?\?n?�?�?�?�?�? �?�?�?O"O��/ gO)/�O�O�O�O�O�O �O__0_B_T_f_%? w_�_�_�_�_�_�_o o,o>oPoboto3O�o WO�o{O�o�o( :L^p���� ��o� ��$�6�H� Z�l�~�������Ə�o 珩o��o2�D�V�h� z�������ԟ��� 
���@�R�d�v��� ������Я����� ׏9���]��!����� ��̿޿���&�8� J�\�n�-��Ϥ϶��� �������"�4�F�X� j�)���M����߅��� ����0�B�T�f�x� ������������ �,�>�P�b�t����� ����{��ߟ����� :L^p���� ��� ��6H Zl~����� ��/����;/e/ '�/�/�/�/�/�/�/ 
??.?@?R?d?#�? �?�?�?�?�?�?OO *O<ONO`O/1/C/U/ �Oy/�O�O__&_8_ J_\_n_�_�_�_�_u? �_�_�_o"o4oFoXo jo|o�o�o�o�o�O�O �O	�O0BTfx �������� �_,�>�P�b�t����� ����Ώ������o �o�o[��������� ʟܟ� ��$�6�H� Z��k�������Ưد ���� �2�D�V�h� '���K���o�Կ��� 
��.�@�R�d�vψ� �ϬϾ�Ͽ������ *�<�N�`�r߄ߖߨ� ��y��ߝ�����&�8� J�\�n������� ���������4�F�X� j�|������������� ����-��Q� ������� ,>Pb!��� �����//(/ :/L/^//A�/�/ y�/�/ ??$?6?H? Z?l?~?�?�?�?s�? �?�?O O2ODOVOhO zO�O�O�Oo/�/�/�O _�/._@_R_d_v_�_ �_�_�_�_�_�_o�? *o<oNo`oro�o�o�o �o�o�o�o�O_�O /Y_����� ����"�4�F�X� o|�������ď֏� ����0�B�T�% 7I��mҟ���� �,�>�P�b�t����� ��i�ί����(� :�L�^�p��������� w���������$�6�H� Z�l�~ϐϢϴ����� ���ϻ� �2�D�V�h� zߌߞ߰��������� 
�ɿۿ�O��v�� ������������ *�<�N��_������� ��������&8 J\�}?�c�� ���"4FX j|������ �//0/B/T/f/x/ �/�/�/m�/��/� ?,?>?P?b?t?�?�? �?�?�?�?�?O�(O :OLO^OpO�O�O�O�O �O�O�O _�/!_�/E_ ?	_~_�_�_�_�_�_ �_�_o o2oDoVoO zo�o�o�o�o�o�o�o 
.@R_s5_ ��mo����� *�<�N�`�r������� gȍޏ����&�8� J�\�n�������c� �џ���"�4�F�X� j�|�������į֯� �����0�B�T�f�x� ��������ҿ����� ��ٟ#�M��tφϘ� �ϼ���������(� :�L��p߂ߔߦ߸� ������ ��$�6�H� ��+�=ϟ�a����� ����� �2�D�V�h� z�����]��������� 
.@Rdv����k�}������$FMR2_GR�P 1���� �C4�  B��	 ��9K6F@� a@�6G� � �Fg�fC��8R�y?�  x��66�X����875t��5���5`+�y�A�  /+BHx�w-%@S339%B�5[/l-6@6! �/xl/�/�/�/�/? �/&??J?5?G?�?k?��?��_CFG �TK�?�? O|O�9NO /
F0FA K@�<�RM_CHKTYP  ��$&�� ROMa@_MsINg@�����@u�R XSSB�3��� 7�O���C�O�O�5�TP_DEF_O/W  ��$W�IRCOMf@_��$GENOVRD�_DO�F��E]TYH��D dbUdKTo_ENB7_ KP�RAVC��G�@ �Y�O�_�?�oyo&oI* ��QOU��NAIRI< �@��oGo�o�o�o��C�p3��O:��B�+sL�i\�O�PSMT��Y�(�@
t�$HOS�TC�21��@s�5 MC���R{��� _ 27.00�1�  e�]�o��� ����K�ď֏���������	anonymous!�O�a�s�D���� �4���� ����D�!�3�E�W� i���������ï柀� .���/�A�S���� ��П����Ŀ��� �+�r�O�a�sυϗ� ����������'� n��������ϓ�ڿ�� ��������F�#�5�G� Y�k���υ������ ����B�T�f�C�z�g� �ߋ������������ 	-P�����u� �����(�:�< )p�M_q���� ����/$Zl I/[/m//�/��� �//�/D!?3?E?W? /?�?�?�?�?�/�? ./OO/OAOSO�/�/ �/�/�?�O?�O�O_ _+_r?O_a_s_�_�_ �O�?O�_�_oo'o��t�qENT 1��hk P!�_no  �p\o�o�o�o �o�o�o�o�o: _"�F�j�� ���%��I��m� 0���T�f�Ǐ��돮� �ҏ3���,�i�X��� P���t�՟��៼�
� /��S��w�:���^� �����������ܯ=�� �QUICC0�J�&�!192.�168.1.10c�X�1��v�8��\��2�ƿؿ9�!R�OUTER:��!���a��PCJ�OG��e�!*� ��0��U�CAMgPRT�϶�!�����RTS���x�� !Softw�are Oper�ator Pan�elU߇���7kNA�ME !Kj!�ROBO����S_�CFG 1�Ki� �Au�to-start{ed�DFTP�Oa�O�_���O���� ������E_�.�@�R� u�c�	����������� cN:�L�^�;r���R �������� %H�[m� ��jO|O�O�O4!/ hE/W/i/{/�/T�/ �/�/�/�//�//?A? S?e?w?�?����? ?�?</O+O=OOO? sO�O�O�O�O�?`O�O __'_9_K_�?�?�? �?�O�_�?�_�_�_o #o�OGoYoko}o�o�_ 4o�o�o�o�of_ x_�_g�o��_�� ���o��-�?�Q� tu��������Ϗ� (:L^`�2��q� ����������ݟ�� �%�H�ʟ[�m���� ������� �ί4�!� h�E�W�i�{���T��� ÿտ�
�Ϟ�/�A��S�e�w����_ER�R ��ڇϗ�P�DUSIZ  j�^6����>��?WRD ?(�����  guest���+��=�O�a���SCD_�GROUP 3��(� ,�"�IF�T��$PA��OM�P�� ��_S�H��ED�� $C��COM��TTP�_AUTH 1���� <!iPendanm�x�#��+!KAREL�:*x���KC������VISION SET��@(����?�-�W�R� ��v������������������G�CTRL K���a�
��FFF9E3���FRS:D�EFAULT��FANUC W�eb Server�
tdG����/�� 2DV��W�R_CONFIGw ���������IDL_C_PU_PC� �sB���� BH��MIN����GNR_IO���������HMI_EDI�T ���
 ($/C/��2/k/V/�/ z/�/�/�/�/�/?�/ 1??U?@?y?d?�?�? ./�?�?�?�?OO?O QO<OuO`O�O�O�O�O��O�O�O__;_�N�PT_SIM_D�O�*NSTA�L_SCRN� ��\UQTPMOD�NTOL�Wl[�R�TYbX�qV�K�E�NB�W�ӭOL_NK 1����� o%o7oIo[omoo�R_MASTE��Y�%OSLAVE ���ϮeRAMCOACHE�o�ROM�O_CFG�o�S�c�UO'��bCMT�_OP�  "��5sY�CL�ou� _AS�G 1����
 �o������ �"�4�F�X�j�|���\�kwrNUM�����
�bIP�o�gRTRY_CN@uQO_UPD��a���1 �bp�b��n��hM��аP}T?��k ��._������ ɟ۟퟈S���)�;� M�_�q� �������˯ ݯ�~��%�7�I�[� m��������ǿٿ� ����!�3�E�W�i�{� 
ϟϱ��������ψ� ��/�A�S�e�w߉�� �߿���������+� =�O�a�s���&�� ����������9�K� ]�o�����"������� ��������GYk }��0���� �CUgy� �,>���	// -/�Q/c/u/�/�/�/ :/�/�/�/??)?�/ �/_?q?�?�?�?�?H? �?�?OO%O7O�?[O mOO�O�O�ODOVO�O �O_!_3_E_�Oi_{_ �_�_�_�_R_�_�_o o/oAo�_�_wo�o�o �o�o�o`o�o+ =O�os���� �\n��'�9�K� ]����������ɏۏ�i�c�_MEMBE�RS 2�:�   $:� ���v����1���RCA_AC�C 2���   [~��R 	* �  (�0 5+�Pl�l�l��( �@�����  l���a�B�UF001 2��n�= ��u0�  u0����U
�
�+
�9
�UJ
�X
�j
�z�߈ � Q���J� J�/J�@J�O�J�`J�pJ��J���J��u0�e����u0X�ho��u0��ܲ���¤¤#�¤3¤C¤R¤V�0��Q��f���m�I������t���u0��bX�����u�0�UP�|R�@�H������u0�[�[������Z��Z�}�R�h[Ȇ�U�%�4�F�U�g�v�!��U�����������ߙ2���s�P������ !��)��1��9�� A��I���Q�R�X��� a���i���q���y��� ������������������t(������ ïկ���������R� ��)�L�(��0�s��8�s���@�Rh xH�U  P�\�Y��k�}�������ſ׺!��S@ߙ3����  ����'��)� 7��9�G��I�W�^� Y�g�^�i�w�^�y��� ^≢��^♢��^⩠ ^�1���^���l����� ���������������� ������l� ���� ����/����8�l� @�N�I�g�Q�N�b�N� j�N�r�N�z���� ����������� �������3��� �������ٲ��~ݖCFG 2�n�� 4l��
l�Jl�<l�47ۘ�HIS钜n� ��� 2025�-11-3�l��    #� &f  'c "珪�  ��*6X�`�hl��}pl�$  x {��8 �l�;W� � 7 �� �-ɔ/l�[}�p29}	7v�����������   % �� �  -�R ' *� l��B��aN/`/r/�/�/�/ �/�/�/�/'/9/&?8? J?\?n?�?�?�?�?�? �/?�?O"O4OFOXO jO|O�O�O�?�?�O�O �O__0_B_T_f_x_ �O�O�O�_�_�_�_o o,o>oPo�O��[Tm
8 c� 8� ��o�o�6d� �b�� �b� +  X��  X�  dT!qc	,: J�� 1r�oO=O�_���������":$�a 2�a ,*q 1  \�_�_m� �������Ǐُ��� ��_X�E�W�i�{��� ����ß՟��0��� /�A�S�e�w������� ��������+�=� O�a�s��������� ߿���'�9�K�]πoρ�J�Ѐo�o

eq� �������� ��� ��� ��� eq� G^�## o�]o������� �����#�5����2��� Z� �־�п ������������ &�8�o��n������� ����������G�Y� FXj|���� ��1�0BT fx�����	 //,/>/P/b/t/��/�/�Ϙ�I_CF�G 2��� H�
Cycle �Time�Bu{sy�Idl�"^�min�+1�Up�&�R�ead�'Do�w8?�` 1�#C�ount�	Num �"����<��zb�qaPROG�"�������)�/softpar�t/genlin�k?curren�t=menupa�ge,1133,1�/OO/OAO3b5�leSDT_ISO_LC  ���p��/J23_DSP_ENBL�vK0~�@INC ��M|�ӄ@A   ?&p�=���<#�
<�A�I:�o���N`_���O<_�GOB�0�C�CF�1�FVQG_�GROUP 1�vvK	r<�P�C�٢_D_?���?�_��Q�_o.o@o�_ dovo�o�o��,_NY�G_IN_AUT�ODԫMPOSRE�^_pVKANJI_�MASK v�HqR�ELMON ��˔?��y_ox������.6r�3��7ĲC���u�o�DKCwL_L�`NUML���EYLOGGINGDЫ���Q�E�0�LANGUAGE� ��~���DEFAULT� ����LG�!���:2�?�W��80H  ���'~��  � 
���囊�GOUF ;���
��(UT13:\��  �-� ?�Q�h�u���������ϟ�����(g4�8�i�N_DISP ���O8�_�_��L�OCTOL����D�z`�A�A��GBO_OK ���d�1
�
�۠#���� �#�5�G�Y�i���3{�W�	��쉞QQJ�¿Կ1��_BU�FF 2�vK 	���25
�ڢVB�&�7 Coll�aborativ �=�OΗώϠϲ��� ������'��0�]�T��fߓߊߜ��DCS ��9�B�Ax����Rh�%�-�?�Q���I�O 2��� ���Q���� ����������*�<� N�b�r����������������&:e�E_R_ITMsNd�o ������� #5GYk}����������hS�EV�`�MdTYPsN�c/u/�/
-��aRST5���SC�RN_FL 2�
s��0����/??`1?C?U?g?�/TPK��sOR"��NGNA�M�D��~�N�UPS�_ACR� �4D�IGI�8+)U_�LOAD[PG �%�:%T_NO�VICEt?��MA?XUALRM2��a����E
ZB�1_�P�5�` ��y�Z@CY��˭�O+���ۡ��D|PP 2�˫ �Uf	R/_
_C_ ._g_y_\_�_�_�_�_ �_�_�_oo?oQo4o uo`o�o|o�o�o�o�o �o)M8qT f������� %��I�,�>��j��� ��Ǐُ�����!�� �W�B�{�f������� ՟����ܟ�/��S� >�w���l�����ѯ�� Ư��+��O�a�D����p���RHDBGDEF ��E�ѱO���_LDXDIS�A�0�;c�MEMO�_AP�0E ?�;
 ױ��3� E�W�i�{ύϟϱ�Z@�FRQ_CFG k��G۳A ���@��Ô�<��d%��� ������B��K{��*i�=/k� **:tҔ� g�y�ߔ��߱����� �����J�Es��J d�����,( H���[�����@�'� Q�v�]����������������*NPJI�SC 1��9Z� ������ܿ������	Zl_MST�R �#-,SC/D 1�"͠{ �������� //A/,/e/P/�/t/ �/�/�/�/�/?�/+? ?O?:?L?�?p?�?�? �?�?�?�?O'OOKO 6OoOZO�O~O�O�O�O �O�O_�O5_ _Y_D_ i_�_z_�_�_�_�_�_ �_o
ooUo@oyodo �o�o�o�o�o�o�o�?*cN�M�K���;љ$�MLTARM��u�N��r ���հ��İMETP�U��zr��CN�DSP_ADCO�L%�ٰ0�CMNT6F� 9�FNb�f�>7�FSTLI��x�4 �;ڎ�s�����9�POSCFz��q�PRPMe���STD�1�;; 4�#�
v��q v�����r�������� ̟ޟ ���V�8�J� ��n���¯��������9�SING_CH�K  ��$MODA���t�{�~~2�DEV 	��	MC:f�HS�IZE��zp�2�T�ASK %�%�$1234567�89 ӿ�0�TR�IG 1�; lĵ�2ϻ�!�bϻ�F��YP����H�1��EM_INF 1��N�`)AT&FV0E0g����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ��2��H6�^���R����A�߶�q�������� ��5������ ߏ�B߳�������� ���1�C�*�g��,� ��P�b�t������ R�?���u0�� ������������� M q���Z� ��/�%/��[/  2�/�/h�// �/�/�3?�/W?>?{? �?@/�?d/v/�/�/O �//OAOx?eO?�ODO��O�O�O�O_�NIT�ORÀG ?z� �  	EXESC1~s&R2,X3,XE4,X5,X��.V7,X8,X9~s'R�2�T +R�T7R�TCR�TOR�T [R�TgR�TsR�TR�TT�R�S2�X2�X2�XU2�X2�X2�X2�XU2�X2�X2h3�X�3�X37R2�R_G�RP_SV 1��� (꡿i���?�4������>��4����>؋�a���_�D�B���cION_�DB<��@�zq W �zp�zp�Y��1u'�>w��p���p�Y��@N 2pZ2p>{n�poY�-ud1������8�PG_JOG� �ʏ�{
�2��:�o�=���?����@0�B��~\�n����@����H�?��C�@eqpȏڏ���  ������qL_NAM�E !ĵ8���!Defaul�t Person�ality (from FD)qp�0�RMK_ENOgNLY�_�R2�a� 1�L�XL��8�gpl d����şן���� �1�C�U�g�y����� ����ӯ���	���� 
�<�N�`�r�������p��̿޿� :� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w���������������+��<�Se w�������x��A�a��AB�Bw��Pf ������/!/ 3/E/W/i/{/�/�/�/ ���/�/??/?A? S?e?w?�?�?�?�?�? �?�?�/�/+O=OOOaO sO�O�O�O�O�O�O�O __'_9_&O�S��#�x_�]�rdtS�� �_�]�_�_�W�����S�"oe_oXoa  ��qogoyo�o�o�o�o@�ouP�p"|����	`[oUgy8qK��A\����s� AA��y@h�Q�Q��e"���Tk\$���  ��P��PE�xC�  �I�@oa�<o��p��� ����ߏ
f�Q*������0��PCr� �� 3r �.� �@D�  A�?��G�-�?.I�.@I��A����  ;��	lY�	 ��X  ������� �,? � ������uPK�o������]K��K]�_K	�.��w��r_	����@
��)�b�1�����I��Y�����T;�fY�{S���3����I�>J���;�Î?v�>��=�@�����E��R ѯעZ���wp��u��� D!�3���7pg  �  ��9�͏W���	'�� � u�I�� �  ���u��:�È��ß�=��ͱ���@��ǰ�3��\�"3�E�&���N�pC�  'Y�&�Z�i�bb�@f�i�n�C��D��I�C����b��r���`����B�p�Ŕq���}ر�.DzƏ<ߛ�`�pK�pߖ����������А G4P����.z���d  �Pؠ?�ff�_��	��C 2p>�P���8.f�t�>L���U���	(.��P���������
ĉ��� x��;e��m��KZ;��=g;�4�<�<����%�G���3����p?fff?�ذ?&S���@==0e�?��q�+ �rN�Z���I���G��� 7���(�����!E 0iT����+��F�p���# ��D��w�� �����//=/ (/a/L/�/p/��/� p�6�/Z#?�/ ?Y? k?}?��?�?>?�?�?@�?�?�?1O�����KD�y^KCO�OO�O���ذO�O�O�Oai����J��}�DD1���.�D��@�AmQ�a��9N,ȴA;��^@��T@|�j@$�?��V�>�z�ý���=#�
>�\)?��
=��G�-]�{=����,��C+�?�Bp���P���6��C98R����?N@��(���5-]G��p�Gsb�F��}�G�>.E��VD�Kn����I�� F��W�E��'E����D��;n����I��`E��G��cE�?vmD���-_�o Q_�o�o�o �o$ H3X~i��� ������D�/� h�S���w�������� я
���.��R�=�v� a�s�����П����ߟ ��(�N�9�r�]��� ������ޯɯۯ��� 8�#�\�G���k����� ��ڿſ���"��F� 1�C�|�gϠϋ��ϯϠ��������P(�Q3g4�] �����Q��	�9�Oߵ53~�m8m��aҀ5Q�߫ߎaғ����ߵ1�������1��U�PC�y�g��%P�P���!�/��'���
���<.������4�;� t�_������������� ��:%��/�/d������ ��7%[I m���027��  B�S@J@�C%H#PzS@�0@ZO/�1/C/U/g/y/�-�#���/�/�/�/�/�3?Y�3�� @�3�%�0�0�13��5
 ?f?x?�? �?�?�?�?�?�?OO�,O>OPO�Z@1 ����ۯ�c/�$M�R_CABLE �2ƕ� ��TT�����ڰO�� �O�)�@���C_��� _O_u_7_I__�_�_ �_�_�_o�_�_oKo qo3oEo{o�o�o�o�o �o�o�o�oGm/�K!�"���O�����ذ�$�6����*Y�** �CO�M ȖI�����92�%%� 2345678'901���� ��Ï���� � !� �!
���Mn�ot sent �b��W��T�ESTFECSALGR  eg�*"!d[�41�
k�������$pB����������� 9UD�1:\maint�enances.�xmlğ�  �C:�DEFA�ULT�,�BGRP� 2�z�  �����%  �%!�1st clea�ning of cont. v��ilation +56��ڧ�!0�����+B��*������+��"%��me�ch��cal c�heck1�  ��k�0u�|�� ԯ����Ϳ߿�@���?rollerS�e�w�ū��m�ϑϣ����@�Basic� quarterCly�*�<�ƪ,\��)�;�M�_�q�8�MXJ��ߓ "8��� ���ߕ �����+�=��C�g�ߋ�ʦ�߹���������@�Overha�u�ߔ��?� x� I�P����}���������� $n���� ���)l�ASew� ����� � +=O�s��� ����/R�9/ �(/��/�/�/�/�/ /�/�/N/#?r/G?Y? k?}?�?�/�???�? 8?OO1OCOUO�?yO �?�?�O�?�O�O�O	_ _jO?_�O�Ou_�O�_ �_�_�_�_0_oT_f_ ;o�__oqo�o�o�o�_ �oo,oPo%7I [m�o��o�o� ���!�3��W�� ������ÏՏ�6� ���l����e�w��� ������џ�2��V� +�=�O�a�s���� ��ͯ����'�9� ��]�������⯷�ɿ ۿ���N�#�r���Y� ��}Ϗϡϳ������ 8�J��n�C�U�g�y� ���ϯ������4�	� �-�?�Q��u����� �ߞ���������f� ;������������ �����P���t�I [m����� �:!3EW� {��� ��� //lA/��w/���/�/�/�/�/X*�"	� X�/?.?@?�)B a/o?m/o%w?�?�? }?�?�?OO�?�?OO aOsO1OCO�O�O�O�O �O__'_�O�O]_o_ �_?_Q_�_�_�_�_�_��\ Џ!?� ; @�! M?Ho Zolo�&4o�o�o�o�(�*�o** F�@ �Q�V�`o�'9�o]o�����/^&�o��� ��/�A�S�e��� #�����я����� +�q�����7������� k�͟ߟ��I�[��� K�]�o���C�����ɯ���o$�!�$M�R_HIST 2���U#�� 
 �\7"$ 2345?6789013�;���b2�90/���� [���./����ǿٿ F�X�j�!�3ρϲ��� {��ϟ�����B��� f�x�/ߜ�S����߉� �߭��,���P��t����=��$�SKCFMAP  �U�&��b
�� ����ONREL  �$#�������EXCFENB��
����&�FNC�-��JOGOVL�IM�d#�v���K�EY�y���_�PAN������R�UNi�y���SFSPDTYPM�<���SIGN���T1MOTk�����_CE_GRP7 1��U��+� 0�ow�#d�� ����&�6 \�7y�m� ��/�4/F/-/j/ !/t/�/�/�/{/�/�/�/?�+��QZ_E�DIT
����TC�OM_CFG 1����0�}?�?�? }
^1SI �NB����?�?���?�$O����?XO78T__ARC_*��X�T_MN_MO�DE
�U:_S�PL{O;�UAP_�CPL�O<�NOCHECK ?��/ �� _#_ 5_G_Y_k_}_�_�_�_��_�_�_�_oo��N�O_WAIT_L�	S7> NTf1�����%��qa_ERMRH2������� ?o�o�o�o��O�Gj�@O�cӦm| �	.GA�f��A�;?�
[��>����e^B/Aq���<���?���)��n�b_PARAM�b����vHO��w
�.�@� = n�]�o� w�Q�����������`Ϗ�)���w�[��m� �����ODRD�SP�C8�OFFSET_CARI0��OǖDISԟœS;_A�@ARK
T9�OPEN_FIL�E��1T6�0OPTION_IO�����K�M_PRG ;%��%$*�����'�WO��N	��
��ǥ��w ����r����	 ������>d���R�G_DSBL  �����jN���R�IENTTO�f��C�����A ���U�@IM_DS����r��V��LCT �{mP2ڢ�3̹���d��%���_P�EX�@���RAT��G d8��̐UOP װ�:�����S�e�Kωϗ��$��r2G�L�X�LȚ�l 㰂�������'�9� K�]�o߁ߓߥ߷��� �������#�5�G���2��v������� ������e�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?�q1�~?�?�?�? �?�?�?�?O O2ODO^�yA�a�m? ~N��~O�O�P�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�O �Oo$o6oHoZolo~o �o�o�o�o�o�o�o  �_oVhz�� �����
��.��@�R�d�QOES��(����Ԣd�ӏ� ʏ��������Y�D�}�0��r������� ��ԟڟ���p���=�4M��q�	`����x����c�:�o��¯ԯ����A�C  �k�C�C�ڰe"ڰ���O���  ����-���)�C�  �t�k���g�����Կ ��ѿ
�5���_:�ĳ��OU������H��n��� � ^��\� @D�  &p�?�v�\�?:px��:qC4r�p�(�� � ;�	l��	 ��X � ������ ��, � �x������Hʪ�������H���Hw�zH����ϝ�8�B���B��  Xѐ�`�o�*��'3����t�>u����fC{ߍ��:pB\��
�Ѵ9:qK�t�� �����$���*��� D�P�^��b�g  �  �h������)�	'� �� ��I� ��  ��'�=��������t�@����!�b��^;bt�U�(�N��r� ' '��E�C�И�t�C�И��ߗ���jA��@�����%�B �� ��,���H:qDz�k�ߏz����������А 4P���:uz:���	�f��?�faf'�&8� ]��m�8:p��>!L�����$�(:p�P��	������:�� x�;e�m�"�KZ;�=g�;�4�<<�0��E/Tv��b����?fff?�?y&� )�@=0�%?��%_9��}! ��$�x��/v��/f'�� W,??P?;?t?_?�? �?�?�?�?�?O�?(O OLO�/�/�/EO�OAO �O�O�O�O_�O_H_ 3_l_W_�_{_�_�_1� �_A���eO+o�ORoo Oo�o�o�oK/�o�omo �o*'`+�,�zt���CL�H<��}?����X�
������u�����D1�/n�t�x�p�q��@I�h~�,ȴA;�^@���T@|j@�$�?�V�n��z�ý��=�#�
>\)?��
=�G�����{=��,���C+��B�p����6���C98R����?}p��(��5���G�p�G�sb�F�}�G��>.E�VD��KL����I��� F�W�E���'E���D���;L����I���`E�G���cE�vmD���\�՟��ҟ� ��/��S�>�w�b��� ����ѯ������� =�(�:�s�^������� ��߿ʿ�� �9�$� ]�Hρ�lϥϐϢ��� ������#��G�2�W� }�hߡߌ��߰����� ���
�C�.�g�R�� v��������	��� -��Q�<�u�`�r��� ����������'�M�(�34�]O!���8h~�%3~�m���ǀ5Q��������!���   `N�r��J	eP@"P��Q�_�/V/9/$/]/H)����c/j/�/�/�/ �/�/�/�/!??E?0? i?T?"&�_�_�?�?�8��?�?O�?OBO 0OfOTO�OxO�O�O�O��O2f?_  B���pyp$QCHR�z�p@�N_`_r_�_�_�_�]c�O�_�_0oo+o?�Bc�� @d4��QJc�D
 2o�o�o�o�o�o�o %7I[m���oa ������c/�$PARA�M_MENU ?� � � DEF�PULSE��	�WAITTMOU�T�{RCV� �SHELL_�WRK.$CUR�_STYL�p�"�OPT8Q8�PT�BM�G�C�R_DECSN�p����� ���������-�(� :�L�u�p��������q�SSREL_ID�  ��̕U�SE_PROG �%�z%���͓C�CR�pޒ��s1�_HOST !�z#!6�s�+�T�=����V�h���˯*�_�TIME�rޖF�~�pGDEBUGܐ��{͓GINP_F�LMSK��#�TR\2�#�PGAP� ���_b�CH1�"�TWYPE�|�P�� ������0�Y�T� f�xϡϜϮ������� ���1�,�>�P�y�t� �ߘ��߼�����	�� �(�Q�L�^�p��%�WORD ?	�{
 	PR��p#MAI��q"3SUd���TE��p#��	1���COL�n%��!���L�� �!��F�d�T�RACECTL �1� �q }� �#�����_�DT Q�� ��z�D �� �^a����c`�������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O__/_A]B_T_v_ �_�_�_�_�_�U��� oo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�.�oP�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/Dϒ/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D��V�h�z�����������$PGTRACE�LEN  �� � ������Ά_UP _�����������΁_CFoG ����*��
���*�:�D��O���O�  ��O��DEFSPD� ��������΀H_CONF�IG ����� ����dĔ�&݂ ��ǑP^�a�l㑹��΀IN�?TRL ��=��8^���PE��������*�ÑO��΀LID���	~T�LLB 1ⳙ_ ��BӐsB4��O� �𼧶��Q� <<7 ��?��� ����M�3�U���i� ��������ӿ��	�7�T�Ϣk�b�tϡπ诚��������S�G�RP 1爬����@A!���4�I���A �C�u�C�OCWjVF�/��Ȕ`a�zي�ÑÐ�t�0�ޯs���´�ӿ���B������������A�S�&�B3�4�_������j���������	� B�-���Q���M�������  Dz����.� ����&L7p[ ��������6!Zh)w�
V7.10be�ta1*�Ɛ@��*�@�) @ߺ+A Ē?���
?fff>�����B33�A�Q�0�B(���A���AK��h����//('/9/P�p*�W�ӑ��n/�/�%���R��fh���� *���P2�LR��/�/@�/�/�/H?�Ĕ�I�u�&:���?��x?��?A���P!\3 Bfu�B��?�5BH�3�[4��o��4�I�[45��/B\3x3Dx�?YO�?aOkO}O�<<�R@��O�C�O�O��O�O�DA�X�KNO?W_M  Z�%��X�SV 賚ڒ]��_�_�_?��_�_�_o����W�M�+�鳛 ��	~@�3#���_��o�\A��
]bV4�@u��u��e��o�l,�X�MR+��JmT3?��W�1C{��OADBANFW�DL_V�ST+�1 k1����P4C� ��[��i/��� ��?�1�C���g�y� �������ӏ�*�	�@�`�?�Q�c��w2�|8Va�up�<ʟ����p3��Ɵ؟Ꟃw4 ��+�=��w5Z�l�~����w6����ѯ㯂�w7 ��$�6��w8`S�e�w����wMAmp�������OVL/D  ��yo���rPARNUM � �{+þ�?υqS[CH�� �
��pX���{s��UPDX��)ź��Ϧ�_CMPa_@`���p|P'yu~�ER_CHK���yqbb3��.��RSpp?Q_MO�m��_}ߥ�_REWS_G�p쩻
� e�����0�#�T�G�x� k�}��������������׳�������� �:�Y�^���Y�y��� ���Ӭ����������� ����R�6UZ��ӥ�u����V �1�FvpVa@k��p��THR_ICNRp��(byudoMASS Z)�MNGMON_�QUEUE �P�uyvup\!��N��UZ�NW��ENqD��߶EXE�����BE���O�PTIO��ۚP�ROGRAM %z%��~Ϙ?TASK_I��.OCFG �zx+�n/� DATACcm�+�0P�up 2 �?�?/?A?S?]51  s?�?�?�?�?�6p1�?��?�?O"O,F�!IN+FOCc��-��bd lO~O�O�O�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_�_�_�/A@FD���, 	��!��K�_�!�)fN!fECNB��0m��Pf2Yo�khG�!2�0k �X,		d�=���·o���e�a$��pd��i�i�g_E?DIT ��/%�7����*SYS�TEM*upV9.�40107 cr7�/23/2021� A��Pw���PRGADJ_�p  h $X|[�p $Y�xZ�xW�xқtZқt?SPEED_�p�p�$NEXT_CYCLE�p��q�{FG�p ��p�ALGO_V ��pNYQ_FRE�Q�WIN_TYuP�q)�SIZ1�O�LAP�r!�[���M+����qCRE�ATED�r�IF�Y�r@!NAM�p�%h�_GJ�STA�TU��J�DEBU�G�rMAILTI:����EVEU���LAST�����tE�LEM� � ?$ENAB�rN��EASI򁼁AX;IS�p$P߄������qROT_R9A" �rMAX ��qjE��LC�AB
�y��C D_LVՁ`�BAS��`�1�{�r��_� ��$x����RM� RB�;�D�IS����X_SP8o�΁�� ��t�P�� | 	� �2 \�AN�� �;������Ӓ�� �0�P�AYLO��3�V�_DOU�qS���p�t�PREF� ( $GRID��E
���R���Y:����OTOƀ�q�  �p��!��p��k�OXY�� � $L��_�PO|�נVa�S�RV��)���DI?RECT_1� �U2(�3(�4(�5(��6(�7(�8��qFꔑA�� $V�ALu�GROU�P�����F�� !��@!��q�����RAN�Ĳ���R��/���TO�TA��F��PW��I=!%�REGEN#�8�������/���ڶnTzЉ���#�C_S����8�(�V[�p'���4���GRE���w���H��D�����V�_H��DAY3�V���S_Y�Œ;�S�UMMAR��2� $CONFIG_SEȃ���ʅ'_RUN�m�C�С�_$CMPR��P�GDEV���_�I��ZP�*��q��EN_HANCE�	��
���1���IN	T��qM)b�q�2�K����OVRo�P�Gu�IX��;���O�VCT�����v�
 �4 ����a˟���PSLG"�� \ �;��?�1�ⷁSƁϕc�U@�����Ò�4�U���]�Tp� (�`�-��rJ<�O� C�K�IL_MJ���V�N�+��TQn{�N45���C�ULȀD�5V(�C6�P_�຀�@�MW�V1V�V1�d�2s�2d�3s�3
d�4s�4d��'�	�`������p	�IN	�VIB1qp1� 2P!pq/,3 3,4 4,�p?��;� �A���N�������;PL��TORr3�p	��[�SAV���d�MC_�FOLD 	�$SL�����Mb,�I��L� �p�L�b��KEEP__HNADD	!K�e�UCCOMc��k��
�lOP����pl��lREM�k��΢�Կ�U��ekHP�W� KSBM���ŠCOLLAB�|�Ӱn��n�+�I�T�O��$NO�L�FCALX� �D�ON�r����� ,��FL���O$SYNy,M��C=����UP_D�LY�qs"DEL�A� ����Y(�AD���$TABTP�_R�#��QSK;IPj% �����OR� �E�� P_ ��� �)���p7�� %9��%9A�$:N�$:[��$:h�$:u�$:��$:9�q�RA�� �X�����MB�N�FLIC]��0"�Ux!�o���NO_H� ��\�< _SWIT�CHk�RA_PA�RAMG� i��p��U��WJ���:Cӣ�NGRLT� OO�U�����X�<A���T_Ja1F�rA}PS�WEIGH]��J4CH�aDOR��aD��OO��)�2�"_FJװ���sA�AV�L�C�HOB.�.����J2�0�q$�EX2��T$�'QIT��'Q��pG'Q-�G��RD�C�m" � ��<��
R]��
H���RGEA��4��U�FLG`g��H��sER	�SPC6R��rUM_'P��2T�H2No��@Q o1 @ED�����  D ��وIi�2_P�2�5cS�ᰁ+�L10�_CI�WQd� �pk����UՖ�D��zaxT�p�Q (�;a��c��޲+�i���pe��` P>`DESIGRb$�VL1:i1Gf�c�g;10�_DS��D�|��w�POS11�q l�pr��x1C�/#AT�B��U
WusIND��}�mq�Cp�mq`B	�HOMME�r 	aBq2GrM_q���`!
@s3Gr��� �(�$�6�4GrG�Y�0k�}����� �a�q5Grď֏����(���?t6GrA�S��e�w�����0�7Gr���П�����6�8Gr;�M�_�q������uS �q    �@sM��P6��K@��! T`M��&M�IO��m�I��2�OK _OPy��� �ػQ�2�pWE"� 7�x EQAE� � #s%Ȳ$D;SBo�GNA�b� C�P�bd�RSw232S�$ �iPr��xc�ICE<@�%�PE`2� @IT���P�OPB7 1�F7LOW�TRa@2��U$�CUN��`�A�UXT��2Ѷ�ER�FAC3İUU�o����CH��'% t<_9�E���A$FREEF'ROMЦ�A�PX q�UPD"YbA�3PT.�pEEX0����!�FA%bҲ���RV�aG� &�  ��E�" 1�AL�  �+�jc�'��D�  2& ��S\PcP(
 ' �$7P�%�R�24SP��T�`AXU���DSP���@�W���:`$��RNP�%�@��z��K��_MIR������MT��AP����P"�qD�QSY�z������QPG7�B�RKH���ƅ AXI�  ^��i�����1 ����BSO�C���N��DUM�MY16�1$S�V�DE��I�FS�PD_OVR7d9� D����OR��֠N"`��F_����@�OV��SF�RU�N��"F0�����U�F"@G�TOd�LC�H�"�%RECOV��9@�@W�`&�ӂ�H��:`_0��  }@�RTINVE��.ѡOFS��CK�KbFWD������1B,��TR�a�B �FD� ��1= B1pBL� �6� A1L�V��Kb����#��@+<�AM:��0��j��_M@ ~�@h���T$X`x ��T$HBK���F���A�����PPA�
��	����~��DVC_DB�3�@pA�A"��X1`�X3`��S�@��`�0��Uꣳ�h�CABPP
R�S #���c�B�@���GUBCPU�"��S�P�` R��11)ARŲ�!?$HW_CGpl�11� F&A1Ԡ@8p��$UNITr�|l e ATTRIr@�y"��CYC#b�C�A��FLTR_2_FI������z2bP��CHK_���SCT��F_e'F1_o,�"�*FS�Jj"CHA�Q�'91Is�82RSD����1���_Tg�`�L i�EM�NPMf�T&2 8p&2- �6�DIAGpERAI�LACNTBMw�L�O@�Q��7��PSı�� � ��PRRBSZ`�`BC4�&�	��FUN5s��RIN�PZaߠ�0�7Dh�RAH@���`�� `C�@�`C�Q�C�BLCURuH�DA0�K�!�H�HDAp�aA�H�C�ELD�������C��jA�1�CTI�BUu�8p$CE�_RIA�QJ�AF� P��>S�`DUT�2�0C��};OI<0DF_LC�H���k�LMLF�aH�RDYO���RG��@HZ0��ߠ�@�UM�ULSE�P�'3.iB$J��J�����FAN_ALM��dbWRNeHA#RD��ƽ�P��k@!2aN�r�J�_}��AUJ R+4�TO_SBR��~b�Іj�e 6?A�cMPIN�F��{!�d�A�cREG�NV��ɣZ�5D��NFLW%6r$M�@� ��f� ��0 h'uCM4NF�!�ON	 e!e�#�(b*r3F�3 �h	 ���q)5�$�g$Y�r�� u�|_��p*$ �/��EG������qAR��i���2�3�u�@<�wAXE��ROB��7RED��WR��c�_���SY`��q� :?�SI�WRI���vE STհ�ӭ d���%Eg!���t8��^a"��B����9�3� �OTO�a����ARY��ǂ�1������FIE���$LI�NK�QGTH���T_������390���XYZ����!*�OFF������ˀB��,B`l������m�FI� ���C@Iû�,B��_J$�F�����S`����3-!$1�w0��d�R��C��,�DU��r��3�P�3TUR`!XS.�Ձ�bXX�� ݗFL�d���pL��0���34���� +1)�K��M��5�5%B'��ORQ�6��fC㘴��0B�O;�D�,������aN�OVE��rM�� ���s2��s2��r1���`0���0�g /�AN=! �2�DQ�q���q�} R�*��6����s��V����ER��jA	�2E���.�C��A���0���XE�2Ӈ�A��AAX��F��A�N!�S� �1_��Q_Ɇ�^ʬ�^� ��^��0^ʙ�^ʷ�^�1&�^ƒP[ɒPkɒP {ɒP�ɒP�ɒP�ɒP �ɒP�ɒP�����ɪ ��R>�DEBU=#�$8ADc�2����
�A!B�7����V� <" 
��i�q��-! ��%��׆��׬��״� ���1�י��׷�JT���DR�m�LAB��8ݥ9 FGRO� ݒ=l� B_�1�u� ��}��`����ޥ��qa��AND�����qa� �Eq��`1��A@�� �NT$`��c�VEL�1��m���1u���QP��m�NA[w�(�CN1� ��3�줙���SERsVEc�p+ $@@�d@��!��PO�
�� _�0T !�p�𗱬p, w $TRQ�b�
(� -DR2�,+"P�0_ .� l"@!�&ERR���"I� q���~TOQ����L�p]�e���0G��%�����|	 �@ / ,��/I -��RA� �2. d�&�! 0�p$�&��2tPM� OC|�A8 1  p�COUNT�� ��qFZN_CFG�2 4B �f�"T��:#��Ӝ� x��`�s3 ���M:0�R�qC@��/�:0��FA1P��?V�X������r���� �P:b�pHEL�pe4 5���B_BAS�cRSSR�f @�S�!�QY 1�Y 2|*3�|*4|*5|*6|*72|*8�L!RO������NL�q �AB����0Z ACK��I-NT_uUS`�Pta9_PU�>b%ROU��PH@�h9#��u`w�9�TPFWD�_KAR��ar R�E���PP��A�QUE�i&��	�f�>`QaI`��9#�j3r��f�SEME��6��PA�STY4SO�0�DI'1�`���18�rQ_TM�cM�ANRQXF�EN�D�$KEYSWITCHj31:A��4HE	�BEATmM�3PE�pLE�(���HU~3F�42�S?DDO_HOM�BPO:a0EF��PARr��*�v�uC�@�O�Qo �OV_Mtϒ��Eq�OCM��d�7��p8%HK�qG5 D��g�Uj��2M�p�4R��FO�RC�cWAR���	:#OM�p 6� @�Ԣ�v`U|�P��p1�V'p�T3�V4���*#O�0L�R7<��hUNLOE0h�dEDVa  s�S�@d8 <p�AQ9�l1MSUP�G�UaCALC_�PLANcc1��A�YS1�1���@�9 '� X`��P � q;a�թ�w��2��j�M$P�㣒�fyt$��rSC�M�pm�q ����aq��0�tYzZ�zEU�Q�b�� T�!�Hr�pPv,NPXw_ASf: 0g �ADD��$S{IZ%a$VA��~�MULTIP�"�ns�PA�Q; � $T9op�B����rS��j!C~ �vF'RIF�2S�0�Y�T�pNF[DODB�UX�B��u&�!���CMtA�Е������������Z ��< �3 �p�TEg���^��$SGL��T���X�&{���㰀��S�TMTe�ЃPSE�G�2��BW���S�HOW؅�1BAN�`TPO���gᣥ��Ԣ���9`V�_Gv�= ��$PC��X�O�FB�QP\��SP�0A&0^���V�DG��>� �cA00�����P����P���P���P��5���6��7��8��9��A��b`���P��w���S`��F����h����1��v�h�י1�1��1��1�1�1�%�12�1?�1L�1�Y�1f�2��2��2���2ʙ2י2�2��2��2�2�2�%�22�2?�2L�2�Y�2f�3��3��3���3ʙ3י3�3P�����3�3%�U32�3߹3L�3Y�U3f�4��4��4��U4ʙ4י4�4�U4��4�4�4%�U42�4߹4L�4Y�U4f�5��5��5��U5ʙ5י5�5�U5��5�5�5%�U52�5߹5L�5Y�U5f�6��6��6��U6ʙ6י6��6�U6��6�6(�6%�U62�6߹6L�6Y�U6f�7��7��7��U7ʙ7י7��7�U7��7�7(�7%�U72�7߹7L�7Y��7f�ORV�`_UP�D��? �c� 
�PV���@ x $TOR�1T�  �cOP �, 6ZQ_7RE^��(� J��SsC�A���_U�p�7bY�SLOA"A � �u$�v��w�@��x�@��bVALUv�10�6�F�ID�_L[C:HI5I~�R$FILE_X3�eu4$�C7 �S;AV��B hM �?E_BLCK�3�|ȁ�D_CPU���p��p5hz�pY���R3R C � PW��� 	�!;LAށSR�#\.!'$RUN�`G@% $D!'$�@G%e!$e!�'%HR03$� '$��T�2Pa_LI�RD w � G_O�2}�0P_EDI�R�@�T2SPD�#�E�"i0ȁ�p	����DCS9@G)�F � 
$JPQC71��� S:C;}C9$MDL73$5P>9TC�`@7�UF�@?8S� ?8COBu �@�"|�L�G�P;;� 9�:;8`TAB'UI_�!L�HGb�%r�0FB3G$�3�A�sR�LLB_AwVAI�B  d�4��!��I $� SE�L� NẼ�@RG�_D N��TaOQ�3S=C�PJ �1/A�B�PT�R`�1_M]`L�K \M f/Q�L_��FMj��PG�i�U9R�6��PS�_�P\� �p�EE�7B�TBC2�eL� ���``�`b$�!FT�P'T�`
�TDCg�� BPLp�sLNU;WTH��qhT�gtWR�2$�pERVE.S�T;S�Tw��R_ACkP MX -$�Q�`.S �T;S�PU@�`IC�`7LOW�GF1�QR�2g�`��p�S�ERTIA�d^0iP��PEkDEUe�LA7CEMzCC#c��V�BrpTf�edg�aT�CV�l�adgTRQ �l�e�j|�Scc��edcBc�J7_ 4
�J!���Se@qde�Q2��0���1�PRcuPJKlvVK<�~qcQ~qw�bspJ0��q�sJJ�s;JJ�sAAL�s�p �s�p�v���r5sS�`N1�l�p�k�`5dXA�_́IDXQC�F�BN `M GRCOU ��bh�NP�C0sD�REQUI9R�R� EBU�C�Qz�6g0 2Mz�X�Pd�QSGUO�@��)APPR0C�7@� 
$� N��CLO� ǉS^U܉Se�
Q�@A�"P �$PM]P�`�`sR�_MGa!�C���+���0�@,�BRK*�N�OLD*�SHOR�TMO�!m�Z��JWA�SP�tp`�sp`�s�p`�sp`�sp`�A��7���8sQ �!�PTQ�� m��R.Qx�cQ�PATH��*� �*��X&���P�NT|@A�"p���6 �IN�RUC4`aZ��C�`UM��Y
`�)p��>�Q��cP����p��PAYLO�Ah�J2L& R_	Am@�L ������+�R_F2LS3HR�T/�LO���p0���>���ACRL0 z�p�y�ޤsRH5b�$H+���FLE�X����JVR P��_._�_�_���>�US :�_�V d`0�G��_tQd`�_�_lF1G��ũ�o0o BoTofoxo��E�o�o �o�o�o�o�o �� ��wz3lt����3EHWF�^zT!��X� ��ju��uu~�W؁ ���p�u�u�u�u������(�T ��P5�G�Y�� ' AT��l�pEL0�_B��js�J�Sz�JEW�'CTR7B`NA���d�HAND_VB�����TUO@h`+�`TSW��"�A�V� $$M��e G�AV� Qs�De�oAA��@�	$�A5�G�AU�Ad�� 6��G�UDU�Dd�PD�G/ �-STI�5V�5Ng�DYF ��+�x� ���P&�G�&�A��lw�o�Q�k�P������ ʕӕܕ��	�T�W 7 �� ���3%�?!ASYM$T��m�T�V�o�A�t�_SH�~��� ���$����Ưد�J񬢐�#39"���_VI��`8�q0V_UNIrS�4��.�Jmu�2��2A��4 X��4�6a�pt��������&E_�����!�E���CH( Xc ̱���TOc�PP�VsSvD�US�RU�P�����z@�D�A}@_5�U��P�EyA�a��RPROG_N�A��$�$LAsST���CANs��ISz@XYZ_SP�u�DW]R@Ͱ,VS�V@�E1QENc��DC�UR�H�P��HR_�T��YtQ9S�d��O�T��uP?�Z ��I�!A �D���Q���#�S�������3�vP [ �[ ME�O�h�R#B�!T�PPT0 F@1�a��̰� �h1a%iT0� �$DUMMY1���$PS_��RMF��  1�lfװ7FLA*�YP�b�c$GLB_T�I �U�e`gA��LIF(!\����g`�OW�P��eVOL2#qb �a_2��[d2�[`����b�P�c�Z`TC��$BA�UDv��cST��B|�2g`ARITY0soD_WAItAIyYCJ2�OU6�Zq>yyTLANS�`�{�S�SZc��BUF�_�r�fиx�PyyCwHK_�@CES���� JO`E�axA�x�bUBYT�� ���r�.�.� ��aA��M�������Q�] Xʰ����ST�����SBR@M�21_@��T$S�V_ER�b����C)L�`��A1�O�BpP�GLh0EW(!^ o4 $a$Uq;$�q$W�9���A�@R����ՁU�م_ "��D$�GI��}$ف �^҄�(!` qL�.��"}$F�"=E6�NEAR��B'$F}��TQ���PJ�@R� a��$JOINT�a�)�ӃMSE]T(!b  +�Ec��2�^�Se�G�_�(!c��  ��U�?����LOCK_F�O@� �PBGLV���GL'�TE�@X9M���EMP����qK��b�$U��؂a�2_���q�`�<� �q�^��CE�/�?��� $KAR�b�M�STPDRA8܀����VECX���֪�IUq�av�HE��TOOL���Vv��REǠIS3�2�6��ACH̐m Mb^QONe[d3����IdB�`@$RAIL_BOXEa���ROB�@D�?����HOWWAR�0Aa�i`-�ROLM tb��$�*���T��`��n��O_FU�!��HTML58QS��@ e�"Հ�(!d��G  ��@�(!e���������І}p(!f t��m�^a��t��B�PO��AIPE�N���O�����q��AORDED0�m �z�XT`��A�)MBPMO�P �g D �`OB �����ǯ�Uc�`���� ��SYS��AD�R��pP`U@^  �h ,"��f$A���E��E�TP�VWVA�Qi Ǥ �@ق�UPR|�B�$EDI�A�d�VSHWRU��z���IS�Uq�pN�D�P7���G�HEA�D�! @���!i�K�EUqO`CP)P��J�MP��L�U�PRA[CE�Tj����IL�S��C��NEx���TICK�ʓ!MKQ�Q��HNr�k @���HW�C��PHVF��`STYYeB+�LO�a�b(��[�C�l3�
�@�FS%$A��D=��S�!$�1�p a�e�qr�ePv HVSQU���#LO�b_1TER�C`���TS?�m 5���R�m@3����ܡ�O`	c IZ�d�A�eha�qtb�}�hA}pP~r��_D)O�B�X�pSSQ�S'AXI�q��v�bS��U�@TL���RE3Q_ܠ��ET���`��CY%��FY'��A,f\!\d9x�P� g�SR$$nl-�w �����c
�uV
Qh(�AA���dC`�A�@�	�Y��D���p�E"�	CC�C`��/�/�/	4� ��SC�` o h�5�DSmడ[`SPL�@�AT� 
R��xL��XbADDR�s3$Hp� IF�Ch�O_2CH���pO��\��- �TUk�Ir7 p��CUCp*F�V��I�Rq�4�(��c��
K�
h@]!����Pr \z�D�� ��|,K� P�"CN���*CƮ��!�TX_SCREE��s�Pp@�INA˃<�4��Dg�����`t Tᫀ�b����O Y6`���º�U4h�RR��������R1�TMAUE���u �j �qz`S�́��RSML��U`����V�1tPS_���6\��1�9G\���C8��2@4 2��0�Ov�R��&F�AM_TN_FL*�`Q���W� ��BBL�_/�WB`�Pw �ԫ��BO ��BLE�"�Cg�R"�DRIG�HtRD��!CKGRB`�ET���G�AWIDTHs���R�B��a�r<@I��EYհRx d�ʰ�����`y�BACKЍ�tb>U���PFO܉�QWLAB�?(��PI��$UR�m�~P�PP�PHy1 y 8 $�PCT_��,"�R�PRUp@�s5�da�`�QO%!Jt�zV�ȇ�pU�@r�SR ���LUM�S�� ERVJ�h�P�P��T{ � " GE�Rh� �¯ГLPAeE��)�^g�lh�lh�ki5
ik6ik7ikpP`� Z�x����$u1��p��Q zQUS=Rل| <z��P1U2�a#2�FOO 2�PRI*m9�[�@p�TRIPK�m�oUNDO��})���Yp��y���'`i����p ~�Rp�qG ��T���-!&�rOS2��vR��2�s�CA�����r�`�R_�sUIaCA�����3Ib_�sOF�FA�D@���O�b�r�5�L�t��GU��Ps������n+QSUB`� ��_E_EXE��V
�v�sWO� �#��w��WAl�p΁�fP
 V_DB���҃RT�pO�0V░���3OR/�5�'RAUa 6�TK����__���� |�j �OWNj�34�$SRC�0`���DxA���_MPFI�����ESP��T�$0 ��c��g��qq�zЎE!� `%�ۂ34�J���COP��$`��p_���/�+�6���CT�Cہ�ہ����DCS��P;4�COMp�@�;��O`�=����K�^�/�VT��q'���Y٤Z���2���@p�w#SAB����2�\0˰_��qM��%!]�DIC#池AY�3G�PEE2�@T�QS�VR1���"eQL�� a��P� D ��f�z��f�> ����6�xAA�t�b# ��L2SHADOW���#ʱ_UNSC�Ad�׳OWD�˰D�GDE#LEGAyC)�q'�VC\ }C��� v����だm�RF07����7d`C2`7�DRI%Vo���ϠC�A]��(�` ���MY_UBY�d?Ĳ��s��1@��$0�����_ఴ����L��BM�A�$�DEY	�EXXp@C�/�MU��X���,��0US����;p_�R"1�0p#�2�G>PACIN*���RG��c�y�:�y��sy�C/�RE�R"!�q��y�D@� L !�G�P�"��Tp�R�pD@�&P�Px1dQ��	.���RE���SWq�_Ar�u@$+�{�Oq�AA/�3��hEZ�U���� Y�p�HK���P�J��_/�Q0{�EAN��ۀ2�2����MRCVCA� ��:`ORG��Q�dR	p��L�����REFoG �����!�+`	�p ��������<���q�A_����r��� S�`�C��Ú�W��@D� ��0�!��#q�š��OU����?� ��Վ2�J@0� 1�*p����0� UL�@��C�O�0)��� NT�[��Z�Qf�af% L飏��Q|��a�VIAچ7� �ÀHD7 6P�$JO�`oB?�$Z_UPo��2Z_LOW��$�QiBn��1$EP �s�y�� 1!f� � 1¦4�� 5�PA�A ��CACH&�LO �w�В�1B����Cn�I#F^��T8m����$HO2�32!{��Uÿ2O�@����Ro��=a��ƐV�P��X@A"_SIZ&�K$Z$�F(�G'��v�CMPk*FAIo�5G��AD�)/��MRE���"P'GP��0е�9�ASYNwBUFǧRTD�%��$P!�COLE_2D_4�5W�sw�~��UӍQO��%EC;CU��VEM��v<]2�VIRC�!5�#�2�!_>�*&�pWp���AG	9R�XYZ@�3�W���8���4+Qz0T"��IM�16�2`�GRA�BB�q��;�LERrD�C ;�F_D��F�f50MH�PE�R�Z��� ��KQL�AS�@��[_GEb� �H൑~23�ET����"���b���I�D�ҙ6m�BG_gLEVnQ{�PK|�X�6\q��GI�@N\P�4���P��!g��dr�S� �NRT
'�VLʁc�Ų���#a��c"!D�qDE�����Xа�X��P�Җ1��d��pzZP���d�c���D4q_���2pT���U&�� $�IT�Pr9p[Q��ՓV�VsSF$�d�  fp�/�f�UR&�  �R`MZu�dr��AcDJ`C�� ZDVfg� D�XAL� x� 4 PERIKB$MSG_Q3$Q!o%[���p'���dr:g�qQ� ��XVR\t��B�pT�_\��R_�ZAB�C"����Sr���
|W��aACTVS'� � � $x|u�0�cCTIV�Q�!IOu¥s&D�I�T�x�DVϐ
Hx�P���!���pPS���� �#��!8���q!LSTD�!ع  �_ST����aq�CHx�� L-�@��u�Ɛ*���P GNA#�C�<!q�_FUN��  ��ZIPu�3�HR�$L���}XZMPCF"���`bƀ�rX�ف��L�NK��
Ă�0#�� $ !��ބ�CMCMk�C8�C�"����P{q '$J8�2�D6!>� O�H���T���2������M���UX�1݅UXE1Ѡ��1C���Y���ੑ����˗7�FTFpG>�����C�Z���� �k�� �"8�YD'@ �� 8n�R� U�ӱ$HEIGH�d�:h?(! 'v���@���� � Gd��qp$B% � E���SHIF��hR�Vn�F�`�HpC � 3�(�8H`O�ѡ�ȭC��+%D	�"�CE�pV�1
�SPH�ERs� � ,�! M�c�u��$P�OWERFL  )�p|����|�p��RG�`  �������/A�  ��?�p����pd��NSb ����?_�  Bz|� l�_  <@�|��%���˃���涜ŵ�� 2ӷ�� W	H��l&����>���A �|��t$��*z��/�� **:�� �p�ϥ��͘�����#����ɘ��|� ����5�������%� ��I�[߉�ߑ��� ��������w�!�3�a� W�i����������� O����9�/�A���e� w�������'���� �=O}s� ������k 'UK]���� ��C/��-/#/5/ �/Y/k/�/�/�/?�/ �/?�/?�?1?C?q? g?y?�?�?�?�?�?�?�_O	OOIO?OQO�� 	 �O�O�O_�E ��3_���O`_�O�_�_�÷PREF �Ӻ�p�p
��IORITY a|���2�p����pSPL`z�����WUT�VqÈ�O�DU~����,�_?�OG��Gx��R\��,fHIBqOy��|kTOENT 1���yP(!AF�_b�`�o�g!�tcp�o}!�ud�o)~!iccm�0bXY̳��k �|�)�a �����p�� ��u������ N�5�r�Y�������̏H�����*/c̳ӹ����E�W�|�>�U�F��/��4����|��,�7�A��,/  ��P���P�%�|�'���Z���h�z�����|��E�NHANCE )	#�7�A9�d������  �,f�T
�_�S����POR�Te�rb�@�U���_CARTRE�P�Pr|brSKSTyAg�kSLGS�`��k����@U�nothing ������Ϳ>�P��b�To��TEMP �?isϨE/�_�a_seiban m_��i_�����0�� T�?�x�cߜ߇ߙ��� ��������>�)�N� t�_��������� ����:�%�^�I��� m����������� �� $H3lWi� ������ D/hS�w����uϪ�VERSI��P=g  d?isable��SAVE ?j�	2670H7K05��k/!�0m//*�/ 	�(%b$�O�+�/�Se?6?H?Z?l?z:%<�/�?t4�*'_j` 1�kX �0ubuE�?O�qG�PURGE��Bp`�ncqWF<@�a�T�Ӓ*fW�`]Daa�W�RUP_DELA�Y z�f�B_?HOT %?e'b���OnER_NORMAL�HGb�O%_�GSEMI_*_i_�Q_QSKIP�3.��3x��_��_�_�_ �]?eo+goKo]ooo 5o�o�o�o�o�o�o�o �o5GYi� }������� 1�C�U��y�g����� ����я����-�?��7%�$RACFG� �[ќ�3�~]�_PARAM�Q�3y��S @Иs@`�G�42C۠5��2��CbFB�=B]�BTIF���J~]�CVTMOU������]�DCR��3�Y ���Q@��uC��1BEH@����?�y<;��]�	���;�5��l���V���_��o;e��m���KZ;��=g;�4�<�<���f@����� �5�G�Y�k�}� ������ſ׿���xU�RDIO_TYP�E  �V�5��E�DPROT_a��&>��4BHbbCEސSǆQ2c�7 ��B�ꐪ� ����ϐ����&�� ��W�V_~�o����� ����������A�O� m�r���9����� ���������=�_�d� �������������� ��'I�Nm�� ������� #EJi+k� �����//4/ F//g//�/y/�/�/ �/�/�/	?+/0?O/? c?Q?�?u?�?�?�?�?��??;?,O��S�INOT 2�I���l�G;� jO|K���<�O�f�0 �O�K �?�O�?___N_<_ r_X_�_�_�_�_�_�_ �_�_&ooJo8ono�o fo�o�o�o�o�o�o�o "F4j|b� ���������B�O�EFPOS1� 1"�  xO��o×O���� ݏ鈃���Ϗ0��T� �x����7���ҟm� �������>�P���� 7�������W��{�� ���:�կ^������ ����S�e��� ��$� ��H��l��iϢ�=� ��a��υ�� ߻��� �h�Sߌ�'߰�K��� o���
��.���R��� v��#�5�o������ �����<���9�r�� ��1���U��������� ��8#\���� ?��u��"� FX�?��� _��/�	/B/� f//�/%/�/�/[/m/ �/?�/,?�/P?�/t? ?q?�?E?�?i?�?�? O(O�?�?OpO[O�O /O�OSO�OwO�O_�O 6_�OZ_�O~_�_+_=_ w_�_�_�_�_ o�_Do��_Aozocf�2 1r�o.oho�o�o
 o.�oR�oO�# �G�k���� �N�9�r����1��� U����������8�ӏ \���	��U�����ڟ u�����"����X�� |����;�į_�q��� ���	�B�ݯf���� %�����[���ϣ� ,�ǿٿ�%φ�qϪ� E���i��ύ���(��� L���p�ߔ�/�A�S� ��������6���Z� ��W��+��O���s� �������V�A�z� ���9���]������� ��@��d��# ]���}�* �'`���C �gy��&//J/ �n/	/�/-/�/�/c/ �/�/?�/4?�/�/�/ -?�?y?�?M?�?q?�? �?�?0O�?TO�?xOOx�O�o�d3 1�o IO[O�O_�O7_=O[_ �O__|_�_P_�_t_ �_�_!o�_�_�_o{o fo�o:o�o^o�o�o�o �oA�oe �$ 6H�����+� �O��L��� ���D� ͏h�񏌏�����K� 6�o�
���.���R��� ퟈����5�ПY��� ��R�����ׯr��� ������U��y�� ��8���\�n������ �?�ڿc�����"τ� ��X���|�ߠ�)��� ����"߃�nߧ�B��� f��ߊ���%���I��� m���,�>�P���� �����3���W���T� ��(���L���p����� ������S>w� 6�Z���� =�a� Z� ��z/�'/�$/ ]/��//�/@/�/�O�D4 1�Ov/�/ �/@?+?d?j/�?#?�? G?�?�?}?O�?*O�? NO�?�?OGO�O�O�O gO�O�O_�O_J_�O n_	_�_-_�_Q_c_u_ �_o�_4o�_Xo�_|o oyo�oMo�oqo�o�o �o�o�oxc� 7�[���� >��b����!�3�E� ���ˏ���(�ÏL� �I������A�ʟe� ������H�3�l� ���+���O���ꯅ� ���2�ͯV���� O�����Կo������ ���R��v�Ϛ�5� ��Y�k�}Ϸ���<� ��`��τ�߁ߺ�U� ��y���&������� ��k��?���c��� ����"���F���j�� ��)�;�M������� ��0��T��Q�%��I�m��/�$5 1�/���m X���P�t� /�3/�W/�{// (/:/t/�/�/�/�/? �/A?�/>?w??�?6? �?Z?�?~?�?�?�?=O (OaO�?�O O�ODO�O �OzO_�O'_�OK_�O �O
_D_�_�_�_d_�_ �_o�_oGo�_koo �o*o�oNo`oro�o �o1�oU�oyv �J�n���� ���u�`���4��� X��|�ޏ���;�֏ _������0�B�|�ݟ ȟ���%���I��F� ����>�ǯb�믆� �����E�0�i���� (���L���翂�Ϧ� /�ʿS�� ��Lϭ� ����l��ϐ�ߴ�� O���s�ߗ�2߻�V� h�zߴ�� �9���]� �߁��~��R���v�����#�	6 1&����������� ����}���<�� `����CUg ��&�J�n 	k�?�c�� /���	/j/U/�/ )/�/M/�/q/�/?�/ 0?�/T?�/x??%?7? q?�?�?�?�?O�?>O �?;OtOO�O3O�OWO �O{O�O�O�O:_%_^_ �O�__�_A_�_�_w_  o�_$o�_Ho�_�_o Ao�o�o�oao�o�o �oD�oh�' �K]o�
��.� �R��v��s���G� Џk�􏏏���ŏ׏ �r�]���1���U�ޟ y�۟���8�ӟ\��� ���-�?�y�گů�� ��"���F��C�|�� ��;�Ŀ_�迃����� �B�-�f�ϊ�%Ϯ� Iϫ����ߣ�,���xP�6�H�7 1S� ���I��߲������ ��3���0�i���(� ��L���p�����/� �S���w����6��� ��l�������=�� ����6���V� z� 9�]� ��@Rd�� �#/�G/�k//h/ �/</�/`/�/�/?�/ �/�/?g?R?�?&?�? J?�?n?�?	O�?-O�? QO�?uOO"O4OnO�O �O�O�O_�O;_�O8_ q__�_0_�_T_�_x_ �_�_�_7o"o[o�_o o�o>o�o�oto�o�o !�oE�o�o>� ��^����� A��e� ���$���H� Z�l�����+�ƏO� �s��p���D�͟h� 񟌟���ԟ�o� Z���.���R�ۯv�د ���5�ЯY���}�c�u�8 1��*�<� v���߿��<�׿`� ��]ϖ�1Ϻ�U���y� ߝϯ�����\�G߀� ߤ�?���c����ߙ� "��F���j���)� c����������0� ��-�f����%���I� ��m������,P ��t�3��i ���:��� 3��S�w / ��6/�Z/�~// �/=/O/a/�/�/�/ ? �/D?�/h??e?�?9? �?]?�?�?
O�?�?�? OdOOO�O#O�OGO�O kO�O_�O*_�ON_�O r___1_k_�_�_�_ �_o�_8o�_5ono	o �o-o�oQo�ouo�o�o �o4X�o|� ;��q���� B����;������� [�������>�ُ�b�����!�������M�ASK 1 ��⤒���ΗXNO�  ݟ���MO�TE  ���S�_?CFG !Z����N�����PL_RGANGV�N������OWER "���Ϡ��SM_DRYPRG %����%W��եTAR�T #Ǯ�UME_PRO���q����_EXEC_E�NB  ����G�SPDJ�����Ρ�TDB����RM�п��IA_OPTgION��������NGVERS���`�řI_AIRPUR��� R�+���ÛMTE_֐T X���ΐ�OBOT_ISO�LC��������^��NAME8��H��ĚOB_CATEG�ϣ,��S�[��.�ORD_NUM� ?Ǩ���H705  �N��ߨߺ�ΐPC_TIMEOUT��{ xΐS232s��1$��� L�TEACH PENDAN��o����)��V�T��Maintena�nce Cons�N�&�M�"B�P�?No Use6�r� 8��������̒��GNPO$��Ҏ�"Ž��CH_LM��Q���	a�,�!OUD1:��.�RՐ�VAILw���|��*�SR  t�� ���5�R_I�NTVAL��� ���V_DA�TA_GRP 2�'���� D��P�������	� �����B 0RTf���� ��/�/>/,/b/ P/�/t/�/�/�/�/�/ ?�/(??L?:?p?^? �?�?�?�?�?�?�?O  O"O$O6OlOZO�O~O �O�O�O�O�O_�O2_  _V_D_z_h_�_�_�_ �_�_�_�_o
o@o.o�Povodo�o��$S�AF_DO_PU�LSW�[�S���i�S'CAN��������SCà(�����+S�S�
����P��q�q�qN� � L^p���5���� ��$���+��r2M�qqd�Y�P�`�J�	t/� @��������ʋ|�� r ք��_ @N�T ��'��9�K�X�T D��X���������ɟ۟ ����#�5�G�Y�k��}�������䅎������Ǧ  ="�;�oR� ����p"�
�u��Di���q$q�?  � ���u q%�\�������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$�6�H�Z����珈�� �����������g� ;�D�V�h�z�������@��������(�Ӣ0� r�i�y���$�7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/?r�+? =?O?a?s?�?�?�?�? �?8��?OO'O9OKO ]OoO�O��$�r�O �O�O�O	__-_?_Q_ c_u_�_�Y�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|�c�路g����� ��0�B�T�f�x����������ҏ����p��:�Ҧ��y��3�	�	123�45678��h�!B!�� +\��p0�� ��Ο�����(�:� @��c�u��������� ϯ����)�;�M� _�q�����R���ɿۿ ����#�5�G�Y�k� }Ϗϡϳ����ϖ��� ��1�C�U�g�yߋ� �߯���������	�� -���Q�c�u���� ����������)�;� M�_�q���B������ ����%7I[ m������� �!3EWi{ �������/ ///�S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?D/�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O*����O	_�E�?5_�G_Y_�yCz  �A��z   ���x2�r }��)�
�W_�  	�*�2�O �_�_ oo"l�#\��_hozo�o�o�o�o �o�o�o
.@R dv����Mo� ���*�<�N�`�r� ��������̏ޏ��� �&�8�J��X #P$Pt�Q�R<u� k�~�Q  �������S�P���Q�Qt�  �PÙ۟�P(� `,b����]��PFl�$SCR_�GRP 1*�+4� �� �,a ��U	 v��~������ d���%���ɯ���h]���P�D1� D7n��3��Fl�
CRX-10�iA/L 234�567890�P�d� r��Pd�L ��,a
1o�����Z���[ ¶~� +fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@��R�d�t���H�~�Ă�m��ϴ�8����,a@�N�����,a��1���U�[��G�imXhuP,[~��V��B�  B!ƠߞҷԚ�A�P��0�����Ԛ�@�����' ?���H�����ښ�F@ F�`A�I�@�m�X��|� �������������р���:�%�7�I�[�B�i������������ ����-Q<u` ��En�ٯ���W�P�"��_�5��h1`b���x�� ��ͣ�O�,dA���H����Fa�,a �#!"/4/E-�!Z(f/x/G/ 	(�P�!(� �/�/�/ ��/�/?#9b�����S7س�M�ECL�VL  ,a���ݲ�Q@f1L_DEFAULTn4�b1�1`~�3HOTSTR�=���2MIPOWEKRFm0pU�5�4oWFDO�6 �5�L�ERVENT �1+u1u1�3 L�!DUM_EI�P#?5H�j!AF_INE�0SO,dO!FT)O�NIOr�O!���O ��O��O!RPC_M'AIN�O�H��O>_NSVIS_�I�-_~�_!OPCUf̦_�Wy_�_!�TP�PPU�_<Id��_"o!
PMON?_PROXY#o?FAeono�R<o8Mf]o��o!RDM_S�R���oADg�o!#R��"=Hh�oRK!
PM�o9LiA��!RLSYN�C��y8��!�ROS(O��4��6�!
CE�PMOTCOM7�?Fk%����!	K�CONSd��>Glq�Ώ!K��WASRC�o?Fm콏�!K�USB��=Hn	�f�!S#TM�0��;JoU�����O֟�c����CICE_KL ?%K� (%SVC�PRG1��G�1�2�G�L�6�3o�t�6�4�����6�5��į6�6��6�7��6���$;�5�9_�d�3� ��6�9���6�a�ܿ6� ���6���,�6�ٯT� 6��|�6�)���6�Q� ��6�y���^����^� ʿD�^��l�^�ϔ� ^�Bϼ�^�j���^��� �^���4�^���\�^� 
߄2���6�� /����V��<�'�`� K���o����������� ��&J5nY ������� �4F1jU�y �����/�0/ /T/?/x/c/�/�/�/ �/�/�/�/??>?)?�P?t?_?�?
�_DE�V I��MC:�84��~�4GRP 2/E��0+�bx 	_� 
 ,@�0�?OD8OJO1OnO UO�O�O�O�O�O�O�O �O"_	_F_-_j_|_c_ �_�[O�_�_�_o�_ ,ooPo7oIo�omo�o �o�o�o�o�o(:8!^�_  �1i @�������  �=�$�a�s�Z���~� �������؏�l
� K���qp�W��Q��� 	�Ο�����(�� L�3�E���i�����ʯ ܯ�_ ��ɯ6��Z� A�~���w�����ؿ� ѿ���2�D�+�h�O� ��s�9���]����ϳ� �ߙ�'��v�]ߚ� �߾��߷������*� �N��r��;��� ���������&�8�� \�C���g�y������� ����g�4-j Q�u����� B)fx_ ����)��/ ,//P/7/t/[/m/�/ �/�/�/�/?�/(??�L?^?E?�?�7d ��[~
�6 s� 	 A;*�=� 6?�=����D�>�����g�:�0���ī��|@��-�@�5_�e�A5�-�=B�G+h�&����6)AB�m����`x��=��?7O%TELE�OP8OcN[~y���5�o�ʾT�F�����������|��?ҝ����E�1��E@�*��A`�~�n�!���$�A����M�Y<T�������C=��J����Gc��McO��IJO/_��[~��6r �_�1<�׻���y;��	A`��ʛ1bP��N	V��A�&@в�@���@)E��]�1������0ד� x����Q��U?�Q��O�__ _o DS�I�I2o oVoDozoho�o�o%�o�o�_ �o�o0TBx �o��oh�d�� �,��P��w��@� ����Ώ��ޏ��(� j�O������p����� ʟ��ڟ �B�'�f�� Z�H�~�l�����Ư� �����د�� �V�D� z�h����ſ����� ��
��R�@�vϸ� ��ܿf��Ͼ������ ��Nߐ�uߴ�>ߨ� ���ߺ����� �V�|� M��&��n����� ����.��R���F��� V�|�j���������� *���B0Rx f������� >,Nt�� �d����// :/|a/s/*/L/&/�/ �/�/�/�/?T/9?x/ ?l?Z?|?~?�?�?�? �?,?OP?�?DO2OhO VOxOzO�O�OO�O(O �O_
_@_._d_R_t_ �O�O�_ _�_�_�_o o<o*o`o�_�o�_Po �oLo�o�o�o8 zo_�o(���� ����R7�v � j�X���|������ *��N�؏B�0�f�T� ��x�����՟矞��� ���>�,�b�P���ȟ ���v��ί��� :�(�^�����įN��� ��ܿʿ�� �6�x� ]Ϝ�&ϐ�~ϴϢ��� ����>�d�5�t��h� Vߌ�z߰ߞ������ :���.���>�d�R�� v����������� *��:�`�N������ ��t�������& 6\�����L�� ����"dI[ 4|���� �<!/`�T/B/d/ f/x/�/�/�//�/8/ �/,??P?>?`?b?t? �?�/�??�?O�?(O OLO:O\O�?�?�O�? �O�O�O _�O$__H_ �Oo_�O8_�_4_�_�_ �_�_�_ ob_Go�_o zoho�o�o�o�o�o�o :o^o�oR@vd �����6� *��N�<�r�`���� ��Ϗ��������&�� J�8�n�����ԏ^�ȟ ��؟ڟ�"��F��� m���6�����į��ԯ ֯��`�E����x� f���������п&�L� �\���P�>�t�bϘ� �ϼ�����"Ϭ�ߨ� &�L�:�p�^ߔ��ϻ� �τ������ �"�H� 6�l�ߓ���\���� ��������D���k� ��4������������� 
L�1C����d �����$	H �<*LN`�� ��� �//8/ &/H/J/\/�/��/� �/�/�/?�/4?"?D? �/�/�?�/j?�?�?�? �?O�?0Or?WO�? O �OO�O�O�O�O�O_ JO/_nO�Ob_P_�_t_ �_�_�_�_"_oF_�_ :o(o^oLo�opo�o�o �_�oo�o 6$ ZH~�o��n� j���2� �V�� }��F�������ԏ 
���.�p�U������ v���������П�H� -�l���`�N���r��� �����4��D�ޯ8� &�\�J���n����˿ 
��������4�"�X� F�|Ͼ����l����� ����
�0��Tߖ�{� ��D߮ߜ��������� �,�n�S����t� ��������4��+� �����L���p����� �����0���$4 6H~l���� ��� 02D z���j��� �/
/,/��y/� R/�/�/�/�/�/�/? Z/??~/?r??�?�? �?�?�?�?2?OV?�? JO8OnO\O~O�O�O�O 
O�O.O�O"__F_4_ j_X_z_�_�O�__�_ �_�_ooBo0ofo�_ �o�oVoxoRo�o�o�o >�oe�o.� �������X =�|�p�^������� �����0��T�ޏH� 6�l�Z���~������ �,�Ɵ ��D�2�h� V���Ο���|��x� ���
�@�.�d����� ʯT������п�� �<�~�cϢ�,ϖτ� �Ϩ��������V�;� z��n�\ߒ߀߶ߤ� �����������4� j�X��|������� �������0�f�T� �������z����� ��,b����� R����� j�a�:��� ��� /B'/f� Z/�j/�/~/�/�/�/ /�/>/�/2? ?V?D? f?�?z?�?�/�??�? 
O�?.OORO@ObO�O �?�O�?xO�O�O_�O *__N_�Ou_�_>_`_ :_�_�_�_o�_&oh_�Mo�_�P�$SE�RV_MAIL + �U�`��Qvd�OUTPUT�h��P@vdRoV 20f  �`� (a\o�ovdS�AVE�l�iTOP�10 21�i d 6 s�P6r _�a2oX j|������ ���0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(��:�guYP�cF�ZN_CFG 2e�c�T�a��e|�GRP 23���q ,B  � AƠ�QD;� �BǠ�  B4~�SRB21�foHELL�4e�v�`�o��/�>�%RSR>�?�Q��� u�����ҿ������ ,��P�;�t�_Ϙϩ�-���s`�¼�P���Ϸͻ��P�L&�'�ސW��2�P�d��g��HK ;15�� ,ߡ� �ߥ���������@� ;�M�_���������������OMM �6��?��FTOV_ENB�d�au��OW_REG_�UI_��bIMIO/FWDL*�7.�ɥ^��WAIT\�`ِ�����`���d��T�IM������V�A�`����_UNI�T[�*yLCy�T�RY��uv`ME�8���aw֑d ���9� ������<��X�Pڠ6p`?�  ���o+=�`VL�l�fM�ON_ALIAS� ?e.��`he Go������/ )/;/M/�q/�/�/�/ �/d/�/�/??%?�/ I?[?m??�?<?�?�? �?�?�?�?!O3OEOWO O{O�O�O�O�OnO�O �O__/_�OS_e_w_ �_�_F_�_�_�_�_�_ o+o=oOoaoo�o�o �o�o�oxo�o' 9�o]o��>� �����#�5�G� Y�k��������ŏ׏ ������1�C��g� y�����H���ӟ��� 	���-�?�Q�c�u� � ������ϯᯌ��� )�;��L�q������� R�˿ݿ��Ͼ�7� I�[�m��*ϣϵ��� ���ϖ��!�3�E��� i�{ߍߟ߱�\����� ������A�S�e�w� ��4���������� �+�=�O���s����� ����f�����' ��K]o��>� ����#5G Y}����l��$SMON_D�EFPROG �&����� &*SYSTEM*����RECALL ?�}� ( �}�tpconn �1=>192.1�68.56.1:�22712 *.*S/e d!�/�/�/�,�}xyzrate 1R/d"�/}/?� ?2?�"8copy� frs:ord�erfil.da�t virt:\�tmpback\`�/?�?�?�?}/K2mdb:h `?r?{?�OO0O�$3xK4:\�?h/b#�?�O�O�O
� 4KEaSOeO�/	__-_�'
�'g!�O�O �O�_�_�_�/m_�/{_ oo0oC?U?�?y?�o �o�o�?�?no�? ,?OQOd_uO��� �O�O`�_��(�;_ M_��7������_�_ �_o����$�6�I�� ���������ԏf� x�	��-�@�R���� ��������Пb�t�� �)�<�N��򯃿�� ����̯^�p����%� ��J�ܿX� ϑϣϵ�|ȿX'15124i��{���0���J disc 0��������P�ߝ߯���K$0U� b�t���)�<oNo�o �߃���o�og��� {���0�C��h��� ��������X�j��� ��#5H���������������[$880��j|1��K������ ���U�bt//)/ <N����/�/�/����716��z/?0?/?B��/6 �/�/ �?�?�?�T?f?x?	O O-O@/R-�?�?�O�O �O�/�/�/rO__'_:�L�^��O67_�_�_ ����f_�I{_oo0o�CS�$SNPX_�ASG 2:����Va�o  0DQ%�7o�~o  ?�GfPA�RAM ;Ve�`a �	lkP�>TDP>X�d�� ��I`OFT�_KB_CFG � CS\eFcOPI�N_SIM  
Vk�b+=OYs�I`RVNORDY?_DO  �eu�krQSTP_D�SB~�b�>kS�R <Vi �{ &c`ELEO�e��>U>TW`I`TO�P_ON_ERR�xGb�PTN �VeP��D�:�RING_PR�M'��rVCNT_�GP 2=Ve�ac`x 	���DP���я����BgVD�ROP 1>�i�`� Vq؏0�B�T�f�x��� ������ҟ����� ,�>�e�b�t������� ��ί���+�(�:� L�^�p���������ʿ �� ��$�6�H�Z� l�~ϐϷϴ������� ��� �2�D�V�}�z� �ߞ߰���������
� �C�@�R�d�v��� �������	���*� <�N�`�r��������� ������&8J \n������ ��"4[Xj |������� !//0/B/T/f/x/�/ �/�/�/�/�/�/?? ,?>?P?b?t?�?�?�?��?�?�?�?O�PRG_COUNT�fs�P�)IENBe��+EMUC�dbO_UP�D 1?�{T  
ODR�O�O�O�O �O__A_<_N_`_�_ �_�_�_�_�_�_�_o o&o8oao\ono�o�o �o�o�o�o�o�o9 4FX�|��� ������0�Y� T�f�x���������� ����1�,�>�P�y� t���������Ο��	� ��(�Q�L�^�p��� �������ܯ� �)� $�6�H�q�l�~����� ��ƿؿ���� �I��D�V�"L_INFO� 1@�E�@��	 yϽϨ������@6Β����>�л����>�
�����Q*sB|Ӵ���|-A�V8���A������������h� �C�ײ�&���úם�3��@����| ��p߂�-@YSDEBSUG:@�@�o�d�I���SP_PASS�:EB?��LOG� A���A  �o�i�v�  ��Ao�UD1:�\��}���_MPC �ݚEk�}�A&��� �AK�SAV �B��IA���*�i��1�SVB�TEM�_TIME 1C����@ 0A@�=D�{Eo�Y��*����MEMBK  �EA��������X|�@� @��n����������dh�9
�� ��@�`r��������� � @Rdv�����
Le�//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H?Z?��SKV�[�EAj���?�?�?��.o���]2���?i�  0 o�^
:O.@�R�O�O�O}N��B� ��OB��F__p/_#S_D2�Y_@�_�_�_�_�_o�$�_ �_�o'o9oKo]ooo �o�o�o�o�o�o�o�o�#5GYk_?T�1SVGUNSP]D�� '����p�2MODE_LI�M D��Ҋt2̗p�qE�݉uAB�UI_DCS 	H}5���0�G�-���C��|-�X�>���*7���� 
��e��i���r�B������uEDIT �I��xSCRN �J���rS�G 3K�-� �0߅�SK_OPTIO�N��^����_DI~��ENB  ,�����BC2_GR/P 2L������MPC�ʓ�|BC�CF/�N���� 8=����`�>� W�B�g���x�����կ ��������S�>� w�b���������Ͽ�� ���=�(�a�Lυ� ��Ň�϶�������v� �
�/�U�@�yߧ�� `�iМ��߰�����
� ��.��>�@�R��v� �����������*� �N�<�r�`������� ��������̀4 FX��|j��� ����B0 fTvx���� �/�,//</b/P/ �/t/�/�/�/�/�/�/ �/(??L?d?v?�? �?�?6?�?�?�?O O 6OHOZO(O~OlO�O�O �O�O�O�O�O __D_ 2_h_V_�_z_�_�_�_ �_�_
o�_.oo>o@o Ro�ovo�ob?�o�o�o �o<*Lr` �������� &��6�8�J���n��� ��ȏ���ڏ��"�� F�4�j�X���|����� ���֟��o$�6�T� f�x���������ү�� �����>�,�b�P� ��t��������ο� �(��L�:�\ς�p� �ϔ��ϸ������� � �H�6�l�"��ߖߴ� ����V������2� � V�h�z�H������ ��������
�@�.�d� R���v����������� ��*N<^` r������� &8�\Jl�� ������"// F/4/V/X/j/�/�/�/ �/�/�/?�/?B?0? f?T?�?x?�?�?�?�? �?O�?,O�DOVOtO �O�OO�O�O�O�O�O�_ V4P�$TBC�SG_GRP 2�O U� � �4Q 
 ?�  __q_[_�_ _�_�_�_�_�_o%k�8R?SQF\d��HTa?4Q	 H�A���#e>����>$a�\#eAT��A WR�o�h|djma�G�?Lfgr�bp�o�n�ffhfG��ͼb4P|j��o�*}@��Rhf�ff>�33pa#e<q!B�o+=xrRp�qrUy�rt~��H�y0 rIpTv�pBȺt~ 	xf	x(�;���f����N�`���ˏڋ�����	V3.00~WR	crxlڃ	*��3R~t2��HH��� \�.�n]�  cC.�X����8QJ2?SRF]�����CFG -T UPQ SPܚ+��r�ܟ1��1�W�e�	Pe� ��v�����ӯ����� ���Q�<�u�`��� ������Ϳ�޿�� ;�&�_�Jσ�nπϹ� ��������WRq@� 0�B���u�`߅߫ߖ� �ߺ������)�;�M� �q�\������4Q  _���O ���J�8� n�\������������� ����4"XFh j|������ .TBxf� �nO����// >/,/b/P/�/t/�/�/ �/�/�/�/�/?:?(? ^?p?�?�?N?�?�?�? �?�?�? O6O$OZOHO ~OlO�O�O�O�O�O�O �O __D_2_T_V_h_ �_�_�_�_�_�_
o�_ o@o�Xojo|o&o�o �o�o�o�o�o* N`r�B��� ����&��6�\� J���n�����ȏ��؏ ڏ�"��F�4�j�X� ��|���ğ���֟� ��0��@�B�T���x� ����ү䯎o���̯ ʯP�>�t�b������� �������Կ&�L� :�p�^ϔϦϸ��τ� ����� �"�H�6�l� Zߐ�~ߴߢ������� ���2� �V�D�z�h� ������������� 
�,�.�@�v����� ��\�������< *`N����x ���8J\ (������ ��/4/"/X/F/|/ j/�/�/�/�/�/�/�/ ??B?0?f?T?v?�? �?�?�?�?�?OO�� 2ODO�� O�OtO�O�O �O�O�O_�O(_:_L_ 
__�_p_�_�_�_�_ �_ o�_$oo4o6oHo ~olo�o�o�o�o�o�o �o D2hV� z�����
�� .��R�@�b���v��� &OXO֏菒����� N�<�r�`�������̟ ޟ🮟��$�&�8� n�������^�ȯ��� گ��� �"�4�j�X� ��|�����ֿĿ�� ��0��T�B�x�fψ� �Ϝ����������� >�P���h�zߌ�6߼� �����������:�(� ^�p���R�����8�� ���  &�*�� *�>�*��$�TBJOP_GR�P 2U����  ?�/��C*�	V�]��Wd������X  �*��� �,� � ���*�� @&�?��	 ߐA�����C��  DD�����>~v�>\? ���aG�:�o���;ߴAT������A�<��M�X����>��\)�?���8Q�|����L��>�0 ^&�;iG.���Ap< � F�A�ff�v��� ^):VM�.�� �S>o*�@��R�Cр	���������ff�:��6/�?�33�B   ��/�������>):�S���� �/�/@��H�%&/��/��=� <#��
*��v�;/��f�!?���4B�3 ?'?2	��2?hZ?D? R?�?�?�?F?�?�?�? �?OAOO�?`OzOdO�rO�O�O*�C�*����A��	V3.0}0{�crxl��*P��%�%c5Z F� JZ�H F6� F�^ F�� F��f F� G�� G5 G�<
 G^] G�� G���G��*�G�S G��; G��ERD�u�\E[� E�� F( F�-� FU` F�}  F�N F�� F�� F�ͺ F� F��V G� G�z Ga 9'ѷ�Q�LHefJQ4�o,b*�0c�1���OH�ED_TCH Xd�+X2S��&�&�d$�'X�o�o*�1F�T�ESTPARS c ��cV�HRpABLE 1Yd� N`*�����g)$j�g�h�h)�T1��g	�h
�h�hTHu*��h�h�h�%vRDI0n��GYk}��u	�O �#�-�?�Q�c�u�)r	S�l� �z6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ��I���m�Fwͩ�� ȏڏ쏘������x)r��NUM  ���n����2� Ep�)r_CF�G Z��I���@�V�IMEBF_T�TqD��e޶VE�R�����޳R {1[8{ 8�o�*�%�Q� ��د  9�K�]�oρϓϥ� �����������#�5� G�Y�k�}��ߡ߳��� ��������1���E� W�i�{�������� ������/�A�S�e� w���������������@+=O�_����@��`LIF7 \��D`�����DR�(FP
��!p�!p� d�� ��MI_CHA�N� � DB/GLVL��f�ETHERAD S?u��0`1��_}�ROUT6�!�j!��~SNMASKY|�j255.%�S///A/S�`OOLOFS_DIp��CORQCTRL ]8{��1o�-T�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OL�/6O%O�ZOcPE_DET�AI7�*PGL_�CONFIG �c������/c�ell/$CID?$/grp1^O�O �O�O
__|���G_ Y_k_}_�_�_0_�_�_ �_�_oo�_CoUogo yo�o�o,o>o�o�o�o 	-�oQcu� ��:����� )���_�q���������׮}N����%�@7�I�a�KOq�P��M� ����ʟܟ� �G�$� 6�H�Z�l�~������ Ưد������2�D� V�h�z������¿Կ ���
ϙ�.�@�R�d� vψϚ�)Ͼ������� �ߧ�<�N�`�r߄� ��%ߺ��������� &��J�\�n���� 3����������"��� F�X�j�|��������@��User �View �I}}�1234567890����+=�Ex �e����2 ��B������`r��3�Oas@����x4> //'/9/K/]/�~/x5��/�/�/�/�/?p/2?x6�/k?}?��?�?�?�?$?�?x7 Z?O1OCOUOgOyO�?�Ox8O�O�O�O	_�_-_�ON_TR �lCamera���O�_�_�_�_�_�_˂E�_o)o;n���Uogoyo�o�o�o�)  mV�	�_�o#5 GY o}���o�@�����F_�mV =�k�}�������ŏ l����X�1�C�U� g�y���2�D��"�ן �����1�؏U�g� y�ğ������ӯ��� ��D��k��E�W�i�{� ����F�ÿտ�2�� �/�A�S�e��nUY9 ������������	߰� -�?�Qߜ�u߇ߙ߫� ����v�D�If��-� ?�Q�c�u�ߙ��� �������)�;��� D��I����������� ����)t�M_@q���N�`�93 ��0B��S x�1�����(//�J	oU0�U/ g/y/�/�/�/V�/�/ �/�?-???Q?c?u? /./tPv[?�?�?�? OO(O�/LO^OpO�? �O�O�O�O�O�O�?oU �k�O:_L_^_p_�_�_ ;O�_�_�_'_ oo$o 6oHoZo_;%N��_�o �o�o�o�o �_$6 H�ol~���� moe��]�$�6�H� Z�l��������؏ ���� �2��e&� ɏ~�������Ɵ؟� ��� �k�D�V�h�z� ����E�e��5���� � �2�D��h�z��� ׯ��¿Կ���
ϱ�  ��9�K�]� oρϓϥϷ���������   ��5� G�Y�k�}ߏߡ߳��� ��������1�C�U� g�y���������� ��	��-�?�Q�c�u� ���������������);M_q� � 
��(  �>-�( 	 �� �����#3 5G}k����
� �Y�
// ./��R/d/v/�/�/�/ ����/�/�/A/?0? B?T?f?x?�/�?�?�? ?�?�?OO,O>O�? bOtO�O�?�O�O�O�O �O_KO]O:_L_^_�O �_�_�_�_�_�_#_ o o$ok_HoZolo~o�o �o�_�o�o�o1o  2DVh�o�o�� �	��
��.�@� �d�v��������Џ ���M�*�<�N��� r���������̟�%� ��&�m�J�\�n��� �����ȯگ�3�� "�4�F�X�j������� ����ֿ�����0� w���f�xϊ�ѿ���� �������O�,�>�P� ��t߆ߘߪ߼���� ����]�:�L�^�p�p����߻@ ����������� ���"frh:\t�pgl\robo�ts\crx!�1�0ia_l.xml��D�V�h�z�����`�������������� 0BTfx�� �������, >Pbt���� ����/(/:/L/ ^/p/�/�/�/�/�/�/ ��/?$?6?H?Z?l? ~?�?�?�?�?�?�/�? O O2ODOVOhOzO�O �O�O�O�O�?�O
__ ._@_R_d_v_�_�_�_ �_�_�O�_oo*o<o No`oro�o�o�o�o�ot�n �6� ���<< 	� ?��k!�o;i Oq������ ���%�S�9�k����o�����я����(��$TPGL_O�UTPUT f������� �&�8�J�\�n��� ������ȟڟ���� "�4�F�X�j�|�����в�į�p�ր23�45678901 �����1�C�K��� �r���������̿d��п��&�8�J��} T�|ώϠϲ���\�n� ����0�B�T���b� �ߜ߮�����j���� �,�>�P����߆�� �������x����(� :�L�^���l������� ����t���$6H Zlz���� ��� 2DVh  ������ �/./@/R/d/v// �/�/�/�/�/�/�/ۂ? $$��ί <7*?\?N?�?r?�?�? �?�?�?�?OO4O&O XOJO|OnO�O�O�O�O��O�O_�O0_"_T_} �an_�_�_�_�_�_�]�@�_o	z ( 	 V_Do2oho Vo�ozo�o�o�o�o�o 
�o.R@vd �������� �(�*�<�r�`���ܦ��  << I_ˏݏ������� :�L�֪��}���)��� ş�������k��C� ݟ/�y���e������ �������-�?��c� u�ӯ]�����W��� Ϳ��)χ���_�q�� yϧρϓ�����M�� %߿��[�5�Gߑߣ� ߫���s����!��� E�W��?���9��� ������i���A�S� ��w���c�u����/� ����=)s �����U�� �'9�!o	[ �����K�#/ 5/�Y/k/E/w/�/� /�/�/�/�/?�/? U?g?�/�?�?7?�?�?�?�?	OO��)WGL1.XML�_�PM�$TPOFF_LIM ���P����^FN_�SVf@  �T�xJP_MON Mg��zD�P�P�2ZISTRTCHOK h��xFk_�aBVTCOMPA�T�HQ|FVWVA/R i�M:X�D� �O R_�P��BbA_DEFP�ROG %�I�%TELEOP�i_�O_DISPL�AYm@�N�RINST_MSK  �\� �ZINUSsER_�TLCKl��[QUICKMEyN:o�TSCREY`���Rtpsc�Tat`yixB�`�_�iSTZxIRA�CE_CFG Uj�I:T�@	[T�
?��hHNL C2k�Z���aA[ gR -?Qcu�����z�eITEM 2�l{ �%$1�23456789y0 ��  =<
�x0�B�J�  !P�X�dP���[S��� "���X�
�|���W� ��r�֏����.��0� B�\�f�����6�\�n� ҟ��������>�� �"���.�����ίR� ���Ŀֿ:��^�p� 9ϔ�Tϸ�xϊ�� �d���H��l��>� Pߴ�\�������v� � �����h�(�ߞ߰� 4�L��ߦ�����@� R��v�6���Z�l��� �������*���N���  ������������X ���J
n� ��b���� "4F�/|</N/ �Z/���//�/0/ �/?f/?�/�/e?�/ �?�/�?�?�?,?�?P? b?t?�?�?DOjO|O�? �OOO(O�O�O^O_ 0_�O<_�O�O�_�O�_ _�_�_H_�_l_~_Go��dS�bm�oLj�g  �rLj �a�o�Y
 �o�o�o��o{jUD1:\�|��^aR_GR�P 1n�{� 	 @�PRd{�N�r����~� �p���q+��O�:�?�  j�|�f� ���������ҏ��� �>�,�b�P���t���������	e���~\cSCB 2ohk U�R�d�v����������Я�RlUT�ORIAL p�hk�o-�WgV_CONFIG qhm��a�o�o��<�OUT?PUT rhi}�����ܿ� � �$�6�H�Z�l�~ϐ� �ϴ�z�ɿ���� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r �������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/��/�/??0?B? T?f?x?�?�?�?�?�/ �?�?OO,O>OPObO tO�O�O�O�O�?�O�O __(_:_L_^_p_�_ �_�_�_�_f�x�ǿo o,o>oPoboto�o�o �o�o�o�o�O( :L^p���� ���o ��$�6�H� Z�l�~�������Ə؏ ��� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я���� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t�����������������X���#��N �_r������ �&8J��n �������� /"/4/F/X/i|/�/ �/�/�/�/�/�/?? 0?B?T?e/x?�?�?�? �?�?�?�?OO,O>O POa?tO�O�O�O�O�O �O�O__(_:_L_^_ oO�_�_�_�_�_�_�_  oo$o6oHoZok_~o �o�o�o�o�o�o�o  2DVgoz�� �����
��.� @�R�d�u�������� Џ����*�<�N� `�q���������̟ޟ ���&�8�J�\�k���$TX_SCR�EEN 1s%� �}��k�����ӯ���	� ��Z��I�[�m���� ���,�ٿ����!� 3Ϫ�W�ο{ύϟϱ� ����L���p��/�A� S�e�w��� ߭߿��� �����~�+��O�a� s���� ���D��� ��'�9�K������ ����������R���v� #5GYk}�����$UALRM_�MSG ?����� �n��� 	:-^Qc������� /�SEoV  �2&��ECFG uv����  n��@�  Ab!  w B�n�
 / u����/�/�/�/�/�/�??%?7?I?W7>!G�RP 2vH+ 0n�	 /�?� �I_BBL_NO�TE wH*T?��lu����w�T �2DEFP�RO� %� (%�Ow�	OBO-OfO QO�OuO�O�O�O�O�O�_�O,_�<FKEYDATA 1x����0p W'n���?�_�_z_�_�_�Z,�(�_on�(PO�INT Koo ? IRECT@oko��PNDUo�oOcCH�OICE]�onTOUCHUP�o �o�o�o8\n U�y�������"�	�F��Y���/frh/gui�/whiteho?me.pngQ��������ŏ׏�h�pointz���/��A�S��  i�direc��������şןf�/iny��"��4�F�X��m�choicy�������ͯ߯��h�touchup���/�A�S�e���h�arwrg �����ÿտ�n�� �(�:�L�^�p����� �ϸ�������}��$� 6�H�Z�l��ϐߢߴ� �������ߋ� �2�D� V�h�z�	������� ������.�@�R�d� v���_����������� ���2DVhz ������
 �@Rdv�� )����//� </N/`/r/�/�/%/�/ �/�/�/??&?�/J? \?n?�?�?�?3?�?�? �?�?O"O�?4OXOjO |O�O�O�OAO�O�O�O __0_�OT_f_x_�_ �_�_=_�_�_�_oo ,o>o�_boto�o�o�o��oW��k�b�����o}�o8J$v,6�{.�� �������/� �S�:�w���p����� я�ʏ��+��O� a�H���l�������ߟ ���'�9�Ho]�o� ��������ɯX���� �#�5�G�֯k�}��� ����ſT������ 1�C�U��yϋϝϯ� ����b���	��-�?� Q���u߇ߙ߽߫��� ��p���)�;�M�_� �߃��������l� ��%�7�I�[�m��� ������������z� !3EWi���� �����П/ ASew~��� ���/�+/=/O/ a/s/�//�/�/�/�/ �/?�/'?9?K?]?o? �?�?"?�?�?�?�?�? O�?5OGOYOkO}O�O O�O�O�O�O�O__ �OC_U_g_y_�_�_,_ �_�_�_�_	oo�_?o Qocouo�o�o�o:o�o �o�o)�oM_ q���6������%�7�9�}����b�@t���^�������,�� 돞����3�E�,�i� P�������ß����� ����A�S�:�w�^� ������ѯ����ܯ� +�
O�a�s������� �Ϳ߿���'�9� ȿ]�oρϓϥϷ�F� �������#�5���Y� k�}ߏߡ߳���T��� ����1�C���g�y� ������P�����	� �-�?�Q���u����� ������^���) ;M��q���� ��l%7I [������ h�/!/3/E/W/i/ @��/�/�/�/�/�/� ??/?A?S?e?w?? �?�?�?�?�?�?�?O +O=OOOaOsOO�O�O �O�O�O�O_�O'_9_ K_]_o_�__�_�_�_ �_�_�_�_#o5oGoYo ko}o�oo�o�o�o�o �o�o1CUgy ������	� ��?�Q�c�u����� (���Ϗ������ ;�M�_�q�������~ ����~ ���ҟ���Ο�*��,�[���f��� ����ٯ�������3� �W�i�P���t���ÿ ���ο��/�A�(� e�Lωϛ�z/������ ����(�=�O�a�s� �ߗߩ�8�������� �'��K�]�o��� ��4����������#� 5���Y�k�}������� B�������1�� Ugy����P ��	-?�c u����L�� //)/;/M/�q/�/ �/�/�/�/Z/�/?? %?7?I?�/m??�?�? �?�?�?���?O!O3O EOWO^?{O�O�O�O�O �O�OvO__/_A_S_ e_�O�_�_�_�_�_�_ r_oo+o=oOoaoso o�o�o�o�o�o�o�o '9K]o�o� �������#� 5�G�Y�k�}������ ŏ׏������1�C� U�g�y��������ӟ ���	���-�?�Q�c� u��������ϯ��h���0���0���B�T�f�>�����t�,��˿~� �ֿ�%��I�0�m� �fϣϊ��������� ��!�3��W�>�{�b� �߱ߘ��߼�����? /�A�S�e�w��� ������������=� O�a�s�����&����� ������9K] o���4��� �#�GYk} ��0����/ /1/�U/g/y/�/�/ �/>/�/�/�/	??-? �/Q?c?u?�?�?�?�? L?�?�?OO)O;O�? _OqO�O�O�O�OHO�O �O__%_7_I_ �m_ _�_�_�_�_�O�_�_ o!o3oEoWo�_{o�o �o�o�o�odo�o /AS�ow��� ���r��+�=� O�a����������͏ ߏn���'�9�K�]� o���������ɟ۟� |��#�5�G�Y�k��� ������ůׯ����� �1�C�U�g�y���� ����ӿ������-�@?�Q�c�uχ�^P����^P���������ͮ���
���, ��;���_�F߃ߕ�|� �ߠ����������7� I�0�m�T������ �������!��E�,� i�{�Z_���������� ���/ASew ������ �+=Oas� �����//� 9/K/]/o/�/�/"/�/ �/�/�/�/?�/5?G? Y?k?}?�?�?0?�?�? �?�?OO�?COUOgO yO�O�O,O�O�O�O�O 	__-_�OQ_c_u_�_ �_�_:_�_�_�_oo )o�_Mo_oqo�o�o�o �o���o�o%7 >o[m���� V���!�3�E�� i�{�������ÏR�� ����/�A�S��w� ��������џ`���� �+�=�O�ޟs����� ����ͯ߯n���'� 9�K�]�쯁������� ɿۿj����#�5�G� Y�k����ϡϳ����� ��x���1�C�U�g� �ϋߝ߯�����������`����`���"�4�F��h�z�T�,f���^���� �����)��M�_�F� ��j����������� ��7[B� x�����o! 3EWixߍ�� �����///A/ S/e/w//�/�/�/�/ �/�/�/?+?=?O?a? s?�??�?�?�?�?�? O�?'O9OKO]OoO�O O�O�O�O�O�O�O_ �O5_G_Y_k_}_�__ �_�_�_�_�_o�_1o CoUogoyo�o�o,o�o �o�o�o	�o?Q cu��(��� ���)� M�_�q� �������ˏݏ�� �%�7�Ə[�m���� ����D�ٟ����!� 3�W�i�{������� ïR������/�A� Яe�w���������N� �����+�=�O�޿ sυϗϩϻ���\��� ��'�9�K���o߁� �ߥ߷�����j���� #�5�G�Y���}��� ������f�����1��C�U�g�>�i��>>�������� ����������,� �?&cu\�� �����) M4q�j��� ��/�%//I/[/ :�/�/�/�/�/�/�� �/?!?3?E?W?i?�/ �?�?�?�?�?�?v?O O/OAOSOeO�?�O�O �O�O�O�O�O�O_+_ =_O_a_s__�_�_�_ �_�_�_�_o'o9oKo ]ooo�oo�o�o�o�o �o�o�o#5GYk }������ ��1�C�U�g�y��� �����ӏ���	��� -�?�Q�c�u�����p/ ��ϟ�����;� M�_�q�������6�˯ ݯ���%���I�[� m������2�ǿٿ� ���!�3�¿W�i�{� �ϟϱ�@�������� �/߾�S�e�w߉ߛ� �߿�N�������+� =���a�s����� J�������'�9�K� ��o�����������X� ����#5G��k�}���������������&�HZ4,F/�>/���� �	/�-/?/&/c/J/ �/�/�/�/�/�/�/�/ ?�/;?"?_?q?X?�? |?�?�?���?OO%O 7OIOXmOO�O�O�O �O�OhO�O_!_3_E_ W_�O{_�_�_�_�_�_ d_�_oo/oAoSoeo �_�o�o�o�o�o�oro +=Oa�o� �������� '�9�K�]�o������ ��ɏۏ�|��#�5� G�Y�k�}������ş ן������1�C�U� g�y��������ӯ� ��	��?-�?�Q�c�u� ��������Ͽ��� Ϧ�;�M�_�qσϕ� $Ϲ��������ߢ� 7�I�[�m�ߑߣ�2� ���������!��E� W�i�{���.����� ������/���S�e� w�������<������� +��Oas� ���J�� '9�]o��� �F���/#/5/�G/�$UI_IN�USER  ����h!��  H/L/_�MENHIST �1yh% � ( u ���)/SOFTP�ART/GENL�INK?curr�ent=menu�page,1133,1�/�/??�'�/�.71�/{?�?ȟ?�?�+E?�%ed�it�"TELEOPj?OO'O�?D?V?�2�/�O�O�O�O�(<MO�/48,2�O
__._@_��A_f_x_ �_�_�_�_O_�_�_o o,o>o�_boto�o�o�o�o�m�\a�!\o�o /ASVow� ����`��� +�=�O��������� ��͏ߏn���'�9� K�]�쏁�������ɟ ۟j�|��#�5�G�Y� k���������ůׯ� �o�o�1�C�U�g�y� |�������ӿ����� �-�?�Q�c�uχ�� �Ͻ�������ߔ�)� ;�M�_�q߃�ߧ߹� ���������7�I� [�m��� ������ ��������E�W�i� {��������������� ��ASew� ��<��� +�Oas��� 8���//'/9/ �]/o/�/�/�/�/F/ �/�/�/?#?5? �2� k?}?�?�?�?�?�/�? �?OO1OCO�?�?yO �O�O�O�O�ObO�O	_ _-_?_Q_�Ou_�_�_ �_�_�_^_p_oo)o ;oMo_o�_�o�o�o�o �o�olo%7I�[F?��$UI_�PANEDATA 1{����q�  	��}  frh/�cgtp/fle�xdev.stm�?_width=�0&_heigh�t=10�p�pic�e=TP&_li�nes=15&_�columns=�4�pfont=2�4&_page=whole�pmI6?)  rim�9�  �pP�b�t����� �������Ǐ��(� :�!�^�E�����{������ܟ�՟�I6�� �   ?  "�J�O� a�s���������ͯ@� ���'�9�K���o� ��h�����ɿۿ¿�� �#�5��Y�@�}Ϗ�vϳ�&��Ɠs��� ��)�;�Mߠ�q�� �ߧ߹�������V�� %��I�0�m��f�� �����������!�� E�W����ύ������� ����:�~�/AS ew����� � =$as Z�~����d� v�'/9/K/]/o/�/� �/�/*�/�/�/?#? 5?�/Y?@?}?�?v?�? �?�?�?�?O�?1OCO *OgONO�O�/�/�O �O�O	__-_�OQ_�/ u_�_�_�_�_�_6_�_ o�_)ooMo_oFo�o jo�o�o�o�o�o�o %7�O�Om�� ���^_�!�3� E�W�i�{������Ï ���������A�S� :�w�^�������џD V��+�=�O�a��� ����
���ͯ߯�� �|�9� �]�o�V��� z���ɿ���Կ�#��
�G�.�k�ޟ�}��|ϵ����������) ��4ߧ�#�`�r߄ߖ� �ߺ�!���������� 8��\�C���y�� �����������������$UI_POSTYPE  ���� 	 ��s�B�QUICKMEN  Q��`�v�D�REST�ORE 1|���  �	�����������mASew�, ������+ =Oan�� ���//�9/K/ ]/o/�/�/6/�/�/�/ �/�/�??0?�/k? }?�?�?�?V?�?�?�? OO�?COUOgOyO�O 6?@O�O�O.O�O	__ -_?_Q_�Ou_�_�_�_ �_`_�_�_oo)o�O 6oHoZo�_�o�o�o�o �o�o%7I[��o������S�CRE��?���u1sc���u2�3�4�5*�6�7�8��swTATM�� ��<��:�USER�p�2�rT�p�ks���U4��5��6��7���8��B�NDO_CFG }Q������B�PDE���?None��v��_INFO 2~j��)���0%� D���2�s�V������� ͟ߟ��'�9���]�o�R���z��OFFSET �Q�-���hs��p��� ��G�>�P�}�t��� Я��׿ο���� C�:�L�^Ϩ����͘ς��
����av��W�ORK �!������.�@ߢ�u�UFRAME  ����RTOL_A�BRT�����EN�B�ߣ�GRP 1������Cz  A������*�<�N�`�r��֐�U������MSK  ��)���N��%�!��%z����_EVN�����+�ׂ�3�«
 h��UEV��!t�d:\event?_user\�u�#C7z���jpF��n��SPs�x�spo�tweld��!�C6��������! ���G|'��5k Y�����> ���1�Ug ���/��	/^/ M/�/-/?/�/c/�/�/ �/�/$?�/H?�/:J��W�3�����8C?�?�? �?�?�?�? O+OOOOaO<O�O�O rO�O�O�O�O_�O'_ 9__]_o_J_�_�_�_��$VALD_C�PC 2�« ��_�_�  w��qd�R�*o_oqo��
hsNbd�j�`��i �da{�oav�_�ooo 3BoWi{�o�o�o �o��o�PA� 0�e�w������ ����(�=�L�a� s�
�������ʏ��� ��$�ޟH�:�o��� ������ڟ؟�����  �2�G�V�k�}����� ��¯ԯ�����.� �R�S�yϋϚ����� �����	��*�<�Q� `�u߇ߖϨϺ����� ����&�8�M�\�q� ���߶���n����� �"�4�F�[�j���� ������������! 0�B�Wf�{���� �������,> teT����� ��/+/:La/ p�/�/./���� �//'?6/H/?l/^? �?�?�/�/�/�/�/? #O�?D?V?kOz?�O�O �?�?�?�?�?_O1_ @ORO9_vOw_�_�_�O �O�O_�__-o<_N_ `_uo�_�o�o�_�_�_ �_o&o;Jo\oq �o����o�o�o�  �"7�FXj�� ���������!� 0�E�T�f�{������� ßҏ����
�,�A� P�b�����x�����Ο �����(�*�O�^� p���������R�ܯ�  ��Ϳ6�K�Z�l�&� ���Ϸ���ؿ���"�  �2�G���h�zϏߞ� ����������
��1� @�U�d�v�]�ߛ��� �������,��<�Q� `�r���������� ����&�;J�_n� ������������ �$F[j|� ������ 0E/Ti/x��/� �/�/�/�//,/.? P/e?t/�/�/�?�?�? �?�/??(?:?L?NO sO�?�?�O�?�O�OvO  OO$O6O�OZOo_~O �OJ_�O�_�_�_�O_� _F_D_V[�$VA�RS_CONFI�G ��Pxa�  FP�]S�\lCMR_�GRP 2�xk� ha	`�` � %1: SC�130EF2 *H�o�`]T�VU�P�h�`�5_Pa?��  A@%pp*`�NVn No9xC VXdv��a��<u�A�%p�q�_R���_R B���#�_Q'��H�� l�;���{�����؏Ï Տ�e��D�/�A�z��-�����ddIA_W�ORK �xe�ܐ�Pf,		�Qxe���G�P ����YǑRTSY�NCSET  �xi�xa-�WINU�RL ?=�`�����������ȯگ�SIONTMO�U9�]Sd� ���_CFG ��S۳�S۵P��` FR:�\��\DATA\�� �� M�C3�LOG@�  � UD13�EX�d�_Q' B@ ����x�e_ſ�x�ɿ�VW �� n6  ����VV��l�q  =���?�]T<��y�Y�TRAIN؎��N� 
gp?�CȞ��TK���b�xk (g����� _���������U�C� y�g߁ߋߝ߯����߮�_GE��xk�`_P�
�P�R���RE��xe*�`h�LEX�xl`1�-e�VMPHA�SE  xec��ecRTD_FILTER 2�xk �u�0��� �0�B�T�f�x����� VW�������� $�6HZl_iSHI�FTMENU 1��xk
 <�\%�������� ��=&sJ\ �������'/��	LIVE/�SNA�c%vs�fliv��9/���� 7�U�`\"menur/w//�/�/������]��MO���y��5`h`ZD�4�V�_Q<��0���$WAITDIN�END��a2p6OK  �i�<���?�S�?�9TIM�����<Gw?M�?*K��?
J�?
J�?�8RELE��:G6p3���r1_ACTO 9Hܑ��8_<� �ԙ��%�/:_af�BRDI�S�`�N�$XV�R��y��$Z�ABC�b1�S;S ,��j�I�2B_�ZmI1�@VSPT ��y��eG�
�*�/o�*!o7o�W�DCSCHG �ԛ(��P\g@��PIPL2�S?�i��o�o�o�ZMPC?F_G 1��ii��0'¯S;Ms�S���i��p'��g�8�G�8��q��O<��� Z�A���g���4����ٿ�P��	�`�p	9�WS��AC�ײ�&��úםI��?g��i��?��4�����>��� ���>س�ߢ�ui7�p
��p��s��p9��S^�t����*�t��p4�p���� �v�|~��g�Ï��y��3�@���C�|��ۃA���_��|#�҉������*�@�N�x��w������%�r����F��=�^S�*F�׽��j���D?V��C_!��U�I�0�����2[?��A���A�>�P�.+Ǿ��@��Zp���o�_C_YLIND�� {� Х� ,(  *=�N�G�:�w�^����� ��ѯ� ��7����<�#�5�r� ����������޿y�_� ���8�ύ�nπ��r�ã wQ �5 �����S�����(��h��X�זr�A���SPHERE 2���ҿ��"ϧ��� ���P�c�>�P�̿t� ��ߪ�����'�� �]�o�L���p�W�i�������������PZZ�F �6