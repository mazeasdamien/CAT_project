��   �A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����CCSCB3�_GRP_T �  � $FS�_TYP3  �$PS_SBF�RAME3��$�J  $INIT_TOL^�RANGE3_F�_uT~FTR/ATIO^c ��P_H_LIMA��L�FSOF�ST_S^JM3�_f _���$$�CLASS  O������[���[� VERSIO�N�  �XKIRTU�AL��' 3 �[� 6  ������b@��  B ��B A�����Cp  T�aY��B�z��m