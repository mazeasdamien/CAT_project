��   C��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN��/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER��q�C_GRP6�P L$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� )DEX� �5O n�8BUF�7TDP�HG�_@FO�SxAV��7R?EC_TRQX��MFLG�J5�� � � N IU�
@!(UF*����4OSV3EN_CG"��0_�!�AU�SCH2�SMP]L4PEXE���2�!_�SUR}A�`jAaW�@A@bVNE|Y]QnAVA?�UY�T7D�VWWnAF�[V�A�\�WTO�0oH
e7D�f�3
e�U
e�W QT�P�0IR	 DMM��A@  @ �$la�EREG_�OFS�aME�hA1SS1�A !la�RE-   �# �0�b{F�c{ĥd� M�d�b�c$�STD�hq�gFA � �h!q�g�"�f�"�c�/ la7   �$p`TIN�@��0SUL� �R}_@  $}�@ SW@�rO:}rR%	 dp~t�� �@JU� �s �/ FS4D6
 O� $�0PGF`~QC!$FIL�  �@�E�PmA�s�&�DIG4o@SCA��$�INTT?HRS_BI�AZ��SMAL%�CO�L��qATE_T=I�PROG�4U��s�!CMDAp FSOUTENV6�P $HR�Z_AXl�CU3VR2QLB܊�0���H������PNT_MV_AVR�C�S!pLkp�c$L`���fO�\��ST�:d�F�#STO v��FX�LECTEdDCp�Y{���FY��2t�Z{�ړFZc�!R�e��	�/ G#P�X $��c_IV����$!�0B"0�?0F�CC�BDDN=�CCI�c�DUMMY23<G ^�DEBU�A\!4PN�"TO�q9RP" � Q09T6�� �;!��NfBUTTSP� (~@�q֥E40N ڡFS3ՁKQ1�r�9T�I�NEW_�UI��VKP�?Up`��CCOORD8\TCH���01�P���mP��)��l �!�3?$WEIGH���2� s_�aF��Tƿ�WA{Q����NTER�Q��- ޵� �c䮱�AS0�$JnZASTA�� �a���� �,�26�36�W�!Ƨ ��ä"UC��Xw�Yw�Zw�6_�CM��?��D��i�RSLy�u���@~��Ǝ��ƚ�	"_Ϡ�_ҡ)�  E�0c"0VROUN�DCMVPERIO���$F1PUU3F2D�'TM1� ��S�_DcGAMqMc1b�TRX�U�Kt�K�K��CLt�`�&O00ADJ�GA�UPDC0R"�2��E� QRED���GFR_� _@W۲���u�DL_R���@�=�M_�5d�0 n�#��}�"��}�� k�����������}�VLj�"����A� 7���`��L�P5A8@
� 
D�A�����"�8��y"��VIBƦ�OV��DEH�֌� �`,����*�� �: RTZ�MN1SUfwMN2YUFRA q	��ShZA
`-G����OR�P�ҡAL�ҤCJ��
L��"�S8B�I$L .$M"�P30+�Q �)k�}�S"PHCmD�GVz�GV��;GVړJDO°]���S�$R�E����b�]�A�AP�)�DA��3$VF�����1LVu��@IL�A���� #��  "�@fR!��$�DC+�����B #П�5'OBOA@�vYԣW2
�G'	�$�ԍ$!#¿�E�K�`�+�eCNPRGOV6��%'PN�t_TW,��"G�3E�MNV�6c0�4WT�cW�TRL/_SKIj�J�qcMN��GW6�
eR<ENABF��rV!�� A$SB}��xS���{P �tyR*�tX�yRQT$���2_Q��?p����ALARMSE�R�QETOTDFRZCHK1����62�9NC�4N@�5�L`N@�:vJ��vE�22��;2�=NA9E�FFI�X2��BF�䦠@I8�dD���DON�t�9�5PSFW�0_DF1"%BF2/_vJ��H|��4|�Pl��33=��5|�kH|�yJ�Z���U�23�;3�=|�9E�SDIAu �6�RKqB�B�VvEfvC�3GA�@�@���R<i V1<d��sP�VQ�U�Uf�S$��� ��F�U�ED�S_H�A�U�e�d�4GEF�k@�2�`�;�a�@�5!%�UzKq�#�$X�(��s���Y���a=�@rSIW(�� � *�X�R�K��`H7p_CHsCK�!'�INS��@�w <B
U; �zH�NT���v�y�A`&|  ��w�ΰP���쑎�����$���� ����2�=�=� 9'���SIOe�1�wkpXKC��IRTU&@0�B�C|�,SV 2n��� X  Ф������͊@͉	������F�@ �߀��B�O  =�kp5� a�s���������ŕ=�d=�
ݐh����� ���6�X�$�n�W�8� P�b�|���ՒN����� ̯⯨����*�8�f� �n�X�����ҿ���� Ŀ���ڿ��X�j� ��FϘϊ�����߲� ���L�B�p�ߔ�b� �߮�x���6���H���7�I�:�	UD�1: 678  �Afsdt1 �78901234�5r�����  )�y�q�����.0����X�\�'Q���
� l#�5�B�~P1�+�|�o������� ��������0'9 Rx_�����~�DMM P����A U�W�(F�Xj��POR 2]	 [����Z1F���B?��S4D 
!x�	/'���,/>/��v}?��B�l ���)***@/�/#!{/�/��C�pONFIG� n����9�2[� e�$��/ّ�7  �z  D30h25Y��>�P0����C  C�3�h1�2D�D�/B42�3N �#� 3�,�Ӳ?o�?��:�ד�=���As!�=�O<O 3O��rO]OoO�O�O�O�O�O�O_� � :Z#S8_J_\_n_�_ �_�_�_�_�_�Y_!o oEo0oioTo�oxo�ot�o�I�� 3 [��`�g4 A�e�g ���01Bk!t�1C�`0.t���=#�
��Nn{k(EuK��Qu�LE@��eeu=D���qu��;��ʞ�u8I��u��It$ �$�m5@r�I���uFۀ3�uBQOGO�����t��+���E�.����Q���$�=�a�(4$�m�%��7�>�E���B<�~w����8E�y���;�j��ar�{�х>��݅���?s ���BHx�g!s >��� A!@��?E��qJ�b��@�sF��3{Fs�"��E~��b��vC��C��B��B ������j!AAo!k!�Bpp#B6q��f!Ju�@u�@�s @p0@�u�:p73� 	�	��l�c�u�����.pݑ Bo C��?�d��g ݯ��`?��33���a:�o-�?��a��c��������������ڿ�?�Ls�S�c��8< ��Na'����B��� ��̻p0%rk�a��8
/x���
�� <�>�-2��nπ�ߤ� ���������߾�P��J������� �����V�A����@� ��)qݑ��)r����·������	��c)�F������� O�a���ڑ��)rk �v�l�1��_FC�COORD 32 `!�?��� ����r���
 �=�d&�J |���/��*/ �]//2/�/F/�/j/ �/�/�/�/#?�/�/J? ?}?0?R?�?f?�?�? �?�?�?�?CO�?OjO ,O�OPOrO�O�O�O�O �O__�Oc__8_�_ L_�_p_�_�_�_o�_ �_>o$oo�o6oXo�o lo�o�o�o�o7�o ^D2�Vx� ����$��W�
� <�~�d�R�Ïv���� ���Џ�D��w�*� \�����r�㟖���
� ̟=���d�&���J� |����������د*� �]��2���F���j� ��޿Ŀ��#�ֿ��J� �}�0�RϤ�f��ϊ� ��������C����j� ,ߝ�P�r��߆��ߪ� ������c��8�� L��p�������� ��>�$����6�X��� l���������7�� ^D2�Vx� ����$�W
 <~dR�v�� �/��D//w/*/ \/�/�/r/�/�/�/
?� 3�$CC_FS�IW ����>1� �  6M81 Y<w?�?�4