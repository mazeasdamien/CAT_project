��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1�TU4QQ  �AR�x1R� � /$TIT91� �� � �Td�T0�ThP�TU5�V6�V7�V8�V9�W0�W�WOQ�U�W�gQ�U�W1�W1�W1��W1�W2�R�SBoN_CF�!@$<!J� ; ;2�1�_CMNT�$�FLAGS]�C�HEK"$�b_O�PTJB � ELL�SETUP � `@HO8@9 P�R�1%�c#�aREPR�hu0D+�@���b{uHM9 MN�B;16 UTOB�J U�0 }49DEVIC�STI/@�� �@b3�4pB�d�"VAL��#ISP_UNI�tp_DOcv7�yFR_F�@|%u13���A0s�C_WAx�t,q�zOFF_T@]N�DEL�Lw0pdq�1�Vr?^q��#S?�o`Q"U��t#*�QTB��bMyO� �E � �[M�����RE�V�BIL���!X�I� v�R  �!D�`��$NOc`M�|����ɂ/#ǆ� �ԅ��ނ�@Ded �p E RD_E���h�$FSSB�6�`KBD_SEV�uAG� G�2Q"!_��2b�� V!�k5�p`(��C�00q_ED|� � � t2d�$!S�p-D%$� ��#�B�ʀ_�OK1��0] P_C�� ʑ0t��U �`LACI�!�a�Y�� ��qCOMM� # $D
� ��@���J_�\R BIGALL;OW� (Ku2:-B�@VAR���!�AB mPBL�@� �� ,K�q���`S�p�@M_O]˥���CCFS_U	T��0 "�A�Cp'���+pXG��b�0 =4� IMCM ��#�S�p�9���i �_D�"t�b��M�1� h$�IMPEE_F�s��s��0� t����D_���J��D��F��%�q_����0 T@L��L�DI�s@G�^� �P��$I�'�����CFed X@G�RU@��Mb�NF�LI�\Ì@UIR�E�i42� SWIYTn$`0_N�`S 2�CF�0M� 	�#u�D��!��v`(����`J�tV��[ �E��.p�`�ʗELBOF� �շ �p`0���3����� F�2T��A`�rq1�J1��z _To!@��p��g���G�� �r0WARNM�p#tC�v`�ç` �� COR-UrF�LTR��TRAT�9 T%p� $AC�CVq��� ��r$�ORI�_&�RT���S<���HG�0I����TW��A�I�'�T��1D���� �202�a1��HSDR�2��2�2J; �S���3��4��5���6��7��8��9Ə� �׀
 �2� @� TRQ�$�vf��'�1�<�_U�<�G��Oec  <� P�b�t�53>B_�LLEC��!~�MULTI�4�"u�Q|;2�CHILD���;1?�O�@T� "'�STY92	r��=��)2���ױ��ec# |r056$J ђ��`���u�TO���E^	EX�Tt����2��2�2"y����$`@ D	�`&�ᣡ����� (p�"��`%�ak�����s�����&'�E�A�u��Mw�9 �% ���TR�� ' L@U#9 ���=At�$JOB���мP�TRIG��( dp������^'�#j�~�l�CpO�R�) t$�F�L�
RNG%Q@�TBAΰ �v&r�*`1�t(��0 �x!�0�+P`�p�%��`��*�Ё͐U��q�!�;2J��_R��>�C<J��8&<J D`5C�F9���x"�@J��Pq_p�7p+ \@�RO"pF�0��IT�s�0NOM��>Ҹ4Ps�2�� @U<PPg�*��P8,|Pn��0b�P�9�͗ RA����l�?C�� �
$T\ͰtMD3�0T���pU�`�΀+AH,lr>�T1�JE�1\� J���PQ��\Q��hQC�YNT�P��PDB�GD̰�0-���P�U6$$Po�|�u�AqX����TAI�s�BUF,�y��A�1.c ����F�`PI|��-@PvWMuXM�Y�@�VFvWSIM�QSTO�q$KEE�SPA��  ?BP�B>C�B�P��/�`=��MARG�u2��FACq�>�SLEW*1!0����
�6�RMCW$0'����pJB�Ї�qDE�Cj�exs�V%w1 Ħ�CHNR�;MPs�$G_@�g�D�_�@s��1_FP�5�@TC�fFӓC@�Й���qC��+�VK��*��"*�JRx���SoEGFR$`IOh!v�0STN�LIN>�&csPVZ�WQ_�A�D2����r 2��hr�r�?�P��3` +^?���եq�`��q�|`�����t��|aSCIZ#�!� �T�0_@%�I��qRS� *s��2y{�Ip{�pTp�LF�@�`��CRC����CCTѲ�Ipڈp�a���bL�MIN���a1순���D<iC �C/���!uc�OP4�Ln j�EVj���F��_!uF��N����|a(��=h?KNLA�C{2�AVSCAB�@A��R�@�4�  cSF�$�;��Ir �4�@�05��	D-Oo%g��,�,m����ޟ��BR>C�6� n����sυ�U��R�0HA;NC��$LG��ɑ6DQ$t�NDɖ��AR۰N��aqg�����X�ME��^�Y�[PfS�RAg�X�AZ��蟸��rEOB�FCT ��A��`�2t!Sh`0ADI��O��y�s" y�n!�������~#C�qG3t!��BMPmt�@�Y�3�afAES�$�����W_;�BA�S#XYZWPR$��*�m!��	y�U�87  ƀI�@d���8\�p_C�:T���#��R_L\
 � 9 ���C��/�(zJ�LB�$��3�D��5�FOsRC�b�_AV;�'MOM*�q�SaԫBP`Ր�y�HBP�ɀE��F����AYLOAD&$ER�t&3��2�Xrp�!�zR�_FD�� : ET`I�Y3��E�&���Ct��MS�P�U
$(kpD���9 �b�;�B�	EV�Id�
�!_IDX��$���B@`X�X<&�SY5�  �HOPe�<>��ALARM��2W̭rY�R_�0= !hb Pnq�`M\qJ@O$PL`A&�M#�$�`��� 8�	���pV�]�0����CU�P�M{�U��>�TI-Tu�
%�![q���Z_;���? ��B pQk��6NO_HEADE^az��} ѯ��`􂳃���dF� ق�tP ���@�@|��uCIRTR�`$��ڈL��D�CB@4�RJ��
�[Q���cA�2>���OR�r���O����T`UN_OO�Ҁ$����T(�����I�VaCx�=� PXWOY���=B��$SKADR���DBT�TRL
��C��րfpbDs�L�~�DJj4 _�bDQ}��PL�q�wbWA���WcD��A��A=�2�U�MMY9��10L���DB����D;�[QPR�� 
9��D�Z���E lO�Y1$�a$8�/��L)F!/�������0GG/_cP�C�1Hf/x$ENE
A@Tf�I�/��,$��COR`"JH y@ �E$L�#F$#PR���+jp���nq�_D$�qPROSS]�
���R�r�` >u�$TRIG96�PAUS73ltETgURN72�MR:�eU 0Ł0EW$�~�`SIGNALA��QR$LA�З5�1�G$PD�H$PDİ�AI�0�A�C�4�C��DO�D�2�!��6GO_AWA�Y2MOZq�Z��� CS��CSCB�g�K Իa#���E+RI�0Nn�T�`$�����FCBPL�@QBGAGE���P��ED`|BD�wA[CD�OF�q�[F0�FoC��MPM�AB0XoC�$FRCIN��2Dk��@��O$NE�@�FD�L8�� L� �����=��Rw�_��P>� OVR10����lҠ�$ESC_|�`uDSBIO��p��pTe�E�VIB�� `s��Z��V��p�SSW��$�VL��:�Lk��X���ѣ�0bQ����USC�P��qA=�	Q��MP1%e@&S*`�(bt`'c5۳ESUd��-cWg&S Wg?cWd����Wd��Wd<.���AUTO$�Ya҃�ac�SB����-d���&SwB[��GB�f_$VOLT�g ���  �GAOD!��q���@:�ORQ�ҀKra�$DH_THE&0�Rgp� <qtnwALPHnt��o��w0 Vp]�$�.�Ra�[��s�5�`r�CQ�#BUD�S� F1M���sV
��;��L�b�tk���BRTHR��L��T`�Z���Vɖ��D)E  �1��2�⋅ ��������kѯ�a� �Tt0V�ꆸ������@̈Я�-�"�N~���sS2����INHB��ILTG0ɡ�T?� �3$�w��E��PqQxQ��TqPe��0Y�AF}�O�ນ��ڗ ��qPڳē����bPܙ���PL?���3���TMOU��ēS��� � ��s�/�S18���O��Aܙ��I����CDqIƑ˩o�STI��գ�O:ҋ�,0���AN��Qg�S��+r�#x$�����w�1_����PRA�P`�vC����MCN�eQe�����VER�S��r�oPIw�F�PåǲШ۷G.�DEN��G>�����F�2H�Ƿ�M�7�F��_�MN�D̠,���@�d�{ƭa����OB����U˱z���DI ���#���3�����A��w�Fx���3�O�N�5��Q��VAL��CR[�_SIZp��b�;Qn�REQ�R�b��]2b���CH q�΂�ڃ�Ռ�����:�n�S_U��X��wW�FLG���wU$CV�iMGP�QδFLXP�923R�u�L��EAL�P-�C	��+rT��W��� �R��c���NDMS�7� ��K>S�P_M'0h�STWv������AL�P���Q����U���U�IAG@,�o��d�U�-�T"	A-`� ���A��� ��H`��Q`��6��Pq_D&��1s��.�P��F�>2�T�� ?7 1A>���#�#L��?`_=i @@>LD�pc���0�FRI�0 `Ѐ��1}Ѳ�IV\1�*�^1�U�P`��a��C�L!W��
`L=S&-c&&S�C.w��  L���!����d�Q$w!�҇��$w��p��
�P�5RSM��P���V0h � r�l�d^2AW�a_TRp�}�8@NS_PE�A����< ��$�SAVG�8�6G]%���CAR �`�!�$���"CRa���$ d�#qE�@��"STD���!Fpo��'QOF0��%��"RC���&RC۠�(F�2A�R#7����%, gMA�Q_�a��
QQ��al2��%u4I��r7I�R�9�wQ�7�8M/��!C:pR�  �p�2F<�SDN�a0 �  W2QM P $Mi��s$cA �$C�cm�9���4���AT�0CY_ �N LS!IG1@x'yB��y@@H2Y��NO����SDE�VI�@ O@�$�RBT:VSP0�3�CuT�DBY|�A�	W`3CHNDGD�AP H@GRP�HE iXL�U��VSЌFx2� DL1p aQ6ROp��FB�\]�FEN�@��S���ChAR d�@DyOd�PMCS̶��P薇P�R��HOT�SWz42�DMpELE�1/e��C8`�RS T�@���r� hfl��`OL�GHA�Fxk�Fs�� �C��A@T � $�MDLUb 2S@�E���q�6�q	0�i(�c�e�cJ��	uݢ`�#~5t+w�PTO���� �byU DSLA}VS� U  ��INP �	V�ЊyA�_;�ENUAV �$R�PC_�q�2 �1bL�w�0 B�pSH=O+� W ���A�a�q�2�r�v�u�v�S_CF� X�` ,f��r�O�G gE��%D�h�J`eC�Iߣi�MA��,D�x AY?�W� p�gNTV	�D�VE�0.@�SKI��T�`g$?Ň2�� JZs�!� Cꆻ��f�_SyV/ �`XCLU��:H���ONL��'��Y�T��OT:eHI�_V,11 APPL�Y��HI4`;�U�_�ML�� $VGRFY8�	�U�M{�IOC_I���J 1�/��߃O�@X�LS�w"`@$DUMMCY4���ڑ�Cd L_TP���kC��^1CNFf���E���@T�y� D_#UQ_0��ݥ�YPCP��=� � ������uJ >�� Y +�
0�RT_;P�!�N;OCCb Z�r��TE���=�פ�DG��@[ D�P_;BAe`kc��!��_��H��Md��E \�pAb=cARGI&�!$���`[���c�_SGNA] �8�`U��IGN�Տ�,�� ��V����>��ANNUN��&��˳�EU�J'�ATCH��J���u�u^ <@g�����:c$Va����擬��1EF] I�� �_ @@FͲI}Tb�	$TOTi @�C�O�c�u�M�@NI�a`tB��c����A>���DAY@CLOAD�D\�n�������EF7�XIJ�Ra��K���O%���a�ADJ_R�!@b��>�H2�"A[�
 c�%��`a͠�MPI�J��D �A8��?�Ac 0��ѐ��� ��Z�ϡ�U|i ��CTRL� �Yp d��TRA�8 ?3IDLE_PAW  �Ѡ��Q�V�G�V_���`c ��o�;Q@e� 1q$��6`<cTAC-3@��P�LQ�Z�Rz�\ A-u:ɰSW;�A\���/J��`�b�K�OH�(OP9P; �#IRO� �"gBRK��#AB � �O������� _ ���F���`d͠, j@S�oRQDW��MS��P6X�'z��IFEgCAL�� 10^tN��V��豊�V�(0L��CP
��N� 9Yb�0FLA_#�3OVL ��HE���"SUPPO��ޑ\B�L�p��&2X�*$Y-
Z-
W-
��`/��0GR�XZ�q6�$Y2�CO�PJ�SA�X2R��*r�!���:��"~RI�0)�f{ `�@CACHE���c��0�s0LA�Z SUFFI, �C��Ja\���6�o´aMSW�g �8�KEYIMA-G#TM�@S��n�
2j�r�3 @OCVsIE��~�h �a�BGL����`�?�P@� @���i��!`STπ!�����������EMKAI�`N�����Y�'FAU� �j�"Jaa��U�3��� �}�k< $dI#�US�� �IT'��BUF`��DN�B���SUBu$�DC�_���J"��"SAV �%�"k������';�r�P�$�UORD���UP_u �%��8OT�T��_B`��8@LM0l�F4��C7AX@Cv�b��Xu 	��#_G��
 @YN_���lT6���D�E��M��U��T��F��cavC�DI`BEDT)@IC��~�m�rI�G�!"c�&��l`��-�P���FZP n (�pSV� )d\�ρ���~QA��o� �����>"$3C_R�IK��kB��hD{p�RfgE.(ADSPd~KBP�`�IIM�# �C�Aa�A��U�G��4�iCM! IP��KC��� �DTH� �S�B2*�T��CHS�3�CGBSC��� ��V�d�YVSP�#[T_DrcCONV�Grc[T� $�Fu F�ቐd�C�0�j1��SC5�e]CM�ER;dAFBCM�P;c@ETBc mp\FU DUi b��+�~�CD�Ix%P702#��EO��B�qWӏ�SQ��QǀSU��MSS�1ju�4`��T�qAa��A�1r�� "�Й��4�$ZO@s���l�U�6�&��eP���eCN�c�l��l�l�iGRO�U�W)��S c�MN�kNu�eNu�eNpR|b|�i�cH�pi��z
 �0CYC���s�w�c���zDEL�_D��RO�a���qVf���v{�O�2���1� �t��:R�ua�.#� &��AL� �1sˢI1¡�J0�PB���0�ER^�T�Gbt �,!@��5��aGI1L�cR1s 
G�ԠN	O��1u��������R�P����Cڠ	�<����DMA��J0��0vH *	�L U�1#J�Q��V
�[�7A z���z��z��z�Ѩz�Fz�7w�8w�9Pw���y���1��1��U1��1��1Ě1њU1ޚ1�2��2�����2��2��2��2�Ě2њ2ޚ2�3J��3��3����3��U3��3Ě3њ3ޚe3�4���2XTF��1w6�.(�0�f�0�U�0ŷ�e��FDR�5�xTU VE���?1���SR��REr�F���OVM~Cz)�A2�TROV2ɳDT� R�MXa�I�N2���Q�2�IND�p�r�
���0�0�0G@u1��[�G`��{�D_֎[�RIV�P��G�EAR~AIOr�K"N�0�y�p�5`�@�a�Z_MCM܀ ���F��UR��Ryǀ��!?� ��p?nЋ�?n�ER�v�=a�!��P��zI:�PXq�B�RI0%��#ET�UP2_ { ����#TDPR�%T�Bp�����Ցa�"BAC�2| T��"�4E)�:%	`^B��p�WIFI��� Mc����.�PT��!FL{UI�} � ��K UR�c!���Bp�1SPx E�EMP�p�2$��S^�?x��Jق0
3VRT|���0x$SHO��9Lq�6 ASScP=18��PӴBG_��񀐓���F�ORC��g�d~�)"FUY�1�2\�2�
A�h� p� |n��NAV�a��������S!"��$�VISI��#�SC�M4SE����:0E�V�O��$���M����$��I��@��FMR2��� �5`�r� @�� �2�I�9 �F�"�_���LI�MIT_1�dC_�LM������DGC�LF����DY�L	D����5�����ģ�� ���u	 �T�FS0Ed� �P��QC�0$E#X_QhQ1i0�PԪaQ3�5��G�oQ��� ����RS�W�%ON�PX�EBcUG��'�GRBpگ@U�SBK)qO1nL� ��POY �
)��P��M��O,Xta`SM��E�"�a����`_E � �
@��>`TERMrZ%�c&��ORI�1z_ �c' �SMep�O��_ �|)�`�(�~c%�l:�UP>� �� -��F�b���q#� ���yG�*� ELTOQ�p�0�PFIrc�1Y���P�$�$�$UFR�$��1L0Le� OTY7�PT4q��k3NST�pPA�T�q4PTHJ��a`EG`*C�p1ART� !5� y2$2�REL�:)ASHF�TR1�1�8_��R(�Pc�& � $�'@��� ��s�1 @I��0�U�R G�PA�YLO�@�qDYN_k���.b�1|��'PERV��RA��H�� g7�p�2�J�E-�J��RC���ASYM�FLTR�1WJ*7����E�ӱ1�I��aUT�pbA�5�F��5P�PlC�Q1FOR2�pM��GRI!����W��/&�0F0�bs�H��Ed� �m2XN���5`OC1!>?�$OP�����c�����bRE�PR.3�1a�F��3e��R�5e�X�1>(�e$PWR��_���@R_�S�4��et�$3UD�ҸПQ72 ����$H'�!^�`ADDR�fHL!�G�2�a�a�a��R���U�� H��SSC����e-��e���eƪ�SEE��aSC=D��� $���PE_�_ B!rP�������HTTP_���HU�� (�OcBJ��b(�$�f�LEx3Us�� G� ���ะ_���T?#�rS�P��z�K9RN�LgHIT܇5� �P���P�r������P�L��PSS<�ҴJQ�UERY_FLA� 1�qB_WEBS;OC���HW�1�U���`6PINCPU���Oh��q�����d���d���� �IHMI_ED� �T �RH�?$��FAV� d�ŁOLN
� 8�R�@$SL�iR$INPUTM_($
`��P��w ـSLA� ����5�1�8�C��BXKـ6p�F_AS7��C$L%�}w%�A��\b.1�����T@HqYķ������g�wUOP4� `y� ґ�f�¤�������`PCC
`����#��>�QIP_ME��7� Xy�IP�`�U�_NET�9����Rĳs�)��DSaP(�Op=��BG`�p����A��� l��:CTAjB�pAF T�I�-U��Y ޥ�0PmSݦBUY IDI �rF ��P��a�� �&y0�,����Ҥ��NQ�Y R��IR�CA�i� � �ěy0�CY�`EA�����񘼀�CC��¥�R�0�A�7QDA�Y_���NTVA�����$��5 ���S3CAd@��CL�����Q���𵁛8�Y��2,e�o�N_�PCP�q��ⱶ��,�N�����
�xr���:p�N� �2��Ы�(ᵁ�p���xr۠LABy1���Y ��UNIR��Ë ITY듭��e&��IR#�5����R_URL���$AL0 EN��ҭ�t� ;�T��T_U��ABKY_z��2D#ISԐ�C�Jg����P�$���E��g�R��З A�/���J����FLs��7 �Ȁ���
�UJR.� ���F{0G`��E7��J7 �O R$J8I�7���R�d�7��E�8�{�H�APHI�QS��DeJ7Jy8B��L_KE*п  �K��L}M[� � <X��XRl�u���WATCH_VA��o@DўtvFIELc��cy�U ��4� � o1Vx@��-�CT[�9�m��4 �LGH�ߣ� $��LG_SIZ�t�z�2Xy�p�y�FD��Ix� ��+!��w�\ ����v� �S���2��p�����@��\ ���A�0_g�CM]3NzU
RF Q\vv�d(u�"B��2�p����I��+ �0\ ��v�RS���0�  �ZIPDULƣ�aLN=��ސ�p�z6���f�>s�D�PLMCDAUiEAFp���Tu�GH�RE�|�BOO~�a�� C���I�IT+���`��R9E���SCR� �s���DI��SF0�`RGIO"$D������T("�t|�S�s{�Wp$|�X��JGM^'�MNCH;�|�FN���a&K�'uЅ)UF��(1@�(FWD�(H]L�)STP�*V�(�%Г(��(RS9HIP�+��C[T�# R��&p:'^9U=q�$9'��H%C𜓚"Gw)�0PO�7�*��#W}$��v�)EX��TUI�%I���Ï���rCO#8C� *�$S��a	)��B@�NOF�ANA|��Q
�AIp|�t:��EDCS�P�c�C�c�BO�HO�G�S���B�HS�H(IGN�����!O��n�DDEV<7LL��#�-��Ц(�;�T�$��2�p���T=��#A���(�`p�{�Y��POS1�U2�U3�Q���2�@��G� ��{�PtD� ���&q)��0�d�V�VSTӐR�YU��B@ ` �$E.fC.k�p<p=fPf	��4�ѩ LRТ�  ��x�c�p��<�Fp�d�_CrS�_ ������Kq&���c ��MC7� ����CLDPӐ��TRQLI#ѽ�yt�FL��,r�5s8�D�5wS�LD5ut5u�ORG��91HrCRESERV���t���t���d�� �� 	u95t5u��PITp��	xq�t�vRCLMC�������q/M��k�������$DEBUGMAS��ް��?%U8$T@��Ee�g�ޥ�MFRQՔ�� � j�HRS�_RU7��a��A<��k5FREQ� ��$/@x�OVER���n��V#�P�!EFI�%�a��g�8ǒ���t� \R�ԁ�d�$U�P��?�A��PS�P��	�߃C��͢a��U|\�l�?( 	=��MISC� d�@�QRQ��	��TB � Ȗ0A՘�AX����ؗ�EX'CESjҧ�M��\��������ԝ���S}C�P � H��̔_��Ƙǰ]���/
�MKHԳK�J�� m�B_K�FLI�C�dB�QUIR-EG3MO��O˫3���`ML�`MGմ ��`��T��F�aNDU�]��>ș�k�G�Df��IN�AUT���RSM>�a��@N�r]3-��PSTL\�� 4nX�LOC�VRI%�v�UEXɶANGuB�u�R�ODA���b�������MFO� ����Y�b@�e4�2�k�SUP�e��FX���IGG� � �A��c���cQ6 �dD�%�b|�!`��!`���|��3w�ZWa�TI���p;� M��[��[ t��MD��I�A)֟@���HݰM��DIA�����AW,!�wQ�1�D��)�O���]�� -0�CU��VP��p�u�x�!_V��ѻ ����S�X�5�������P��0N���P���KES2���-$qB� ����ND2�����2_TX�dX�TRA�C?�/��M8�|q�`�Pv��X0Ұ�Pt SBq`�U/SWCS��T��	����PULS��A�N�Sޔ��R��JOIN��H��~`j�=��b��b�����P=���$��b$���TA�����S���S�HS�E&��SCF���J��R�ƚ�PLQ�:��LOā�н.���^� ���8�������0�R�R2��� 1���eA�q d$���Iΐ+�G�A2�+/� �PRsIN�<$R �SW0"�a/�ABC�D_J%�¡u���_J3�
�1#SPܠe�u�P���3��р`u��JP/���r�qO8QIF��CSKP"z{�${�J���QLp2LBҰ_AZ�r��~ELQ��O�CMPೕ�T���R1T�����1�+��F�P1��>@�Z��SMG0��=�JG��`SCL�͵SPH_�@��%V�u�= RTER` L �< A_�@G1"�aA�@c��\$DI�n
"23UDF��}!LW�(VEL�qIN�b)@� _BL�@u��$G�q�$�'��'�%`<�� ECH<ZR/�TSA_`�K���E}`<����H5�Bu��1}`_�� �)5D2d%�A4bI��N9t&�DH�tA���ÀP$V `�#>A$��ͲV�$QS�R}�����H �$B�ELvᵆ<!_AC�CE�!c��7/��0I�RC_] ��pNyTT��S$PS�rL�d�/Es��F {�@F
��9gGCgG36B���_�Q�2�@p�A���1_MGăcDD�A]"ͲFW�`����3�EC�2�HDE>�KPPABN>G��SPEE�B�Q%_p�B�QY�Y��11$U�SE_��,`Pk�C�TReTYP�0�q P�YN��Ae�V�)хQM���ѷ��@O8� YA�TINCo�ڱ��B�DՒ�WG֑ENC����u�.A�2Ӕ+@/INPOQ�I�Be���$NT�#�%NT�23_�"ͲIcLO� Ͳ_`��I�_�if�� _�k�? �` ej�C<400fMOSI�A���ОA䃔�PERCGH  �c��B" �g ��c��lb=������oUu@�@	A�B(uL eT	~�1eT�ljgv΂fTRK@%�AY ��"sY��q�B�u�s۰p�]��RU�MOMq�ՒY�MP�^��Ca�s�CJR��DUF ��BS_BCKLSH_C�B)����f����St�H��RR��QDCLALM-d���pm0���CHK���GLRTY���d��pY��)Üd_UM]��ԉC��A!�=PLMT� _L�0��9��E�.� ��#E )�#H� =��Q3po�xPC�axHW�頿E�ׅCMCE��@�GC�N_,ND�Ζ�S	F�1�iVoR��g<!p��0r���CATގSH)�,�DfY���f��7A���܀PALބ�R_P݅�s_� �v���s����JG�T]���Y�����TORQUaP��c�yPOU��b��P%�_W�u�t��1D�P�3C��3C�IK�IY�I�3F�6�����@VC�00RQ�t���1���@ӿ��ȳJRaK�����UpDB �M��UpMC� DL�1BrGRVJ�Cĭ3Cĳ3$�H_��"�j@�q�COS~˱~�LN���µ�ĭ0���@��u����̓��Z���f$�MY��؊��|��>�THET0reNK23�3hҧ3��[CBm�CB�3C! AS� ��u��ѭ3���m�SB�3��x�GT	S$=QC������x�����$DU��@Kw�B�%(��%QqA_��a��x�{�K���b(��\�A`Չ��8p�{�{�LPH~�g�Aeg�Sµ��������@g������֚�V��QV��0��V��V��UV��V��V	�V�V%�H��������G�T����H��H��H	�UH�H%�O��O��OV	��O��O��O���O��O	�O�O�Fg���	������SPBALANC�E_-�LE��H_`�SP!1��A��|A��PFULCE`lTl��.:1���UTO_����T13T2��22N���2 9`�!�qnL�=B�3��qTXpOv 
A4�I�NSEG�2�aREqV��`aDIF�ufS91�8't"1�`COB.!t�M��w2��9`��,�LCHWA�RRCBAB�� �@�#�`-ФQ 5�X�q�PR��&��2�� �
�""��1eROB�͠CR0r5�� ���C�1_��T �� x $W�EIGH�P`$Ȝ�?3àI�Qg`IF�YQ�@LAG�Rq�S��R �RBILx5O1D�p�`V2ST�0V2P!t�W0 �01�&1
/0�30
�P�2�QA�  2řd[6DEKBUg3L_@�2�OMMY9&E Nz��D`$D_A�a�$�0��O� _�DO_@A.1� <B0�6�m�Q��B�2�0N-cdH_�p`�P
�2O�� _�� %��T`�"a��T/!�4)@TI�CKh3| T11@%�C ��@N͠�XC͠R?��Q�"�E�"�E8@_PROMP�SE~�? $IR��Qp��R;pZRMAI)�h�Q�R4U_r02S�; �q�PR8�COD��3FU�Pd6ID_�[�vU R!G_SwUFFu� l34�Q;Q�BDO�G �E�0�FGRr3�"�T �C�T�"�U�"�Uׁ�T�8D�0�B0Hb _F�I�19*cORDf�1 50�236V��+b�Q1@$ZDT�}U���1;E��4 *:!L_NA�mA�@�b�EDEF_I�h�b�F�d�E�2�F��4�F�c�E�e�FIS�P��PAKp�Ds�C��d��44בi��2DP�"�It�3D�O#>OBLOCKEz��S��O�O�Gq�R�PUM �U�b�T�c�T�e�T!r �R�s�U�c�T�d�R�6 �q�S� ���U�b�U@�c�S�Z��X�@P`  t�@qe�)@W�x����sSCH�TE|�<D�( l1�LOMB_��ɇ0�V2VIS;�ITY�V2A��O�3A_FcRI��a SIq��QR�@��@�3�3V2W��W�4���r�_e��QEAS^3��Rϡ��_�[p:R�4��5�6_3ORM_ULA_Iz���wTHR^2 �Gtg��30f��<8�5COEFF_O�A	 �$�A��GR�^3Sg0B#CAnO/C$��]3�ؠ�1GRP� � � $�p�YBX�@TM~w���u�BX�s��bCER, Ttt�sd$`�  �LLt�TSpS~�_SVNt�ߐ��$`�@��$`�� ��SETUsMEA*P�P��W0��1+b/0� � h��  @ڐo�l�o�cqz��b�@cqq	`tP�G��R�� Q�\p*q[p��>�c �NPREC>at� έ0SK_$|��� PB11_USER�e"�{ ���VEL���{ 0�$�Ҍ!I]`u�T�ACF}G���  �@z@ O�"NORE-0Xl@o�V�SI.1�d��6�"UXK�fP!���DE�� $K�EY_�3�$gJOG�� SV��`����!��}�SW�"��a\aS�ՐT|�GI���| ^�� 4� h��'d2�!XY�Zc���31�_7ERR#�� 8Ԡ�AfPV�d��1����_$BUF��X��ܴ��MOR|�� HB0CUd�lA�!���GQ\aB�,"!a	$� ���a��0_��?�G~�� � �$SIՐ���VOx��T� OBJE_���ADJU)B��EGLAY���%�DR�OU.`=ղВQ0b=��T���0���;BDIR���; I�"0DYNW�2��	T��"R���@�0�"�OPWORK����,%@SYSB9Uy�SOP��$ޑ�U�; P�pN�<�PA�t�>�"��+OP�PUd!0�`!z��l�IMAGw�1B0y�2IM�Õ��INe�d��RGO�VRD��-��o�P q��0��J�Os���"�L�pBa���o�PMGC_Ee`���1Ny M A�21�2U����SL_��� � ?$OVSL�ǫň?q�`��2�" -�_ ��k�P��k�Pu���2�C� �`�Ź����_ZER�D��$G��\��>���� @*���%MOh`RI��� 
�JP8+��=!/�L���ح�T� �0AT�US��TRC_T���sB��}fs��9s�1Re`��� DFAm����L���"��00a� ޱ��XEw{�����C0vcUP��+p	qPXPȝj�43 ���PG\���$S�UBe�%�qe9J?MPWAIT z�}%LO��F�A�R�CVFBQ�@x"�!R��� �x"ACC� R�&�B�'IGNR_{PL9DBTB�0Pqy!BWbP�$w��Uy@�%IGT�PI���TNLN�&2R���rL�NP��PE�ED \HADO!W�06�w��E[q4�jO!�`SPDV!� LbAz�`�07��3UNIr��0"!R��LYZ`� o���PH_PK��~e�RETRIE9�{�q����0'PFI�"�� �G`�0D �2�g�DBGL�V�#LOGSIZ,��EqKT�!U��VD�D�#$0_T�G�MBՐCݱ��|@eMRvC|}�3�CHECK0N���PO�V!�kЙI��LE(!��P�ArpT�2K�WӿAP�2V!� h $ARIBiR� c�a/�qO�P8�ӐATT�� 2�IF|@z�Aq4S�3�UX����PLI�2V!� $g���I�TCHx"[�W �AqS9�uULLBV!��� $BAr�DYs��BAM!h���Y9�PJ5���Q��R6�V�Q_KN�OW�Cb��U��A�D�XV��0D�+iPAYLOAt��Ic�_��Rg�RgZOcL|�q��PLCL_�� !7��b�QB�T�d���fF�iC֠P�js��d�I�hRؠH�g�ҢdB����J�¦q_J�a#���AND��Ĳ.t�b�a���r�PL0AL_ �P�0���Qր�C��DNcE���J�3CpWv� TPP�DCK������P�_�ALPHgs�sBE0��gy|�K�1>�� � ���HoWD_1Oj2ydDP�AR�*��;�&���TIA4U�5U�6��MOM��a���n�h��{�Y�B� ADa�p��n���{�PUB���R��҅n�҅{�����2�Wp��W �  �PMsbT� �BxQ���� e$PI��81��TgPJ��niJ�IV�Id�Ir��[��3!��>!���r�Ӫ�U3HIG�SU3�%�4얎4 �%� ���"����!
�<�!�%SAMP����^��_��%�P4s ю���[ 	ӝ�3  ���0���&�C�����^��Sp��H&0	�IN�SpB����뤕"���6��6�V�GAM�M�SyI�� ET�ْ��;�D�tA�
$NZpIBR!62IT�$HIِ_���C�˶E��ظAҾ���LWͽ�
���7����rЖ,0�qC�%CHyK��" �~I_A�����Rr�Rq�ܥ�Ǚ��ԥ���Ws ��$�x 1����I7RCH_5D�!� RN{��#�LE��ǒ!,��x����90MSWFL��$�SCR((100��R@��3]B��ç���a����َ0��PI�3A9�METHO�����%��AXH��XX0԰62ERI���^�3��R�0$u	D��pF{�_���?���1�L�L�_�a�OOP����wᲡ��'APP:���F���@0{���أRT�V�OBp�0T����;��� 1�I��� ��r�6��RA�@MGA1��vuTSV-��P��CURg�;�GRO<[0S_SA�Q��,Y�#NO�pC!" �tY��Zolox��������!b����&�DO�1A���A����Х� �A���A"�WS�c� �2h�*�� � ��YLH�qܧ��SrZ�]B�o�@��ĵq_�C�1��M_W���g���c�M� �`Vq�$p�x1o�3"r�PMJ�,�� �'Aȡ 9�!Wi:�$�LWQ|ai�tg�t@g�tg{t� �N`P���S��SpX�0O�s�RqZ��P� *�� ���M�������� ������X��� ��2�:�q_~R� |�q#( Y����&n��&{�Y�Z� �'�&t��Q��D�#0��qP}`�$P#Q�PMON_QUc�� � 8�@QCsOU��%PQTH��sHO�^0HYS:P3ES�R^0UEI0O�@O|T�  �0P�Gõz�RUN_T�O��0Oْ.�� PE`�5C��A<��INDE�ROG�RAnP� 2g�N�E_NO�4�5ITx��0�0INFO�1�� �Q�:A��s�AB� (��SLEQݖFAѕF@��6� OSy�T�{ 4�@ENAB�>�0PTION.S%0ERVE���G��wFwGCF�A� @R0�J$Rq�2���R��H�O�G "�ED;IT�1� �v��K�ޓʱE�N9U0W*XAUTu�-UCOPY�ِN\�����MѱNXP\[q�PWRUT9� _RN�@wOUC�$G�2|�T���$$CL`�������Q��&�� �P�S�@�Xw�PXK�Q�IRTU��_�PA�� _WRK 2 �e�@ 0  �5�QMoYh�Jo|m |l	 �`�m�o��`��o�o�f�e�l}�a0I[ct'`BS�*�� 1�Y� <7���� ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������sr;CC��LMT�P����s  dѴI�Nڿ�дPRE_EXE��)�Ƅ0`jP��za'`DV���S�@e)�%�select_macro����kϤ�>qtIOCNVVB��k ��P��US�x�w���0V 14kP $$p��a�|�`?��Ɛ >�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p ������� ���$�ѰLARMRECOV ^������LMDG ��Ь�LM?_IF ���d.TPIF-2�80 Remot�e iPenda�nt: 127.�0ހ1 logg?ed out�� � ���9�K�]�o���, 
 �	���8DEF�AULT ȗLI�NE 0ȑAUT�O ABORTE=DȘJOIN�������$���� �A����������ȯ�Ҧ��ѰNGTO�L  @� 	 A   ��Ѱ�PPINFO �� f�L�^�p����  ������ k���ۿſ�����5���Y�C�iϏ�%��� ү����������'߀9�K�]�o߁ߓߙ�P�PLICATIO�N ?t���|�Ha�ndlingTo�olȖ 
V9.40P/17�~��
8834ؒ���F0�	�549���������7DF�5�О�ȓNone���FRA�� �69��_ACoTIVE1�  ��� �  ��ސMO�D��������CH�GAPONL�� ��OUPL[�1	��� >�B�T��f���CUREQ [1
��  /�p�խ��������l��� ����������i3�l�p���^H/�A�t
HTTHKY� FXv|�� *<N`���� ����//&/8/ J/\/�/�/�/�/�/�/ �/�/�/?"?4?F?X? �?|?�?�?�?�?�?�? �?OO0OBOTO�OxO �O�O�O�O�O�O�O_ _,_>_P_�_t_�_�_ �_�_�_�_�_oo(o :oLo�opo�o�o�o�o �o�o�o $6H �l~����� ��� �2�D���h� z�������ԏ��� 
��.�@���d�v���0��������TO������DO_CLEA�N���E�NM  �� p������ɯۯv�DSPDgRYRL���HI��o�@��G�Y�k�}��� ����ſ׿�������MAX��,�呿��=�X,�<�9�<���PLUGG,�-�9���PRC��Bm�"q�6�(ϗ�O���^�SEGF�K�� �� �m��G�Y�k�}�8������LAP$�7� �������+�=�O�a�s����� �T�OTAL_ƈ� �U�SENU$�1� �������RGDI_SPMMC�d��C�O�@@�1�O�"�D��-�_STRING 1��
�M��S���
��_ITE;M1��  n��� ������ $6H Zl~��������I/O SIGNAL���Tryout� Mode��I�npNSimul�ated��Ou�t`OVER�R!� = 100���In cyc�lT��Prog� Aborj��~JStatus���	Heartbe�at��MH F�aul��Aler�!/!/3/E/W/�i/{/�/�/�/  (���(����/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO�/WORИ�~A�/ XO�O�O�O�O�O __ $_6_H_Z_l_~_�_�_�_�_�_�_�^PO ���"`�KoEoWoio {o�o�o�o�o�o�o�o /ASew��bDEV%n�p9o ����#�5�G�Y� k�}�������ŏ׏������1�C�PALT�-j��OD����� ��ȟڟ����"�4� F�X�j�|�������į֯X�GRIB���� ���6�H�Z�l�~��� ����ƿؿ���� π2�D�V�h�z�����R �-��&���������� "�4�F�X�j�|ߎߠ� �������������PREGn�W���0� ~������������ � �2�D�V�h�z���������$�$AR�G_~@D ?	������  	$�$	[]��$:	��SBN_CONFIG�X�WqRCII�_SAVE  �$zm��TCEL�LSETUP �
%  OME�_IO$$%M�OV_H� ��R�EP��#��UTOoBACK� 	�tFRA:\�D� .D�z '�`�D�w� ��s  2�5/11/29 �20:26:16D�;D���#//h��C/j/|/�/�/�/�/D�X/�/?? (?:?L?�/p?�?�?�? �?�?�?g? OO$O6O HOZO�?~O�O�O�O�O��O�O���  c_�F_\ATBCK?CTL.TM�)_�;_M___q_8INI�m��j~CMESSAG� �Qz >�[ODE_D� ��j�XO�p�_@PwAUS6` !�� ,,		� ; :oHg.ohoRoto vo�o�o�o�o�o�o`@*<v��d~`TSK  mxw}_CUPDT�P�Wd�p�VXWZD_ENB�Tf
�v�STA�U�u��X�ISX UNT 2t�vwy � 	� d�S���w�����ԏ�������.�1�ME�T��2@��y P��r����9�SCRDCFG 1;Y ��w�����%�7�I�pD�Q�	ܟ������ ϯ��Z��~�;�M� _�q�������6���F�GR9��p�_ԳPN5A� 	FѶ�_ED�P1��� 
 �%-PEDT-¿ R�v�&��Es� -FE�
D�;9/�>���/  ����2��� ��B� ����{�����j�����3��#� �G� Y���G�ߠ�6�����4������Yި�� Z�l������5K��� ����Y�t���&�8���\���6��d��Yހ@����(��7 �S0wY�w��f���8�W��{�IZ��C/��2/����9{/��//L Zݤ/?V/h/�/�/��CR���?�?Tn?��? ?2?�?V?԰!�N�O_DEL�ҲGE_UNUSE޿�дIGALLOW� 1�   �(*SYST�EM*z�	$S?ERV_GR[�@n`REG�E$�Cz��@NUM�J�C�M�PMU?@z��LAYK�z��PMPAL�PUCOYC10 N3^P<!^YSULSU_�M�5Ra�CLo_�TB�OXORI�ECU�R_�P�MPMC�NVV�P10|I^�PT4DLI�p��_�I	*PROG�RA�DPG_cMI!^Ko]`AL+e�joTe]`B�o�N�$FLUI_RE�SU9W�o�O�o�dMR�N�@�<�?�; M_q����� ����%�7�I�[� m��������Ǐُ돀���!�3�E�W�2BL�AL_OUT ��K���WD_A�BOR:PcO��IT�R_RTN  ��$�빸�NONS�TO�� lHC�CFS_UTIL� �̷CC_�AUXAXIS ;3$� h}�j��|�����ƽCE_R�IA_I`@��נ��FCFGG $�/�#��o_LIM�B2+�w �� � 	��SB\���$� 
Ԡm��)�Z�%�/������[����� !���!�����L��(a
5�����PA�`�GP 1H������A�S�e�w�6�CZC� C7��J���]��p�������W C���������U������é�̩�Uձ�ߩ�����e���;���PCk���������������J�����ɱ���������� D�W D!�!�!�m!� ��&?��{HE@ONFIp�C�G_P�P1H� +EH��ߟ߀�����������C�KoPAUS�Q1H�ף IR�S�H�A� �e���������� ����E�+�i�{�a����A?Iץ�M~ؐNFO 1�;�� �3���$ ´ � Dq�  �D	� �4  �6(�L^�O�� � ��LL/ECT_�!�����EN+`�ʒ��n�NDE�#��/�1234?567890�" �A��/ҵHw��#)j��<i{��; ��/��/`/+/ =/O/�/s/�/�/�/�/ �/�/8???'?�?K? ]?o?�?�?�?�?O�?t��$� �>�IO &��A▒O�O�O�O`G[TR�2'DM(��0^�?�NN�(oM Z���_MOR)q3)H��7ىU3��Y�_ �_�_�_�_�[bR�kQ�*H�,S�?<�<ѠD<cz�KFd���P	,��;ϒo�o�o@˿�o�oœh�UA	�@E�oA ��sja�PDB�.���4cpmidbg3��Рs:��>uqpz��vq ��>x��}�.��}�`��|�<�mgP���t��~f�������@ud�1:�?��XqDE�F -��zC)�*�cO�buf.t�xtJ��|K�[`�/zDM��>���Rl�A��MCiR20_{bRCd���hS21�1���G�ACzA�d )v�%������Я��6f23DLD�	>�z�!� 2��}���yc
�@x9µ�C���= Da I���E����  E%q��F�� E�p��u���F�P E���fF3H ��GM���A	?5�>�33H��?�xn9�q@�QG5����RpA?a�A=L��<#�QU�@���Cϒ����RSMOFST �+i�����P_Tu1Ɠ4DMA =����MODE 5�dm�@��	Q�i;��%��?����<�M>�̽Ͷ�TESTc�2i�`�R�6�O�K�ECa AB�An� 8���\�n�CdB�j��Cu @p������p:d�QS ���մ�������4�IJ7>���>B8m�5$�RT_c�P�ROG %j%�d�1�h@NUSE�R��x�KEY_T�BL  e������	
��� !"#$%&'�()*+,-./�(:;<=>?@�ABCc�GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������>��͓���������������������������������耇���������������������9�4A8�LCK��F�<y��STAT��2�=X�_ALM������_AUTO_D�O�E�FDRw 3:i�2h��AUS�x����$g ��A����� �T*g�2�  bf��/�/9/ ;�*pm�P/z/�~/h/ �/�/�/�/�/?"=� G?Y?k?/|?�?L/�? �?�/�?�?OO�?*O @OvO�O6?�O�O�O~? �O	_�?*_$_BOD_6_ p_~_T_�_�_�_�_�O o)o;o�OLoqo_�o �o�_�o�o�o�o�o�o FXo��No ���o���� @�N�$�b�x�����n ������A��b� \�z�|�n�������ʟ ���(�֏O�a�s�� ����T�ʯį��֯ ����2�H�~���>� ��ɿۿ���ϼ�2� ,�J�L�>�xφ�\Ϛ� �����Ϧ��1�C�� T�y�$Ϛߔ߲ϴߦ� ��������N�`�� ����V߼����� �����H�V�,�j� ������v����� $I��jd���v �����0�� Wi{&��\� ����/&/�:/ P/�/�/F�/�/�/� �/?�:?4?R/T?F? �?�?d?�?�?�? O�/ 'O9OKO�/\O�O,?�O �O�?�O�O�O�O�O
_  _V_h_O�_�_�_^O �_�_�O
oo"_$oo Po^o4oro�o�o�o~_ �o	�_,Q�_r l�o�~���� �&�8��o_�q���. ����dڏԏ���  �.��B�X�����N� ǟٟ럖���!�̏B� <�Z�\�N�����l��� �������/�A�S��� d���4�����¯Ŀ�� ���Կ�(�^�p�� �ϩϻ�f����Ϝ�� �*�,��X�f�<�z� �����߆����#��� 4�Y��z�t�ߔ�� ���������.�@��� g�y���6����l��� ��������(6J `��V������ )��JDbdV ��t���/� 7/I/[/l/�/<�/ �/��/�/�/?�/? 0?f?x?&/�?�?�?n/ �?�?�/OO2?4O&O `OnODO�O�O�O�O�? __+_�?<_a_O�_ |_�O�_�_�_�_�_�_  o6oHo�Ooo�o�o>_ �o�ot_�o�oo�o 0>Rh��^o ����o�1��oR� L�jl�^�����|��� Џ���?�Q�c�� t���D�����ҏԟƟ  ���"�8�n���.� ����˯v�ܯ���"� �:�<�.�h�v�L��� ��ֿ迖��!�3�ޯ D�i���τϢ��ϖ� ���ϴ����>�P��� w߉ߛ�FϬ���|��� ��
����8�F��Z� p���f�������� �9���Z�T�r�t�f� ���������� �� GYk�|�L�� ������* @v�6���~ �	/�*/$/BD/6/ p/~/T/�/�/�/�/� ?)?;?�L?q?/�? �?�/�?�?�?�?�?�? OFOXO?O�O�ON? �O�O�?�O�OO__ @_N_$_b_x_�_�_nO �_�_o�OoAo�Obo \oz_|ono�o�o�o�o �o(�_Oaso ��To���o�� ���2�H�~���> ��ɏۏ����2� ,�J�L�>�x���\��� ��������1�C�� T�y�$����������� ��į��N�`�� ������V���ῌ�� �����H�V�,�j� �϶���v����߾� $�I���j�d߂τ�v� �߾ߔ������0��� W�i�{�&ߌ��\��� ���������&���:� P�����F�������� ����:4R�TF ��d��� �� '9K��\�,� �������
/  /V/h/�/�/�/^ �/�/�
??"/$?? P?^?4?r?�?�?�?~/ �?	OO�/,OQO�/rO lO�?�O~O�O�O�O�O �O&_8_�?__q_�_.O �_�_dO�_�_�O�_�_� o.ooBoXo�otc��$CR_FDR_�CFG ;re��Q
U�D1:�W�TJ�d � �`�\�bHISoT 3<rf  �`  ?�RW@tAtBt�CqpDtEtI*tgtotw�_���bINDT_EN�6p�T��q�bT1_DO�  �U�u�sT2���wVAR 2=ֹg@qh?r ��r��r�l�R�s<4�s<�m�[��RZ�`STOP���rTRL_DEgLETNp�t ���_SCREEN �re�rkc�sc�rUw�MME�NU 1>�� / <�\%�_� �T��R��S/�U��� e�w�ğ������џ� 	�B��+�x�O�a��� ��������ͯ߯,�� �b�9�K�q������� ࿷�ɿ����%�^� 5�Gϔ�k�}��ϡϳ� �������H��1�~� U�gߍ��ߝ߯����� ��2�	��A�z�Q�c� �����������.� ��d�;�M���q�������������YӃ_?MANUAL{��r7ZCD�a?�y�r^G ���R�f�"
�"
?|(���PdTGRP 25@�yAqB� � �s��� �$DwBCO�pRIG����v�G_ERRL�OG A��Q��I[m �N_UMLIM�s���u
�PXWOR/K 1B�8����//�}DBT;B_�� C%��Ap�S"� �aDB__AWAY��Q�GCP �r=���m"_AL�F�_�Yz����p�vk � 1D� , 
��/"�/%?/(c_M�pqw,@�=5�ONTIM���f�t�_6�)
�0~�'MOTNENFp�F�;RECORDw 2J� �-?�SG�O��1�?" x"!O3OEOWO�8_O�O �?�OO�O�O�O�O�O (_�OL_�Op_�_�_�_ A_�_9_�_]_o$o6o Ho�_lo�_�o�_�o�o �o�oYo}o2�oV hz��o��C �
��.��R��K� �������Џ?��ߏ �*�����+�b�t�� ������Ο=�O��� ��:�%���p�ߟ񟦯 ��O�ǯ�]������ H�Z���������#��5����ϩ�i"TO�LERENCv$B�ȿ"� L��� C�SS_CCSCB� 2K�\0" ?"{ϰϟ���7�� 
����@�R�d�3߈���"�x�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C�Ugy��� �������R�LL]�La�m1T#2� C�C�p�F�^ A�C�%pC���#�0�? 	 A����B���?�  ��$����\0����0��B��`#sߠK/]/o/�ϓ/��/�/s/�/�/�K��K8Lg�����\1� 1�?3�Ȧ��/�Q�/`?;�@���O?�?�?�?Ȏ0A0F��?{F�A OO��7�1���9M	AB 
AZOdBAE�9$O�O�O��Oi:P��`�@0��DJCA� @5��
X-.
[N#_   M?�>O� ڴ�q_�_�_�_:W�A<o:[<ǲ/o�/�_+oPobotoL�eACHC�V�W-B$�Dz�cD�`�a =/�o�oo�oW�a.+	!��2=t,y�J? �.s�s�js�w�yj �������Q�Qs�@`��$���� �A����Bމ�o�� '�9��_]�o�N���r� ��ɟ۟_�B�ʄ���YZ>`,`:�B���B��@���=
j�1	Ĝ�Z�l�~����`_м¯��� 
���̯9�,�]�o���  �H�����ٿ뿊�� ƿ3�E�W�iϬ���$� ������ Ϟ����/� A�S߶�w�V�h߭ߌ�0�S���ߐ�_�f 	��H�?�Q�~�u�� ����������� D��-�g�q������� ������
@7�Icm��߾�  �����) M@qdv��� ����//I/P� m/�v/�/�/�/�/�/ �/�/?3?*?<?i?`? r?�?^/�?�?�?�?�? O/O&O8OJO\O�O�O��O�O�O�O�O�g	 � Q�P��s �PC4
p*p�p6U6P\�C9p/p��Q ]V^PM]�6P�:P��>P�VJ_�^P��bP�fP�Vr]v���p Q
k���_oob�id1Q&oNo ;o�_co�oˏUUA  � �o�k1Q@�  ��o�k�b�������p �� 1��b6��1C���C�cP�fL��?#�c>�/{���`�cP��@@�d��r�`BȲcP>�s�qC��p���b�t<�o�?�PH�)S�B�tq�q�p�r�`CB���eIC�&��Q�4( �oz�UU+`�; =��9��=��A��0N�*U���=��7P\�OB�x�b�<�`ځ`  ?�p�x��U�[?���}t���$���$DCS�S_CLLB2 {2M��p��P�^?�NSTCY� 2N���  ����� ��ʟ؟���� �2� D�Z�h�z�������¯�ԯ��SA�DEVI_CE 2O��!�$��4&V�h����� ��˿¿Կ���
�7� .�[�R�ϑϣϵ������4(A�HNDGDg P��*�Cz�A�LS 2Q�� _�Q�c�u߇ߙ߽߫����?�PARAM �RP��1�`�&�R�BT 2T�� �8�P<C�'p# �qi�l��s@"��R��(qI�X��y0�pB CW  ��B\x�N��Z����%��)���X�j� �p����zq�����B 	�(s,�F�p�V���q���b��B ��4&c �S�e�l�4+�����H1~���{�D�C�$Z���b���A,� 4��u@�X@���^@w���]Bߣ��B�cP%���C4�C3:_^C4��nЬ ���p8�-B�{B��A������ l��C��C3�JC4�jC3��yn+��3 Dff 2��A PB W4+@ :�]o�W��� ��/�/P/'/9/ K/]/o/�/�/�/�/? �/�/�/?#?5?�?Y? k?�?�?�o�?�?O�? 6O!OZOlOWO�O�Es �?�?�?�O�O_�O�O L_#_5_G_Y_k_}_�_ �_�_ o�_�_�_oo 1o~oUogo�o�o�o�o �owO D/Az e����O�o�o
� �o��R�)�;���_� q����������ݏ� <��%�r�I�[�m��� �����ǟٟ&�8�� \�G���k�������گ ů�����F��/� A�S�e�w�Ŀ������ ѿ�����+�x�O� aϮυϗϩϻ����� ,���b�t�ﯘ߃� �ߧ���������:� �C�U߂�Y�k��� ���������6��� l�C�U�g�y������� ���� ��	-? Q������� @+dvQ� �������*/ //%/r/I/[/�// �/�/�/�/�/&?�/? \?3?E?�?i?{?�?�? U�?�?"O4OOXOCO |OgO�O{��?�O�? �O�O0___f_=_O_ a_s_�_�_�_�_�_o �_oo'o9oKo�ooo �o�o�o�o�o�O: %^I�������H�$DCSS�_SLAVE �U���	����z_4D � 	��AR_M�ENU V	�  �j�|�������ď�B�Y�� ��~?�SH�OW 2W	� � �b�aG�Q�X� v���������П֏���� @�:�d�a�s� ���������߯�� *�$�N�K�]�o����� ��̯ɿۿ���8� 5�G�Y�k�}Ϗ϶��� ��������"��1�C� U�g�yߠϝ߯����� ���	��-�?�Q�c� ��s����������� ��)�;�M�t���� ������������ %7Ip�m���� ������!3 ZWi���J� ���//DA/S/ e/��/��/�/�/�/ �/?./+?=?O?v/p? �/�?�?�?�?�?�?? O'O9O`?ZO�?�O�O �O�O�O�OO�O_#_ JOD_nOk_}_�_�_�_ �_�O�_�_o4_.oX_ Uogoyo�o�o�o�_�o �o�ooBo?Qc u���o:����CFG X)��3�3q5p�_FRA:\!�L+��%04d.CSVj|	p}� �q[A g�CHo�zv��	����3q������́܏� ���4���JP����q�p1� �RC_O�UT Y���C��_C_F�SI ?i� .������� ͟�����>�9�K� ]���������ίɯۯ ���#�5�^�Y�k� }�������ſ���� �6�1�C�U�~�yϋ� �����������	�� -�V�Q�c�uߞߙ߫� ���������.�)�;� M�v�q������� �����%�N�I�[� m��������������� ��&!3Eni{ ������� FASe��� �����//+/ =/f/a/s/�/�/�/�/ �/�/�/??>?9?K? ]?�?�?�?�?�?�?�? �?OO#O5O^OYOkO }O�O�O�O�O�O�O�O _6_1_C_U_~_y_�_ �_�_�_�_�_o	oo -oVoQocouo�o�o�o �o�o�o�o.); Mvq����� ����%�N�I�[� m���������ޏُ� ��&�!�3�E�n�i�{� ������ß՟����� �F�A�S�e������� ��֯ѯ�����+� =�f�a�s��������� Ϳ�����>�9�K� ]φρϓϥ������� ����#�5�^�Y�k� }ߦߡ߳��������� �6�1�C�U�~�y�� �����������	�� -�V�Q�c�u������� ��������.); Mvq����� �%NI[ m������� �&/!/3/E/n/i/{/ �/�/�/�/�/�/�/3��$DCS_C_�FSO ?����71 P ??T?}? x?�?�?�?�?�?�?O OO,OUOPObOtO�O �O�O�O�O�O�O_-_ (_:_L_u_p_�_�_�_ �_�_�_o oo$oMo HoZolo�o�o�o�o�o �o�o�o% 2Dm hz������ �
��E�@�R�d��� ������ՏЏ��� �*�<�e�`�r����� ����̟�����=��8�J�\�������?C/_RPI4>F?�� �����3?�&�o�X���� >SLү@d� �����%�7�`�[� m�Ϩϣϵ������� ���8�3�E�W߀�{� �ߟ����������� �/�X�S�e�w��� ����������0�+� =�O�x�s��������� ����'PK ]o������ ��(#5Gpk }�����Q��� /6/1/C/U/~/y/�/ �/�/�/�/�/?	?? -?V?Q?c?u?�?�?�? �?�?�?�?O.O)O;O MOvOqO�O�O�O�O�O �O___%_N_I_[_ m_�_�_�_�_�_�_�_ �_&o!o3oEonoio{o �o�o�o�o�o�o�o FASe������>�NOCO�DE ZU���?�PRE_?CHK \U��p�A �p�< ��pU�]�o�U� 	 <Q������ ��ۏ�Ǐ�#���� Y�k�E�����{�şן ��ß����C�U�/� y�����s���ӯm��� 	���?��+�u��� a�������ɿ�Ϳ߿ )�;��_�q�K�}ϧ� �������ω���%��� �[�m�Gߑߣ�}߯� �߳����!���E�W� 1�c��g�y������ �������A�S�-�w� ��c����������� ��+=asM_ ������' �]o	�� ����/#/�G/ Y/3/e/�/i/{/�/�/ �/�/?�/?C?9K y?�?%?�?�?�?�?�? 	O�?-O?OOKOuOOO aO�O�O�O�O�O�O�O )_____q_K_�_�_ a?�_�_�_�_o%o�_ Io[o5oGo�o�o}o�o �o�o�o�o�oEW 1{�g���_� ���/�A��M�w� Q�c����������Ϗ �+���a�s�M��� ������ߟ���'� ��3�]�7�I������ ɯۯ�������G� Y�3�}���i���ſ�� ������1�C���+� yϋ�eϯ��ϛ����� ����-�?��c�u�O� �߫߅ߗ�������� )��M�_�U�G��� A������������� I�[�5����k����� ��������3E Q{q���]� ���/Aew Q������� /+//7/a/;/M/�/ �/�/�/�/��/?'? ?K?]?7?�?�?m?? �?�?�?�?O�?5OGO !O3O}O�OiO�O�O�O �O�O�/�O1_C_�Og_ y_S_�_�_�_�_�_�_ �_o-oo9oco=oOo �o�o�o�o�o�o�o __M_�ok�o �������� I�#�5����k���Ǐ ��ӏ��׏�3�E�� i�{�5c���ß��� ��ӟ�/�	��e�w� Q�������ѯ㯽�ϯ �+��O�a�;����� ���Ϳ߿y���� !�K�%�7ρϓ�mϷ� �ϣ���������5�G� !�k�}�W߉߳ߩ��� ���ߕ��1���g� y�S�������� ���-��Q�c�=�o� ��s��������� ����M_9��o �����7 I#mYk�� ����!/3/)/ i/{//�/�/�/�/�/ �/�/?/?	?S?e??? q?�?u?�?�?�?�?O O�?%OOOE/W/�O�O 1O�O�O�O�O__�O 9_K_%_W_�_[_m_�_ �_�_�_�_�_o5oo !oko}oWo�o�omO�o �o�o�o1Ug AS������ 	����Q�c�=��� ��s���Ϗ�o���� ��;�M�'�Y���]�o� ��˟����۟�7� �#�m��Y������� �����!�3�ͯ?� i�C�U�������տ� ������	�S�e�?� �ϛ�uϧ��ϫϽ�������$DCS_SGN ]	��E��-����29-NOV-�25 20:27� ��N� x�x�� [}�t��q��т�xҚك�JѨ��EƼÞ� �ۈǖ�  1�HO�W ^	�� x�/�VE�RSION �=�V4.5.�2��EFLOGI�C 1_���  	�����C���R�%�PROG_E_NB  ��:��{�s�ULSE  �X��%�_AC�CLIM������d��WRSTgJNT��E��-�EMO|�zя�$���INIT `2�����OPT_S�L ?		�	�
 	R575��V]�74b�6c�7c�50��1���C��|�@�TO  L��� �V�DEXҞ�dE�x�PA�TH A=�A�\k}��HCP�_CLNTID y?�:� D���ռ��IAG_G�RP 2e	�����z�	 �@�  
ff�?aG���BG�  2��/�8�[I@c�ς!��7@�z�@^��@
�!���mp2m15 �89012345�67���� � ?��?��=q?��
?���R?�Q�?ѯ�?�����?(�?�z����x�@�  A_�A�p !7A�8�8_�B4�� ��L�x�
�@����@��\@~��R@xQ�@q���@j�H@c��
@\��@U�@Mp��//�'$�; �O)H���@Ct >d 9���@4�/\)@)�� #t {@��/�/�/�/�/P'�?���?����_ ?}p�?u?n{?s ;?\�Q�? ?�2?D?V?h8�
=?�����0w5�z��H?p�h��?^�R�?�?�?�?��?h8��t0����@�?��0� ;@&O8OJO\OnOP' �$_�_Y_k_�O?_ �_�_�_�_�_s_�_�_ 1oCo!ogoyoo�o���Bj"� �2{1�@"?���f�t0�d"�5!�
u4V��u"�B3t�A>u��U?@[q��@`,�=q�=b���=�E1>�J��>�n�>��H�"<�o �z�s��q��� �x�C��@<(�Uz� �4�� ����A@x�?*�o��m*� P�b���tn���2����Ώ�����i>J���&�bN2�"�'�G�N��o@�@v�奈0����@f�fr!l ��33����(��"C��� ƒI�CH��)C.dB؃�"8"����' ���"~�A?�&"K���,�pf�B��@�p�� �����p�Ľ�ϯ�x� �����0��N�T� ��e�=�������̿�� �ۿ���A*B��!��o��CT_CON�FIG f�|�|�egY���STBF_TTS��
����О�}�:��1�MAU����~��MSW_CF���g�  # ��OCoVIEW��h!�-����s߅ߗߩ� ���ߟ�a�����,� >�P���t����� ��]�����(�:�L� ^�������������� k� $6HZ�� ~������y  2DVh��������v�RC�i���!��/ S/B/w/f/�/�/�/���SBL_FAUL�T j*6��!G�PMSK���'��TDIAG k���-�������UD1: 6789012345I2��=1���%P\υ?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�Od6�96�I�r
t?�O|�TORECP"?4:
B4 4_[77[s?p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�O�O�O��o7�UMP_OP�TIO=��.�aT�R����)uPM�E��Y_TEM�P  È�3�BC�gp�B�QtU�NI����gq�YN_BRK lL�~7�EDITOR�a��a@�r_
PENT� 1m)  ,&�/��d�3�8� "�_�F���j������� ݏď����7��[� m�T���x�������� ҟ����E�,�i�P� ������ï���������A�(��pMGDI_STAzuV�gq��uNC_INFO� 1n!��b����X���������n�1o!� ��o���
�
�d�oU�g�y� �ϝϯ���������	� �-�?�Q�c�u߇ߙ� �߽��� u����
�� *�B�*�P�b�t��� �����������(� :�L�^�p��������� 2�������9�C Ugy����� ��	-?Qc u�������� //1;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?��?�?�?O)/O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�?�?�_ �_o�_3O=oOoaoso �o�o�o�o�o�o�o '9K]o�� ��_�_����+o 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y��������ӟ ���	�#�-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� �7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߹��� �������%�/�A�S� e�w��������� ����+�=�O�a�s� �������������� �'9K]o�� ������# 5GYk}�	�� ����/1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?��?�?�?�? /O)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�? �_�_�_�_O�_!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew��_�_��� �o�+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o���� ���ɟ۟���#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� ���߹���������� %�7�I�[�m���� �����������!�3� E�W�i�{��߇����� �����/AS ew������ �+=Oas ����������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?���?�? �?�?��?OO1OCO UOgOyO�O�O�O�O�O �O�O	__-_?_Q_c_ u_�?�_�_�_�_�?�_ oo)o;oMo_oqo�o �o�o�o�o�o�o %7I[m�_u� ���_���!�3� E�W�i�{�������Ï Տ�����/�A�S� e��������u�� ����+�=�O�a�s� ��������ͯ߯�� �'�9�K�]�w����� ����ɿ�����#� 5�G�Y�k�}Ϗϡϳ� ����������1�C� U�g߁��ߝ߯���ۿ ����	��-�?�Q�c� u����������� ��)�;�M�_�y߃� ������������ %7I[m�� �����!3 EWq�c����� ����////A/S/ e/w/�/�/�/�/�/�/ �/??+?=?O?i{ �?�?�?�?��?�?O O'O9OKO]OoO�O�O �O�O�O�O�O�O_#_ 5_G_�?s?}_�_�_�_ �?�_�_�_oo1oCo Uogoyo�o�o�o�o�o �o�o	-?Qk_ u����_��� ��)�;�M�_�q��� ������ˏݏ��� %�7�I�cQ������ ���ٟ����!�3� E�W�i�{�������ï կ�����/�A�[�� �$ENETM�ODE 1p����  
k�k�f�����j��OATCFG �q�����Ѵ��C���DAT�A 1rw�Ӱ�.��*	�*��'�9�K�]�l�dlύ�e��ϻ�������� �'ߡϳ�]�o߁ߓ� �߷�1���U����#� 5�G�Y����ߏ��� ��������u��1�C� U�g�y������)��� ����	-����c�u�����j�RPOST_LO��	t�[
׶#5�Gi�RROR_P-R� %w�%L��XTABLE  w�ȟ�����RSEV_NUM� ��  ����  �_AUT�O_ENB  ����X_NO5! �uw���" W *�x �x �x 	�x + +w �/�/�/�Q$FLTR=/O&H�IS#]�J+_A�LM 1vw� e�[x,e�+�/�Q?c?u?�?�?�?�/_\"W   w�v!����:j�TCP_V_ER !w�!x޻?$EXT� _R�EQ�&�H)BCSsIZKO=DSTKhI�f%�?BTOL�  ]Dz�"��A =D_BWD��0�@�&�A���CDI�A wķ���]�KSTEP�O�Oj�>POP_DO�Oh��FDR_GRP s1xw��!d 	�?x�_��yPs�Y�Q�'�M"����l��T� ����VyS�_�] �_o�_&ooJo5ono�Yoko�o�o�o�j?��L%@&��?���?o"�n
 F@]�a�o ���3:�o^I�mxyAp�u@S33�uh}@�q�g��yP�q��|yPG�  �@�Fg�fC�8RL��}?��`i��~�6�X����87�5t��5����5`+��������n[PEATUROE y���@���Handl�ingTool ��]Engl�ish Dict�ionary�4�D St��ard���Analog� I/O>�G�gle ShiftZ��uto Soft�ware Upd�ate�mati�c Backup����ground� Edit ��C_ameraU�FY��CnrRndIm����ommon �calib UI���nˑ�Monoitor$�tr�?Reliabn���DHCP �[�at�a Acquis�3�\�iagnos���R�v�ispla�yΑLicens�Z�`�ocument Viewe?��^�ual Che�ck Safet�y��hance�d���s�Fr�ܐ�xt. DI�O /�fi��@�e�nd�Err>�L(��\�4�s[�rP�K�� �@
�FCTN /Menu��vZ����TP In��faycĵ�GigE־��Đp Mask� Exc�g=�H�T԰Proxy �Sv��igh-wSpe�Ski��� Ť�O�mmuni�c��onsV�ur໰��q�V�ײcon�nect 2��n{crְstru!�$�ʴ�eۡ��J����KAREL Cmod. L�ua�~��Run-Ti<��Env�Ȟ�el u+��s��S/W��ƥ���r�Book�(System)�
�MACROs,~M�/Offseu��p�HO���o�u�MR�8�4���MechStop+�t����p�im�q���x�R������odo�witc�h�ӟ�.��4�O�ptmF��,�fi�l䬳�g��p�ul�ti-T�Γ�P?CM fun�Ǽ��o��������Regeie�rq���riݠ�F���S�Num �Sel��/�:� Adjua�*�W�q�h�tatu��ߪ��RDM Robo}t�scove'���ea��<�Fre�q Anlyq�Rem��O�n5�����ServoO�!��?SNPX b-�v�;SN԰Cliܡ?r�Libr&�_��Q ��q +oJ�t���ssag���@ 0����	�@/Iս��MILIB��P� Firm���Pλ�AccŐ͛TPsTXk��eln���������orq}uo�imula=�4�|u(�Pa&���ĐX�B�&+�ev.̸��ri��TU�SB port ��iPf�aݠ&R� EVNT� n?except�����%5��VC�rl�c���V���"�%4q�+SR SCN�/gSGE�/�%UI	�?Web Pl��>���A43��ۡ��ZDT Applj�<
�{1EOAT�����&0?�7Gridp�񾡬=�?iR�"�.5� F���/גRX-10iA/L�?�Alarm Caouse/��ed(��All Smoo�th5���C�sciyi+�V�Load�ΌJUpl�@w�to�S ��rityA_voidM(�s7�1t�@�ycn��0���_�CS+���g. c��XJo� ��-T3_H�.RX��U����Xcollabo����RA�:�.9����in���N�RTHI
�On��e Hel����ֿ������1trU�ROS Eth$��A� �����;,�G �B�,|HUpV�%�W�3t ԰�_iRS�ݐ��64MB DRsAM�o�cFRO8���L8F FlD���d��2M �A:�opm�bԕex@V�
�sh�qD��wce�u��p��|tyn�sA�
�%�Ar����J��^�.v� P)Q/sbS�`���8O�N��mai��U����R�q�T1��^FC+Ԍ%̋Fs�9�ˌk̋��Typ߽FC%�hױV�N Sp�ForްK��Ԇ��lu!����cp�P'G j�֡�RJ�[L`Sup"}���֐f��crFP��lu� ��al�����r��i�
q�4@�ް�uest,IMPLE ׀6*|H�Z���c0�BTeap(�|���$rtu���V�9HMI�¤��wUIFc�pono2D��bC�:�L�y�p� ��������ʿܿ	� � �?�6�H�u�l�~ϫ� �ϴ���������;� 2�D�q�h�zߧߞ߰� �������
�7�.�@� m�d�v������� �����3�*�<�i�`� r��������������� /&8e\n� �������+ "4aXj��� �����'//0/ ]/T/f/�/�/�/�/�/ �/�/�/#??,?Y?P? b?�?�?�?�?�?�?�? �?OO(OUOLO^O�O �O�O�O�O�O�O�O_ _$_Q_H_Z_�_~_�_ �_�_�_�_�_oo o MoDoVo�ozo�o�o�o �o�o�o
I@ Rv����� ����E�<�N�{� r�������Տ̏ޏ� ��A�8�J�w�n��� ����џȟڟ���� =�4�F�s�j�|����� ͯį֯����9�0� B�o�f�x�����ɿ�� ҿ�����5�,�>�k� b�tφϘ��ϼ����� ���1�(�:�g�^�p� �ߔ��߸������� � -�$�6�c�Z�l�~�� �����������)� � 2�_�V�h�z������� ��������%.[ Rdv����� ��!*WN` r������� //&/S/J/\/n/�/ �/�/�/�/�/�/?? "?O?F?X?j?|?�?�? �?�?�?�?OOOKO BOTOfOxO�O�O�O�O �O�O___G_>_P_ b_t_�_�_�_�_�_�_ oooCo:oLo^opo �o�o�o�o�o�o	  ?6HZl�� �������;� 2�D�V�h�������ˏ ԏ���
�7�.�@� R�d�������ǟ��П �����3�*�<�N�`� ������ï��̯��� �/�&�8�J�\����� ������ȿ�����+� "�4�F�Xυ�|ώϻ� ����������'��0� B�T߁�xߊ߷߮��� ������#��,�>�P� }�t��������� ����(�:�L�y�p� �������������� $6Hul~�����  ?H552���21R785�0J614AwTUP'545'�6VCAMC�RIbUIF'2�8cNRE52�VR63SCH�LIC�DOC�V�CSU86�9'02EIOC��4R69VEgSET?UJ7U�R68MASK^PRXY{7OCO#(3?+ �&3j&J6%53��H�(LCHR&O�PLG?0�&MH�CRS&S�'MCS�>0.'552MD�SW+7u'OPu'M�PRv&��(0&PCMzR0q7+ 2l� �'51J51�8�0JPRS"'69�j&FRDbFRE�QMCN93�&SNBA��'SHLBFM1G�8�2&HTC>TMsIL�TPA�oTPTXcFELF�� �8J9�5�TUTv'95�j&UEV"&UEC�R&UFRbVCC�
XO�&VIPnFC;SC�FCSG���IWEB>HTT>R6��H;RV�CGiWIGQWIP�GS�VRCnFDGvu'H7�7R66J�5'R�8R51*
(6�(2�(5V�)J8�86�L=I%� �84g662R�64NVD"&R�6�'R84�g79ڎ(4�S5i'J7�6j&D0�gF xR�TSFCR�gCR�Xv&CLIZ8IC�MS�Sp>STY:nG6)7CTO>���7�NNj&ORqS�&C &FCB��FCF�7CH>F�CR"&FCI�VF�C�'J�PO7GBfMv�8OLaxENDS&�LU�&CPR�7L�WS�xC�STxT�E�gS60FVmR�IN�7IHaF �я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� !3EWi{� ������ /ASew��� ����//+/=/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]? o?�?�?�?�?�?�?�? �?O#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �_�_�_�_�_	oo-o ?oQocouo�o�o�o�o �o�o�o);M _q������ ���%�7�I�[�m���������Ǐُ��  H55�2��21�R7�8�50�J61�4�ATUP7�5�457�6�VCA�M�CRI��UI�F7�28��NREv�52v�R63�wSCH�LICƚ�DOCV�CSU��8697�0F�E�IOCǛ4�R6=9v�ESETW�u��J7u�R68�M�ASK�PRXY���7�OCO��3�W����6�3�J6�5�536�H$�LC�HƪOPLGW�0^�MHCRǪS���MCSV�0��55�F�MDSW���OP��MPR���6��06�PCM��R0`E˓�F���6�51f��51��0f�PRSv��69�FRD���FREQ�MCN��936�SNBA�כ%�SHLB�M�E��ּ26�HTC�V�TMIL�6�T{PAV�TPTX��#ELړ�6�8%�#���J95��TUTv��95�UEV��wUECƪUFR���VCCf�O��VI�P��CSC��CS�Gƚ$�I�WEBnV�HTTV�R6՜���S���CG��IG���IPGS'�RC���DG��H7��RK66f�5�u�R��WR51f�6�2�I5v�#�J׼��6���LU�5�s�v�4��6�6F�R64�NV�D��R6��R84֦79�4��S5n�J76�D0u�FRTS&�CR�CRX��CLI&�e�CMSV�sV��STY��6�CT�OV�#�V�75�NN��ORS����6�F�CBV�FCF��C�HV�FCR��FC-IF�FC��J#�˵G
M��OL�E�NDǪLU��CPUR��Lu�S�C$��StTE�S60n�FVRV�IN��IH���m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s�@��������͏ߏ��STD�LANG���0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰����RBT
�OPTN������'�9�K� ]�o�����������DPN	���)� ;�M�_�q��������� ������%7I [m����� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	-?Qcu� �������� )�;�M�_�q������� ��ˏݏ���%�7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w� ��������ѿ���� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� ������1�C�U�g� y���������������@	-?Qc�f�������9�9��$FEAT�_ADD ?	����  	�#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������DEMO y?   �L� B�T߁�xߊ߷߮��� ��������G�>�P� }�t��������� ����C�:�L�y�p� �������������� ?6Hul~� �����; 2Dqhz��� ��� /
/7/./@/ m/d/v/�/�/�/�/�/ �/�/?3?*?<?i?`? r?�?�?�?�?�?�?�? O/O&O8OeO\OnO�O �O�O�O�O�O�O�O+_ "_4_a_X_j_�_�_�_ �_�_�_�_�_'oo0o ]oTofo�o�o�o�o�o �o�o�o#,YP b������� ���(�U�L�^��� ��������ʏ��� �$�Q�H�Z���~��� ����Ɵ����� � M�D�V���z������� ¯ܯ��
��I�@� R��v���������ؿ ����E�<�N�{� rτϱϨϺ������ ��A�8�J�w�n߀� �ߤ߶��������� =�4�F�s�j�|��� ����������9�0� B�o�f�x��������� ������5,>k bt������ �1(:g^p ������� / -/$/6/c/Z/l/�/�/ �/�/�/�/�/�/)? ? 2?_?V?h?�?�?�?�? �?�?�?�?%OO.O[O ROdO�O�O�O�O�O�O �O�O!__*_W_N_`_ �_�_�_�_�_�_�_�_ oo&oSoJo\o�o�o �o�o�o�o�o�o "OFX�|�� �������K� B�T���x�������ۏ ҏ����G�>�P� }�t�������ןΟ�� ���C�:�L�y�p� ������ӯʯܯ	� � �?�6�H�u�l�~��� ��Ͽƿؿ����;� 2�D�q�h�zϔϞ��� �������
�7�.�@� m�d�vߐߚ��߾��� �����3�*�<�i�`� r������������ �/�&�8�e�\�n��� ��������������+ "4aXj��� �����'0 ]Tf����� ���#//,/Y/P/ b/|/�/�/�/�/�/�/ �/??(?U?L?^?x? �?�?�?�?�?�?�?O O$OQOHOZOtO~O�O �O�O�O�O�O__ _ M_D_V_p_z_�_�_�_ �_�_�_o
ooIo@o Rolovo�o�o�o�o�o �oE<Nh r������� ��A�8�J�d�n��� ����яȏڏ���� =�4�F�`�j������� ͟ğ֟����9�0� B�\�f�������ɯ�� ү�����5�,�>�X� b�������ſ��ο�� ��1�(�:�T�^ϋ� �ϔ��ϸ������� � -�$�6�P�Z߇�~ߐ� �ߴ���������)� � 2�L�V��z���� ��������%��.�H� R��v����������� ����!*DN{ r������� &@Jwn� ������// "/</F/s/j/|/�/�/ �/�/�/�/???8? B?o?f?x?�?�?�?�? �?�?OOO4O>OkO bOtO�O�O�O�O�O�O�__0]   'XF_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o o&o8oJo\ono�o�o �o�o�o�o�o�o" 4FXj|��� ������0�B� T�f�x���������ҏ �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ����������
��.�  /�)�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?V?h?z?�?�? �?�?�?�?�?
OO.O @OROdOvO�O�O�O�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|� �������� 0�B�T�f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�\�n� ���������������� "4FXj|� ������ 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<N `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������P ��$�4�8�+� N�`�r߄ߖߨߺ��� ������&�8�J�\� n����������� ���"�4�F�X�j�|� �������������� 0BTfx�� �����, >Pbt���� ���//(/:/L/ ^/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?l? ~?�?�?�?�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�o&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�`�r����������� ����&8J\ n������� �"4FXj| �������/ /0/B/T/f/x/�/�/ �/�/�/�/�/??,? >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO ^OpO�O�O�O�O�O�O��O __$_6Y�$F�EAT_DEMO�IN  ;T��fP�<PNTIND�EX[[jQ�NPI�LECOMP �z����Q�iRIU�PSETU�P2 {�U~�R�  N �Q��S_AP2BCK� 1|�Y  #�)7Xok%�_8o<P�P&oco9U�_�o o�oBo�o�oxo�o 1C�og�o��, �P�����?� �L�u����(���Ϗ ^�󏂏�)���M�܏ q������6�˟Z�؟ ���%���I�[��� �����D�ٯh���� ��3�¯W��d���� ��@�տ�v�Ϛ�/� A�пe����ϛ�*Ͽ� N���r���ߨ�=��� a�s�ߗ�&߻���\� �߀��'��K���o� ��|��4���X����� ��#���G�Y���}�� ����B���f������1�Y�PP�_ 2>�P*.VR8���*��������l PC���OFR6:�2�V�TzPz�w�]PG���*.Fo/��	�:,q�^/�STMi/ �/ /�-M/�/�H�/?�'?�/�/g?�GIFq?�?�%��?D?V?�?�JPG �?O�%O�?�?oO�
#JSyO�O��5C�O�MO%
JavaS�cript�O�?C�S�O&_�&_�O %�Cascadi�ng Style SheetsR_���
ARGNAMOE.DT�_��� �\�_S_�A�T�_�_>�PDISP*�_���To�_�QLaZoo�CLLB.ZIXwo2o$ :\�a\�o��i�AColla�bo�o�o
TPEINS.XMLƱ_:\![o�QCu�stom Too�lbarbiPA?SSWORDQo��?FRS:\�d�B`Passwor�d Config ���/��(�e��� �����N��r��� ��=�̏a������&� ��J���񟀟���9� K�ڟo�������4�ɯ X��|���#���G�֯ @�}����0�ſ׿f� �����1���U��y� �ϯ�>���b���	� ��-߼�Q�c��χ�� �߽�L���p��ߦ� ;���_���X��$�� H�����~����7�I� ��m���� �2���V� ��z���!��E��i {
�.��d� ���S�w p�<�`�/� +/�O/a/��//�/ 8/J/�/n/?�/�/9? �/]?�/�?�?"?�?F? �?�?|?O�?5O�?�? kO�?�OO�O�OTO�O xO__�OC_�Og_y_ _�_,_�_P_b_�_�_ o�_oQo�_uoo�o �o:o�o^o�o�o) �oM�o�o��6 ��l��%�7�� [����� ���D�ُ h�z����3�,�i� �������ßR��v�������$FIL�E_DGBCK �1|������ < ��)
SUMMA�RY.DG!�͜�MD:U���ِ�Diag Sum�mary����
C?ONSLOG��n����ٯ���Con�sole log����	TPACC�N�t�%\������TP Accou�ntin;���F�R6:IPKDM�P.ZIPͿј
��ϥ���Exception"�ӻ���MEMCHECKЏ�������-�Me�mory Dat�a����&n )��RIPE�~ϐ��%ߴ�%�� Packet L:����L�$�c���S�TAT��߭�� %A�Sta�tus��^�	FTAP����	��/��mment TB�D2�^� >I)ETHERNEw��
�d�u�﨡Et�hernJ�1�fi�guraAϩ��DCSVRF&����7����� verify all:�����4��DIFF/��'���;�Q�diff��r�d���CHG01������`A����it�2���270���fx�3���I ��p�VTR�NDIAG.LS�u&8���� �Ope��L� ��n�ostic��/�)VDEV�DAT�������Vis�Dev�ice�+IMG@��,/>/�/:�i$�Imagu/+U�P ES/�/FORS:\?Z=���Updates OListZ?��� �FLEXEVEN���/�/�?���1 ?UIF EvM�M����-vZ)CRSENSPK�/�˞�\!O���C�R_TAOR_PE�AKbOͩPSRB?WLD.CM�O͜�E2�O\?.�PS_ROBOWELS���:GIG��@_�?|d_��GigE�(�O��N�@�)>UQHADOW__D_�V_�_��Shad�ow Changye����	dt�R?RCMERR�_�_��_oo��4`CFG� Erroro t�ailo MA��k�CMSGLIBgoNo`o�o|R�e���z0ic�o�a�)�`ZD0_O�osn��ZD�Pad��l �RNOTI��Rd���Notific����,�AG��P�ӟt� ��������Ώ]��� ��(���L�^�폂�� ����G�ܟk� ���� 6�şZ��~������ C�د�y����2�D� ӯh��������¿Q� �u�
�ϫ�@�Ͽd� v�Ϛ�)Ͼ���_��� ��ߧ�%�N���r�� �ߨ�7���[����� &��J�\��߀��� 3����i����"�4� ��X���|������A� ����w���0��= f�����O� s�>�bt �'�K��� /�:/L/�p/��/ �/5/�/Y/�/ ?�/$? �/H?�/U?~??�?1? �?�?g?�?�? O2O�? VO�?zO�OO�O?O�O cO�O
_�O._�OR_d_ �O�__�_�_M_�_q_ oo�_<o�_`o�_mo �o%o�oIo�o�oo �o8J�on�o�� 3�W�{�"�� F��j�|����/�ď�֏e������0��$�FILE_FRS�PRT  ��������?�MDONLY� 1|S�� �
 �)MD:�_VDAEXTP.ZZZ1�⏹�ț�6%NO �Back fil�e ���S�6P �����>��K�t��� ��'���ί]�򯁯� (���L�ۯp������ 5�ʿY�׿ Ϗ�$ϳ� H�Z��~�Ϣϴ�C� ��g���ߝ�2���V� ��cߌ�߰�?����� u�
��.�@���d�������C�VISBC�Kq�[���*.V�D����S�FR:�\��ION\DA�TA\��v�S��Vision VD���Y�k���� y��B�����x��� 1C��g���, �P����? �Pu�(�� ^��/��M/� q/�/>/�/6/�/Z/�/ ?�/%?�/I?[?�/?�?�?2?D?�?9�LU�I_CONFIG7 }S����; $ �3U�/O�AOSOeOwO�O�Ov�$ |x�?�O�O�O_ _%\�OH_Z_l_~_�_ '_�_�_�_�_�_o�_ 2oDoVohozo�o#o�o �o�o�o�o
�o.@ Rdv���� ����*�<�N�`� r��������̏ޏ�� ���&�8�J�\�n��� �����ȟڟ쟃��� "�4�F�X�j������ ��į֯����0� B�T�f����������� ҿ�{���,�>�P� b����ϘϪϼ����� w���(�:�L�^��� �ߔߦ߸�����s� � �$�6�H���Y�~�� �����]������ � 2�D���h�z������� ��Y�����
.@ ��dv����U ��*<�` r����Q�� //&/8/�\/n/�/ �/�/;/�/�/�/�/? "?�/F?X?j?|?�?�? 7?�?�?�?�?OO�? BOTOfOxO�O�O3O�O �O�O�O__�O>_P_ b_t_�_�_/_�_�_�_ �_oo�_:oLo^opo��o�o$h  x��o�c�$FLUI�_DATA ~�����a�(a�dRESU_LT 3�ep �T���o "4FXj|�� �����(a"� 4�F�X�j�|�������@ď֏�����?(`0�0`�e?�Q��0ou��������� ϟ����)�;�M� �d�w���������ѯ �����+�=�O�(b�`O�u�3���W��� ο����(�:�L� ^�pςϔϦϷ����� �� ��$�6�H�Z�l� ~ߐߢ�a��߅��ߩ� � �2�D�V�h�z�� ������������� .�@�R�d�v������� ������������9 ����r����� ��&8J	� n������� �/"/4/F/g/) �/�/a�/�/�/�/? ?0?B?T?f?x?�?�? [�?�?�?�?OO,O >OPObOtO�O�OW/�/ {/�O�O�/_(_:_L_ ^_p_�_�_�_�_�_�_ �_�?o$o6oHoZolo ~o�o�o�o�o�o�o�O �O�OA_hz� ������
�� .�@��_d�v������� ��Џ����*�<� �o1��U��̟ ޟ���&�8�J�\� n�����Q���ȯگ� ���"�4�F�X�j�|� ����_�q���忧�� �0�B�T�f�xϊϜ� �������ϣ���,� >�P�b�t߆ߘߪ߼� �����߱�ÿտ7��� ^�p��������� �� ��$�6���G�l� ~���������������  2D�e'� K�����
 .@Rdv��� ����//*/</ N/`/r/�/�/U�/y �/�??&?8?J?\? n?�?�?�?�?�?�?�? �O"O4OFOXOjO|O �O�O�O�O�O�O�/	_ �/-_�/�Of_x_�_�_ �_�_�_�_�_oo,o >o�?boto�o�o�o�o �o�o�o(:�O [_�Uo��� � ��$�6�H�Z�l� ~���Oo��Ə؏��� � �2�D�V�h�z��� K�o��㟥
�� .�@�R�d�v������� ��Я⯡���*�<� N�`�r���������̿ ޿������5���\� nπϒϤ϶������� ���"�4��X�j�|� �ߠ߲���������� �0����%χ�I� ������������,� >�P�b�t���Eߪ��� ������(:L ^p��S�e�w�� �� $6HZl ~�������� / /2/D/V/h/z/�/ �/�/�/�/�/��� +?�R?d?v?�?�?�? �?�?�?�?OO*O� ;O`OrO�O�O�O�O�O �O�O__&_8_�/Y_ ?}_??�_�_�_�_�_ �_o"o4oFoXojo|o �o�_�o�o�o�o�o 0BTfx�I_ �m_��_���,� >�P�b�t��������� Ώ���o��(�:�L� ^�p���������ʟܟ ����!���Z�l� ~�������Ưد��� � �2��V�h�z��� ����¿Կ���
�� .��O��sυ�I��� ����������*�<� N�`�r߄�C��ߺ��� ������&�8�J�\� n��?ω�cϭ���� ���"�4�F�X�j�|� �������������� 0BTfx�� ���������) ��Pbt���� ���//(/��L/ ^/p/�/�/�/�/�/�/ �/ ??$?�� {?=�?�?�?�?�?�? O O2ODOVOhOzO9/ �O�O�O�O�O�O
__ ._@_R_d_v_�_G?Y? k?�_�?�_oo*o<o No`oro�o�o�o�o�o �O�o&8J\ n�������_ �_�_��_F�X�j�|� ������ď֏���� ��o/�T�f�x����� ����ҟ�����,� �M��q�3������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~�=���a��υ����� � �2�D�V�h�zߌ� �߰����ߓ���
�� .�@�R�d�v���� ������������� N�`�r����������� ����&��J\ n������� �"��C�gy =������/ /0/B/T/f/x/7�/ �/�/�/�/�/??,? >?P?b?t?3}W�? �?��?OO(O:OLO ^OpO�O�O�O�O�O�/ �O __$_6_H_Z_l_ ~_�_�_�_�_�?�?�? �_o�?DoVohozo�o �o�o�o�o�o�o
 �O@Rdv��� �������_�_ �_oo�1o������̏ ޏ����&�8�J�\� n�-������ȟڟ� ���"�4�F�X�j�|� ;�M�_��������� �0�B�T�f�x����� ����������,� >�P�b�tφϘϪϼ� �ύ������կ:�L� ^�p߂ߔߦ߸����� �� ��ѿ#�H�Z�l� ~������������ � ���A��e�'ߌ� ������������
 .@Rdv���� ����*< N`r1��U��y� ��//&/8/J/\/ n/�/�/�/�/�/��/ �/?"?4?F?X?j?|? �?�?�?�?��?�	O ��?BOTOfOxO�O�O �O�O�O�O�O__�/ >_P_b_t_�_�_�_�_ �_�_�_oo�?7o�? [omo1_�o�o�o�o�o �o $6HZl +_������� � �2�D�V�h�'oqo Ko�����o���
�� .�@�R�d�v������� ��}�����*�<� N�`�r���������y� Ï����ӏ8�J�\� n���������ȿڿ� ���ϟ4�F�X�j�|� �Ϡϲ���������� ˯ݯ��c�%��ߜ� ������������,� >�P�b�!φ���� ��������(�:�L� ^�p�/�A�Sߵ�w��� �� $6HZl ~���s����  2DVhz� ���������/�� ./@/R/d/v/�/�/�/ �/�/�/�/?�?<? N?`?r?�?�?�?�?�? �?�?OO�5O�YO /�O�O�O�O�O�O�O �O_"_4_F_X_j_{O �_�_�_�_�_�_�_o o0oBoTofo%O�oIO �omO�o�o�o, >Pbt���� {_����(�:�L� ^�p���������woُ �o���o��6�H�Z�l� ~�������Ɵ؟��� ��2�D�V�h�z��� ����¯ԯ���
�ɏ +��O�a�%������� ��п�����*�<� N�`���ϖϨϺ��� ������&�8�J�\� �e�?��߳�u����� ���"�4�F�X�j�|� ����q�������� �0�B�T�f�x����� ��m߷ߑ�����, >Pbt���� �����(:L ^p������ � /��������W/ ~/�/�/�/�/�/�/�/ ? ?2?D?V?z?�? �?�?�?�?�?�?
OO .O@OROdO#/5/G/�O k/�O�O�O__*_<_ N_`_r_�_�_�_g?�_ �_�_oo&o8oJo\o no�o�o�o�ouO�O�O �o�O"4FXj| ��������_ �0�B�T�f�x����� ����ҏ�����o)� �oM�t��������� Ο�����(�:�L� ^�o���������ʯܯ � ��$�6�H�Z�� {�=���a�ƿؿ��� � �2�D�V�h�zό� �ϰ�o�������
�� .�@�R�d�v߈ߚ߬� k��ߏ��߳���*�<� N�`�r������� �������&�8�J�\� n��������������� ������CU�| ������� 0BT�x�� �����//,/ >/P/Y3}/�/i �/�/�/??(?:?L? ^?p?�?�?�?e�?�? �? OO$O6OHOZOlO ~O�O�Oa/�/�/�O�O �/ _2_D_V_h_z_�_ �_�_�_�_�_�_�?o .o@oRodovo�o�o�o �o�o�o�o�O�O�O�O K_r����� ����&�8�J�	o n���������ȏڏ� ���"�4�F�X�) ;��_ğ֟���� �0�B�T�f�x����� [���ү�����,� >�P�b�t�������i� {���￱��(�:�L� ^�pςϔϦϸ����� �ϭ���$�6�H�Z�l� ~ߐߢߴ��������� ���߿A��h�z�� �����������
�� .�@�R�c�v������� ��������*< N�o1�U�� ��&8J\ n���c���� �/"/4/F/X/j/|/ �/�/_�/��/��/ ?0?B?T?f?x?�?�? �?�?�?�?�?�O,O >OPObOtO�O�O�O�O �O�O�O�/_�/7_I_ Op_�_�_�_�_�_�_ �_ oo$o6oHoOlo ~o�o�o�o�o�o�o�o  2D_M_'_q �]_����
�� .�@�R�d�v�����Yo ��Џ����*�<� N�`�r�����U�y ßퟯ�&�8�J�\� n���������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ迧��� ˟ݟ?��f�xϊϜ� ������������,� >���b�t߆ߘߪ߼� ��������(�:�L� ��/ϑ�Sϸ����� �� ��$�6�H�Z�l� ~���Oߴ���������  2DVhz� �]�o�����
 .@Rdv��� ������/*/</ N/`/r/�/�/�/�/�/ �/�/�?�5?�\? n?�?�?�?�?�?�?�? �?O"O4OFOW?jO|O �O�O�O�O�O�O�O_ _0_B_?c_%?�_I? �_�_�_�_�_oo,o >oPoboto�o�oWO�o �o�o�o(:L ^p��S_�w_� �_��$�6�H�Z�l� ~�������Ə؏ꏩo � �2�D�V�h�z��� ����ԟ查�� +�=��d�v������� ��Я�����*�<� ��`�r���������̿ ޿���&�8���A� �eϏ�Q��������� ���"�4�F�X�j�|� ��M������������ �0�B�T�f�x��I� ��mϷ������,� >�P�b�t��������� ������(:L ^p������ ������3��Zl ~������� / /2/��V/h/z/�/ �/�/�/�/�/�/
?? .?@?�#�?G�? �?�?�?�?OO*O<O NO`OrO�OC/�O�O�O �O�O__&_8_J_\_ n_�_�_Q?c?u?�_�? �_o"o4oFoXojo|o �o�o�o�o�o�O�o 0BTfx�� �����_��_)� �_P�b�t��������� Ώ�����(�:�K� ^�p���������ʟܟ � ��$�6��W�� {�=�����Ưد��� � �2�D�V�h�z��� K���¿Կ���
�� .�@�R�d�vψ�G��� k��Ϗ�����*�<� N�`�r߄ߖߨߺ��� �ߝ���&�8�J�\� n���������� ����1���X�j�|� �������������� 0��Tfx�� �����, ��5��Y�E��� ���//(/:/L/ ^/p/�/A�/�/�/�/ �/ ??$?6?H?Z?l? ~?=�a�?�?��? O O2ODOVOhOzO�O �O�O�O�O�/�O
__ ._@_R_d_v_�_�_�_ �_�_�?�?�?�?'o�? No`oro�o�o�o�o�o �o�o&�OJ\ n������� ��"�4��_ooy� ;o����ď֏���� �0�B�T�f�x�7�� ����ҟ�����,� >�P�b�t���E�W�i� ˯�����(�:�L� ^�p���������ʿ�� ۿ ��$�6�H�Z�l� ~ϐϢϴ����ϗ��� ���߯D�V�h�zߌ� �߰���������
�� .�?�R�d�v���� ����������*��� K��o�1ߖ������� ����&8J\ n�?����� �"4FXj| ;��_������/ /0/B/T/f/x/�/�/ �/�/�/��/??,? >?P?b?t?�?�?�?�? �?��?�O%O�/LO ^OpO�O�O�O�O�O�O �O __$_�/H_Z_l_ ~_�_�_�_�_�_�_�_ o o�?)OOMowo9O �o�o�o�o�o�o
 .@Rdv5_�� ������*�<� N�`�r�1o{oUo��ɏ �o����&�8�J�\� n���������ȟ�� ���"�4�F�X�j�|� ������į�������� �ݏB�T�f�x����� ����ҿ�����ٟ >�P�b�tφϘϪϼ� ��������(���� �m�/��ߦ߸����� �� ��$�6�H�Z�l� +ϐ����������� � �2�D�V�h�z�9� K�]߿�������
 .@Rdv��� �}���*< N`r����� �����/��8/J/\/ n/�/�/�/�/�/�/�/ �/?"?3/F?X?j?|? �?�?�?�?�?�?�?O O�?O/cO%/�O�O �O�O�O�O�O__,_ >_P_b_t_3?�_�_�_ �_�_�_oo(o:oLo ^opo/O�oSO�owOyo �o $6HZl ~�����_�� � �2�D�V�h�z��� �����o㏥o�� �@�R�d�v������� ��П������<� N�`�r���������̯ ޯ���ӏ���A� k�-�������ȿڿ� ���"�4�F�X�j�)� �Ϡϲ���������� �0�B�T�f�%�o�I� �߽��������,� >�P�b�t����� {�������(�:�L� ^�p���������w߉� �߭���6HZl ~������� ��2DVhz� ������
// ������a/#�/�/�/ �/�/�/�/??*?<? N?`?�?�?�?�?�? �?�?OO&O8OJO\O nO-/?/Q/�Ou/�O�O �O_"_4_F_X_j_|_ �_�_�_q?�_�_�_o o0oBoTofoxo�o�o �o�oO�o�O�O, >Pbt���� �����':�L� ^�p���������ʏ܏ � ���o3��oW� ~�������Ɵ؟��� � �2�D�V�h�'��� ����¯ԯ���
�� .�@�R�d�#���G��� k�m������*�<� N�`�rτϖϨϺ�y� ������&�8�J�\� n߀ߒߤ߶�u��ߙ� �����4�F�X�j�|� ������������� ��0�B�T�f�x����� ������������� ��5_!���� ���(:L ^������� � //$/6/H/Z/ c=�/�/s�/�/�/ ? ?2?D?V?h?z?�? �?�?o�?�?�?
OO .O@OROdOvO�O�O�O k/}/�/�/_�/*_<_ N_`_r_�_�_�_�_�_ �_�_o�?&o8oJo\o no�o�o�o�o�o�o�o �o�O�O�OU_| �������� �0�B�T�ox����� ����ҏ�����,� >�P�b�!3E��i Ο�����(�:�L� ^�p�������e���ܯ � ��$�6�H�Z�l� ~�������s�տ���� �� �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ���������ſ'�� K��r������� ������&�8�J�\� ߀������������� ��"4FX�y ;�_�a��� 0BTfx�� �m����//,/ >/P/b/t/�/�/�/i �/��/?�(?:?L? ^?p?�?�?�?�?�?�? �? O�$O6OHOZOlO ~O�O�O�O�O�O�O�O �/?�/)_S_?z_�_ �_�_�_�_�_�_
oo .o@oRoOvo�o�o�o �o�o�o�o*< N_W_1_{�g_� ����&�8�J�\� n�������coȏڏ� ���"�4�F�X�j�|� ����_q����� �0�B�T�f�x����� ����ү������,� >�P�b�t��������� ο���ß՟�I� �pςϔϦϸ����� �� ��$�6�H��l� ~ߐߢߴ��������� � �2�D�V��'�9� ��]���������
�� .�@�R�d�v�����Y� ��������*< N`r���g�������	�$FMR�2_GRP 1���� ��C4  B�.��	 ��9K^6F@ a@��6G�  �Fg?�fC�8R�y�?�  ��66��X���875�t��5���5�`+�yA�  �/+BH�w-%@'S339%�5[/l-6@6!�/xl/�/ �/�/�/?�/&??J?�5?G?�?k?�?��_�CFG �T�K�?�? OO�9NO� 
F0�FA K@�<RM_C�HKTYP  ���$&� RO=Ma@_MINg@��W���@�R X�SSB�3�� 7�O���C�O�O�5TP_D�EF_OW  ��$WIRCO�Mf@_�$GENOVRD_DO�F���E]TH��D �dbUdKT_ENB�7_ KPRAVC���G�@ �@Y�O�_�?oyo�&oI* �QOU*�NAIRI<�@��oGo��o�o�o��C�/� /��O<��q�+sL�i�O�PSM�T��Y(�@
t��$HOSTC�21���@��� 5	�x�{������e,�]�o� ������K�ď֏��������	anonymous!�O�a�s����� ����� �9���(�:�L�^��� ��������ʯ�#�5� �$�6�H�Z�����ş ןٯƿ����� � 2�y�V�h�zόϞ��� ��	�����
��.�u� ����v߭Ϛ�῾��� ����;��*�<�N�`� �߄��Ϩ�������� 7�I�[�m�o�I��߀� ������������� "4W����|�� ����/��C0 w�Tfx��G� ���/a>/P/ b/t/�/����/ /9?(?:?L?^?� �?�?�?�?�?�/#/5/ O$O6OHOZO�/�/�/ �/�?�O?�O�O_ _ 2_y?V_h_z_�_�O�_ �?�_�_�_
oo��q�ENT 1�hk� P!�_no  �p\o�o�o�o�o�o �o�o�o:_" �F�j���� �%��I��m�0��� T�f�Ǐ��돮��ҏ 3���,�i�X���P��� t�՟��៼�
�/�� S��w�:���^�������������ܯ=� �?QUICC0J�&��!192.16?8.1.10c�X�A1��v�8��\�2��ƿؿ9�!ROUgTER:��!���a��PCJOG|��e�!* ���0��U�CAMPRT�϶�!������RTS���x� !�Softwar�e Operat�or Panel�U߇���7kNAME� !Kj!RO�BO����S_CF�G 1�Ki ��Auto�-started^�DFTP�Oa� �O�_���O�������� ��E_�.�@�R�u�c� 	�����������cN:� L�^�;r���R�� ������% H�[m��� jO|O�O�O4!/hE/ W/i/{/�/T�/�/�/ �/�//�//?A?S?e? w?�?����??�? </O+O=OOO?sO�O �O�O�O�?`O�O__ '_9_K_�?�?�?�?�O �_�?�_�_�_o#o�O GoYoko}o�o�_4o�o �o�o�of_x_�_ g�o��_���� �o��-�?�Q�tu� �������Ϗ�(: L^`�2��q����� ������ݟ���%� H�ʟ[�m�������� ��� �ί4�!�h�E� W�i�{���T���ÿտ �
�Ϟ�/�A�S�e��w����_ERR ���ڇϗ�PDU�SIZ  �^�6����>��WR�D ?(���� � guest���+�=�O��a���SCD_GR�OUP 3�(� u,�"�IFT��w$PA��OMP��w ��_SH�޻ED�� $C��C�OM��TTP_A�UTH 1���� <!iPen�danm�x�#�+!�KAREL:*8x���KC�������VISION SET��(�����?�-�W�R���v� �����������������G�CTRL �Ҧ�a�
�?FFF9E3���FRS:DEF�AULT�F�ANUC Web Server�
 tdG����/�� 2DV��WR_�CONFIG ]���������IDL_CPU�_PC� �B����� BH�MI�N����GNR_�IO������ȰH�MI_EDIT {���
 ($/ C/��2/k/V/�/z/�/ �/�/�/�/?�/1?? U?@?y?d?�?�?./�? �?�?�?OO?OQO<O uO`O�O�O�O�O�O�O��O__;_�NPT_SIM_DO��*NSTAL_oSCRN� �\�UQTPMODNT�OL�Wl[�RTY�bX�qV�K�ENB�W�ӭOLNK 1�����o%o�7oIo[omoo�RMA�STE��Y%O�SLAVE ���ϮeRAMCAC�HE�o�ROM�O_�CFG�o�S�cUO�'��bCMT_O�P�  "��5sYCL��ou� _ASG s1����
 �o �������"� 4�F�X�j�|����kwrWNUM����
�b�IP�o�gRTRY�_CN@uQ_USPD��a��� �bp�b��n��M���ڰP}T?��k ��._������ɟ۟ ퟈S���)�;�M�_� q� �������˯ݯ� ~��%�7�I�[�m��� �����ǿٿ����� !�3�E�W�i�{�
ϟ� ���������ψϚ�/� A�S�e�w߉�߭߿� ��������+�=�O� a�s���&������ ������9�K�]�o� ����"����������� ����GYk}� �0���� �CUgy��, >���	//-/� Q/c/u/�/�/�/:/�/ �/�/??)?�/�/_? q?�?�?�?�?H?�?�? OO%O7O�?[OmOO �O�O�ODOVO�O�O_ !_3_E_�Oi_{_�_�_ �_�_R_�_�_oo/o Ao�_�_wo�o�o�o�o �o`o�o+=O �os�����\ n��'�9�K�]�� ��������ɏۏi�c��_MEMBERS� 2�:�_   $:� ���v���1����RCA_ACC �2���   [}�Q� �Zl������  l�l���+�  d����������a�BUF�001 2�n�=� �L l����u0  u0���
��
��
���
��
��
��
��Z
��
��R�R�U!R�-R�8R�FR�}QR�X9�  �� ������ϯ���� )�;�M�_�q���������˿��2�����B�2X�
�� �!��)��1��9� �A��I��Q�
�X� ]�a�]�i�]�q�]�y� ]�]�]����� ����������,�>� P�b�t߆ߘߪ߼���ؿ�3������� ��!�/��1�?�� A�O��Q�_�f�a�o� f�q��f⁢��f③ �����������%� 7�I�[�m���������������e�CFG ;2�n� 4l��
l�l�<��47]�HIS钜n�� �� 20�25-11-29l� �����������  Ii�;B��� r������� //K]J/\/n/�/ �/�/�/�/�/�/#/5/ "?4?F?X?j?|?�?�? �?�?�/?�?OO0O BOTOfOxO�O�O�?�? �?�O�O__,_>_P_ b_t_�_�O�O�_�_�_ �_oo(o:oLo^oL	 ��[m�o�o�o�o@�o!3!.a< �_�_������ �	��-�dv�u� ��������Ϗ��� �N�`�M�_�q����� ����˟ݟ�&�8�%� 7�I�[�m�������� ǯ������!�3�E� W�i�{�����֯诬� �����/�A�S�e� w�eoR�Ѐo�o�o�� �����"�4�F�X�! w߱�ÿ�Ͽ������� ��+�=�O�ߘߪ� ������������ '�9�p��o������� ����������H�Z� GYk}���� �� 21CU gy�����
 	//-/?/Q/c/u/��/�/��taI_CF�G 2��� H�
Cycle �Time�Bu{sy�Idl�"^�min�+1�Up�&�R�ead�'DoYw8? 2�#�Count�	N'um �"����<���c1qaPROG��"�������(/softpa�rt/genli�nk?curre�nt=menup�age,153,1�/
OO.O@O4b5�leSDT_ISO�LC  ��� ��@�.J23_D�SP_ENB  �vK0�@INC ���M�Ä@A  � ?�  =�̟�<#�
�A�I:�o �A__��X�O<_�GOB�0C�C�5�FVQG_GR�OUP 1�vK{<��d<�P�C��_D_?��?�_��Q�_o.o@o�_ dovo�o�o�,_NY�G_IN_AUT�OcT�MPOSRE�^_pVKANJI_�MASK v�HqR�ELMON ��˔?��y_ox������.6r�3��7ĲC���u�o�DKCwL_L�`NUM�@��$KEYLOGOGING�����Q��E�0LANGUA_GE ��~���DEFAUgLT ����LG�!���:2���x��@�  80H�  ���'0h� +
������GOUF� ;��
��(�UT1:\��  �-�?�Q�h�u����������ϟ�����(�g4�8i�N_DISP ��O8�_��_��LOCTOL����Dz�0A�A���GBOOK ����d�1
�
�۠X����#�5�G�Y�`i���3{�W�	��@쉞QQJ¿Կ1���_BUFF 2�NvK ���25�
�ڢVB&�7 C�ollaborativ�=�OΗώ� �ϲ���������'�� 0�]�T�fߓߊߜ��?DCS ��9�B �Ax�����%�-�?�|Q���IO 2���� ���Q� ������������ �*�<�N�b�r����� ����������&�:e�ER_ITMsNd�o����� ��#5GYk }����������hSEV��M.dTYPsN�c/pu/�/
-�aRST5����SCRN_FLW 2�s��0��� �/??1?C?U?g?�/�TPK�sOR"��NGNAM�D��~�N�UPS_ACR� ��4DIGI�8~+)U_LOAD[P�G %�:%-�INST_PAT�H�@Dt?�EMAXUALRM2��1����E
ZB�1_PD�5�0 ��y�Z@CY��˭�O+���ۡ�D�|PP 2�˫ ��	R/_
_C_._ g_y_\_�_�_�_�_�_ �_�_oo?oQo4ouo `o�o|o�o�o�o�o�o )M8qTf �������%� �I�,�>��j����� Ǐُ�����!��� W�B�{�f�������՟ ����ܟ�/��S�>� w���l�����ѯ��Ư ��+��O�a�D����p���RHDBGDEF ��E�ѱO���_LDXDISA��0�;c�MEMO_{AP�0E ?�;
 ױ��3�EπW�i�{ύϟϱ�Z@F�RQ_CFG ���G۳A ��@i��Ô�<��d%��� ������B��K���*i�/k� **:tҔ�g� y�ߔ��߱������� ���J�Es�J `d�����,(H� ��[�����@�'�Q� v�]����������������*NPJIS�C 1��9Z� � �����ܿ������	Zl_MSTR� �#-,SCD 1�"͠{� �������/ /A/,/e/P/�/t/�/ �/�/�/�/?�/+?? O?:?L?�?p?�?�?�? �?�?�?O'OOKO6O oOZO�O~O�O�O�O�O �O_�O5_ _Y_D_i_ �_z_�_�_�_�_�_�_ o
ooUo@oyodo�o �o�o�o�o�o�o�?*cN�MK����;љ$M�LTARM���:N��r ��հ���İMETPU���zr��CND�SP_ADCOLx%�ٰ0�CMNTF� 9�FNb�f�7�FSTLI��x�4 �;ڎ�s��|��9�POSCF��=q�PRPMe���STD�1�; 4�#�
v��qv� ����r��������̟ ޟ ���V�8�J��� n���¯�������9��SING_CHK�  ��$MODA���t�{�~2��DEV 	�	�MC:f�HSI�ZE��zp�2�TA�SK %�%$�12345678�9 ӿ�0�TRI�G 1�; l ĵ�2ϻ�!�bϻ��YP����H�1�E�M_INF 1��N�`)AT?&FV0E0g����)��E0V1&�A3&B1&D2�&S0&C1S0}=��)ATZ��2��H6�^���Rφ��A�߶�q�������� ��5������� ��B߳��������� ��1�C�*�g��,�� P�b�t������R� ?���u0��� ������������M  q���Z�� �/�%/��[/  2�/�/h�//�/ �/�3?�/W?>?{?�? @/�?d/v/�/�/O�/ /OAOx?eO?�ODO�O�O�O�O_�NITO�RÀG ?z�  � 	EXEC�1~s&R2,X3,X4�,X5,X��.V7,X8
,X9~s'R�2�T+R �T7R�TCR�TOR�T[R �TgR�TsR�TR�T�R��S2�X2�X2�X2��X2�X2�X2�X2��X2�X2h3�X3�X37R2�R_GRP_SV 1���� (�  �����OMO��_D��B���cION_D�B<��@�zq  K�zp%U�1u$:{��zpU��@N ��: U�-ud1�����8��PG_JOG ��ʏk�
�2�`�:�o�=���?����0�B��~\�n�������k0H�?��C�@�ŏ׏����  ������qL_NAME �!ĵ8��!�Default �Personal�ity (fro�m FD)qq1�R�MK_ENONL�Y�_�R2�a 1��L�XLy�8�gpl d�� ��şן�����1� C�U�g�y��������� ӯ���	��n�
�<� N�`�r���������̿޿� :��)� ;�M�_�qσϕϧϹ� ��������%�7�I� [�m�ߑߣߵ����� �����!�3�E�W�i� {������������ ��/�A�S�e�w��� ������������+��<�Sew� ������^��A�a��B�Bw��Pf�� ����/!/3/E/ W/i/{/�/�/�/�� �/�/??/?A?S?e? w?�?�?�?�?�?�?�? �/�/+O=OOOaOsO�O �O�O�O�O�O�O__�'_9_&O�S^Q�(x_�]�rd�d�_�^ �_�_�W���k�o.ooRog Fhqogo yo�o�o�o�o�oE`�ph"|��Fe	`[o Ugy8qK�A\��8��s� A ��y�@h�Q�Q��"����Tk\$�� W ��P�PE�x?C�  �I�@o a�<o��p�������ߏ 
f�Q,������0��P�Cr� � �3r �.� @D��  A�?�G�-�?x.I�.@I�A�����  ;�	l�Y�	 �X?  ������� �, ǀ �����̀K��o�����]K���K]�K	�.��w�r_	��̀@
�)�b�1������I�Y������T;fY�{{S���3�����I�>J���;Î?v߮>��=@�����E�΂ѯעZ����wp��u�� D�!�3��7pg  �  �9��͏W���	'� �� u�I� ��  ��u��:��È��È=�s�ͱ�E�@��@ǰ�3��{3�E��&���N�pC�  'AY�&�Z�i�b�@f��i�n�C����I�Ch����b��r����B�p�Ŕq��0�}ر�.DzƏ<����`�K�pߖ߁�݀������� 4P����.9z��d  �Pؠ??�ff�_��	�� 2p>�P��18.f�t�>L���$U���(.��P�����������É��� xށ�;e�m��K�Z;�=g;�4�<<����%��G��3����p?f7ff?ذ?&S����@=0e�?��q��y�rN�Z���I� ��G���7���(����� !E0iT��0���x��F�p� ��#��D��w ������� //=/(/a/L/�/p/ ��/�p�6�/Z#? �/ ?Y?k?}?��?�? >?�?�?�?�?�?1O��"���KD�y{CO�O8O�O���ذO�OX�O�O�y���J���}�DD1���.�D���@�AmQa��9N,���A;�^@���T@|j@$��?�V�>�z��ý��=#��
>\)?���
=�G�-]��{=���,���C+��Bp����P��6��C98R���?N@���(��5�-]G�p�Gsb��F�}�G�>�.E�VD�K�n���I��� F�W�E���'E���D���;n���I���`E�G���cE�vmD���-_�oQ_�o�o�o  �o$H3X~i �������� �D�/�h�S���w��� �����я
���.�� R�=�v�a�s�����П ����ߟ��(�N�9� r�]���������ޯɯ ۯ���8�#�\�G��� k�������ڿſ��� "��F�1�C�|�gϠ� ���ϯ���������P=(�Q34�] �����Q�	�9�Oߵ53�~�mm��aҀ5qQ�߫�aғ���<�ߵ1������ـ1��U�C�y�g��%P�P���!�/��'����
���.������4�;�t�_������� ��������:%���/�/d��� �����7 %[Im���0y27�  B�S@,J@�CH#PzS@�0@ZO/1/C/U/g/y/�-�#��/�/�/�/��/�3?�3�� @*�35�0�0�!q3��5
 ? f?x?�?�?�?�?�?�? �?OO,O>OPO�Z@1� ���ۯ�c/��$MR_CAB�LE 2ƕ�/ ��TT��& �ڰO���O�Y�@���C _���_O_u_7_I_ _�_�_�_�_�_o�_ �_oKoqo3oEo{o�o �o�o�o�o�o�o�o�Gm/�K!�"�� �O����ذ�$��6���*Y�**} �COM ȖI�����"W�'%% 2345?678901����! ��Ï��� � !5� �!
���M�not segnt b��W���TESTFE�CSALGR  eg)
!d[�41�Y
k�������$�pB���������� 9�UD1:\ma�intenanc?es.xmlğ��  C:�D?EFAULT�,�B�GRP 2�z� � ��(D;  ��%!1st cl�eaning o�f cont. �v�ilatio�n 56��ڧ�!0�����+B��*�`����+��"%���mech��cal� check1�  �k�0u�|��ԯ����Ϳ߿��@���rollerS�e�w�ū��m���ϣϵ�@�Bas�ic quarterly�*�<�ƪ,\�)�;�M�_�q�8�cMJ��ߓ "8��!� ���ߕ ��� ��+�=��C�g��ߋ���߹���������@�Overghau�ߔ��?�C x� I�P����@}���������� $n� �����aIl�ASe w������ � +=O�s� ������/R �9/�(/��/�/�/ �/�//�/�/N/#?r/ G?Y?k?}?�?�/�?? ?�?8?OO1OCOUO �?yO�?�?�O�?�O�O �O	__jO?_�O�Ou_ �O�_�_�_�_�_0_o T_f_;o�__oqo�o�o �o�_�oo,oPo% 7I[m�o��o�o ����!�3�� W��������ÏՏ �6����l����e� w���������џ�2� �V�+�=�O�a�s� �����ͯ���� '�9���]�������� ��ɿۿ���N�#�r� ��YϨ�}Ϗϡϳ��� ���8�J��n�C�U� g�yߋ��ϯ������ 4�	��-�?�Q��u� �����ߞ�������� �f�;�������� ���������P��� t�I[m���� ��:!3E W�{��� � ��//lA/�� w/��/�/�/�/�/X*�"	 X�/?.?@?�)B a/o?�?�?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_�_�_�_�_��_	oo" Џ!?�  @�!  M?HoZolo�&4o�o�oܽo�(*�o** F�@ i!k&�` o'9�o]o�����/^&�o� ����/�A�S�e� ��#�����я��� ��+�q�����7��� ����k�͟ߟ��I� [���K�]�o���C������ɯ��o$�!��$MR_HIST� 2�g%#�� �
 \7"$ 23�45678901P3�;���b2�90/ ����[���./���� ǿٿF�X�j�!�3ρ� ����{��ϟ����� B���f�x�/ߜ�S��� �߉��߭��,���P��t��=��$�S�KCFMAP  ]g%&��b�
�� ����ON?REL  �$#�������EXCFE�NB�
����&�F�NC-��JOGO/VLIM�d#�v���KEY�y���_PAN������RUNi�y����SFSPDTY�PM����SIGN|��T1MOTk�����_CE_G�RP 1�g% ��+�0�ow�#d� �����& �6\�7y� m���/�4/F/ -/j/!/t/�/�/�/{/��/�/�/?�+��QZ_EDIT
�����TCOM_CFG 1���0�}?�?��? 
^1SI 	�N����?�?��!�?$O����?XO~78T_ARC_*��X�T_MN_oMODE
�U:�_SPL{O;�UA�P_CPL�O<�N�OCHECK ?��� ��  _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo���NO_WAITc_L	S7> NTf1�����%��qa_7ERRH2��������?o�o�o�o��POGj�@O�cӦm�| �^GO  �´)<���?����t��n�bPA�RAM�b����t^�8
�.�@� = n�]�o�w� Q�����������Ϗ0�)��7�[�m�� �����ODRDS�P�C8�OFFS?ET_CARI0�O�ǖDISԟœS_�A�@ARK
T9O�PEN_FILE���1T6�0OPT?ION_IO�����K�M_PRG %��%$*����'��WO��N�s�ǥ�� ���u����	 a����Ӧ������RG_DSBL  ����jN���RIENTTO�e��Csp��A ���U�@IM_DS����r��V��LCT �{mP2ڢ�3̹���dҩ��_PEX��@���RAT�G �d8��̐UP Sװ�:����Sϰe�Kωϗ��$�r2�G�L�XL;Ț�l㰂� ������'�9�K�]� o߁ߓߥ߷�������@���#�5�G���2�� v�������������e�B�T�f� x��������������� ,>Pbt� ������ (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? �q1�~?�?�?�?�?�?��?�?O O2ODO�yA�a�tn?~M��~O�OhrP�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�O�Oo$o 6oHoZolo~o�o�o�o �o�o�o�o �_o Vhz����� ��
��.�@�R�d�QOES������B�d�ӏ�ʏ���������Y�D�}�0� �r���������ԟڟ����p���=�M��q�	`��������c�:�o�¯ԯ�|���A�  ��k�C�C�ڰ"ڰ����O��  ���-���)�?C�  �t�k� ��g�����Կ��ѿ
�`5���6z�ĳ�OU����
��
��H��n�� ۷ ^�\� �@D�  p�?��v�\�?:px�:qC4�r�p�(��  ;��	l��	 ��X  ������� �, � ��������Hʪ�����H���Hw�z/H���ϝ�x8�B���B�  X���`�o�*��3����t�>u���fC{ߍ���:pB\�
��{�9:qK�t�� ����$���\*��� DP�^���b�g  �  �h�����)�	'� � ���I� �  ���'�=���8����t�@���� !�b��6{b�t�U��(�N��r�  'D��E�C�И�t�C������ߗ���jA�@�����%�B�� ��`,���H:qDz�k�ߏz���������?А 4P���":uz:���	f��??�ff'�&8� ]�m�18:p��>L���$��$�(:p�P��	�������:� xް;e�m"�K�Z;�=g;�4�<<���E/T�v��b���?f7ff?�?&� )��@=0�%?��%8y��}!��$�x� �/v��/f'��W,?? P?;?t?_?�?�?�?�? �?�?O�?(OOLO�/ �/�/EO�OAO�O�O�O �O_�O_H_3_l_W_ �_{_�_�_1��_A��� eO+o�ORooOo�o�o �oK/�o�omo�o* '`+�,�zt��;CL�H��}?�����
��)����u����D1�/n�t��p�q���@I�h~,ȴ�A;�^@��T�@|j@$��?�V�n�z��ý��=#�
�>\)?��
�=�G�����{=��,��C�+��Bp�����6��C98�R���?}p��(��5���G�p�Gsb��F�}�G�>.�E�VD�K�L����I�� �F�W�E��'�E���D��;�L����I��`�E�G��c�E�vmD��� \�՟��ҟ���/�� S�>�w�b�������ѯ �������=�(�:� s�^���������߿ʿ �� �9�$�]�Hρ� lϥϐϢ��������� #��G�2�W�}�hߡ� ���߰��������
� C�.�g�R��v��� ������	���-��Q� <�u�`�r��������������'M�(��34�]O!����8h~�%3~��m����5Q8�������!���  `@N�r��	eP@"	P��Q�_/V/�9/$/]/H)���� c/j/�/�/�/�/�/�/ �/!??E?0?i?T?"&`�_�_�?�?�8��? �?O�?OBO0OfOTO��OxO�O�O�O�O2<f?_  B��pyp�$QCHR�z�p@ �N_`_r_�_�_�_�]c�O�_�_oo+of?�Bc� @�d4�Q8Jc�D
 2o�o �o�o�o�o�o%�7I[m��oa ������c/��$PARAM_M�ENU ? ��  �DEFPUL�SE
	WAI�TTMOUT�{�RCV� S�HELL_WRK�.$CUR_ST�YL�p"�OP9T8Q8�PTBM�G��C�R_DECSN�p�	������� ����-�(�:�L�u��p��������qSSR�EL_ID  ���̕USE_PROG %�zq%���͓CCR�p�ޒ��s1�_HOSoT !�z!6�s�+�T�=���V�h����˯*�_TIM�E�rޖF��pGD�EBUGܐ�{͓G�INP_FLMS�K��#�TR2�#�P+GAP� ��_b��CH1�"�TYPE
�|�P������ ��0�Y�T�f�xϡ� �Ϯ����������1� ,�>�P�y�t߆ߘ��� ������	���(�Q��L�^�p��%�WOR�D ?	�{
 �	PR�p#MsAI��q"SUd����TE��p#��	1���COLn%��!�Z��L�� !���F�d�TRACECTL 1� ��q ���#���_�DT �Q� ��z�Do � ��� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�U ��oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *� oN�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/Bϐ/�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX j|������ ���0�B�T�f�x�����������$PG�TRACELEN�  ��  �_����Ά�_UP ���������  ���΁_CFG M���烸�
���*�*�D�O���O��  �O��D�EFSPD ܲ������΀H�_CONFIG s���� �����dĔ�݂ ���ǑP^�a�㑹���΀IN�TRL' ��=�8^����PE��೗����*�ÑO�΀LI�D���	T�LL�B 1ⳙ k��BӐB4��O� 䘼����~Q� <<�  ?������ �M�3�U���i����� ����ӿ��	�7�T�Ϣk�b�tϡ�诚���������S�GRP� 1爬���@�A!���4I����A �Cu��C�OCjVF�/��Ȕa�z���ÑÐ�t��ޯ�s���´�ӿߨ�B �����������A��S�&�B34�`_������j�� ��������	�B�-����Q���M�������  Dz����.��� ��&L7p[� ������6�!Zh)w
V�7.10beta�1*�Ɛ@�*��@�) @�+�A Ē?���
?fff>�����B33A��Q�0�B(��A���AK��h ����//'/9/
P�p
�W�ӑ�n/��/�%���R�f?h����
�M +�?�/[��/�/�/�/�C?*��Ĕ�I�u �&:���?��x?�?A����P!\3 Bu�B���?�5BH�3[4b��o��4��[4R5��/B\3x3Dx�?@YO�?aOkO}O�<<� R@��O�C�O�O�O�O��DA�X�KNOW_�M  Z�%�X�SoV 賚ڒ ]��_�_�_?�_�_��_o����W�M+�鮳� ��	<�3#���_�o�\~=��
]bV4�@u��u��e�o�l��X�MR+��JmT�3?��W�1C{�OADBANFWDL_�V�ST+�1 1����P4C��� [��i/����� ?�1�C���g�y����� ���ӏ�*�	��`�?�Q�c��w2�|Va��up�<ʟ���p3 ��Ɵ؟Ꟃw4��+�=��w5Z�l�~�����w6����ѯ㯂w7  ��$�6��w8S�e�Xw����wMAmp�������OVLD � ��yo߄rP�ARNUM  ��{+þ�?υqSCH�� �
��X���{s��UPDX�)ź�|�Ϧ�_CMP_@`����p|P'yu�E�R_CHK����yqbb3��.�RS8pp?Q_MOm���_}ߥ�_RES_G�p쩻
�e��� ��0�#�T�G�x�k�}� �������������������������:� Y�^���Y�y������� �������������� ��R�6UZ�ӥ��u����V 1���FvpVa@k�p���THR_INR�p��(byudMA�SS Z)MN�GMON_QU?EUE �uyvTup\!��N�UZ�qNW��END��߶EXE�����BE���OPT�IO��ۚPROGRAM %z�%��~ϘTA�SK_I��.OCFG �z+�n/^� DATACc�+�1#s2ae?"? 4?F?X??|?�?�?�?��?o?�?�?OO�/IWNFOCc��-�� �?wO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_:GFD���, 	��!��K�_�!�)fN!fECNB��0m��Pf2Yo�khG�!2�0k �X,		d�=���·o���e�a$��pd��i�i�g_E?DIT ��/%�7����*SYS�TEM*upV9.�40107 cr7�/23/2021� A��Pw���PRGADJ_�p  h $X|[�p $Y�xZ�xW�xқtZқt?SPEED_�p�p�$NEXT_C�YCLE�p���q�FG�p ���pALGO_V� �pNYQ_F�REQ�WIN_�TYP�q)�SIuZ1�O�LAP�r�!�[��M+����qC?REATED�r��IFY�r@!NAM��p%h�_GJ�S�TATU��J�DE�BUG�rMAIL�TI����EVE<U��LAST������tELEM� �� $ENAB<�rN�EASI򁼁�AXIS�p$P�߄�����qROT�_RA" �rMAX� ��qE��LC�A�B
���C D_L9VՁ`�BAS��`��1�{���_� ��Y$x���RM� RB��;�DIS����X_cSPo�΁�� �u|�P� | 	�� 2 \�AN�� �;����8�Ӓ�� �0�PAYLO��3�V�_DOU�qS���p��tPREF� �( $GRID*�E
���R���9Y��rOTOƀ�q�  �p��!��p��k�OXY�� � $L��_�PO|�נVa�S�RV��)���DI?RECT_1� �U2(�3(�4(�5(��6(�7(�8��qFꔑA�� $V�ALu�GROU�P�������� !��@!��8�����RAN泲�⚁R��/���TOTaA��F��PW��I=!%�REGEN #�8�������/��фڶnTzЉ���#�_!S����8�(�V[�'�8��4���GRE��w����H��D�����V_]H��DAY3�V���S_Y�Œ;�SU�MMAR��2 �$CONFIG�_SEȃ���ʅ_�RUN�m�C�С�$�CMPR��P�D�EV���_�I��ZP�*��q��ENH�ANCE�	�
����1���INT���qM)b�q�2Kܖ���OVRo�PG�u�IX��;���OV�CT���  ��v�
 4 ����a˟���PSLG"�� \ �;��?��1���SƁϕc��U�����Ò�4�U��q]�Tp� Q(`�-��rJ<�O� =CK�IL_MJ���1VN�+��TQn{�iN5���C�ULȀjD�V(�C6�P_�ഺ�@�MW�V1V�VU1d�2s�2d�3s�3d�4s�4d��'��	�������p	�IN	VIB1qp1� �2!pq/,3 3
,4 4,�p?�� ;��A���N�����v��PL��TORr�3�	��[�SAVޒ�d�MC�_FOLD 	$SL������M,�I��L� �pL�b��KEEP�_HNADD	!xKe�UCCOMc��k��
�lOP���pl��lREM�k��΢����U��ekH�PW� KSB�M��ŠCOLLAAB|�Ӱn��n�+��IT�O��$N=OL�FCALX� ÇDON�rZ���7 ,��FL����$SYNy,M��C=����UP_�DLY�qs"DE�LA� ����Y(�A�D��$TABT�P_R�#��QSwKIPj% �䠆��OR� �E�� P_��� �)���p7 ��%9��%9A�$:N�$: [�$:h�$:u�$:��$:�9�q�RA��c X�����MB�NFLIC]��0"��U!�o���NO_H�� �\�< _SWI�TCHk�RA_P�ARAMG�� ��p��U��WJ���:Cӣ�NGRLT� OO�U�����X�<A��T_Ja1F�r�APS�WEIGH�]�J4CH�aDO1R��aD��OO��)�D2�_FJװ���sA�AV��C�HOB.�.�`��J2�0�q$�EeX��T$�'QIT���'Q�pG'Q-�G�pR�DC�m" � ��<��
R]��
H�<��RGEA��4��U�FLG`g��H���ER	�SPC�6R�rUM_'P��2�TH2No��@Q �1 XPED�����  D q�وIi�2_P�2�5cS�ᰁ+�L10_CI�WQd� �pk����U ՖD��zaxT�p�Q(�;a��c��޲+��i��e��` P>`DESIGRb$�VL1:i1Gf�c�g;10�_DS��D�~�cFPOS11�q l�pr��x1C�/#AT�B��U
WusIND��}�mq�Cp�mq`B	�HOMQE�r`!@s2GrM�_q����!@s3Gr��� ��$�+ >u4GrG�Y��k�}�������5Gr�ď֏������w6GrA�S�e�w�����
6�7Gr��П���(��6�8Gr;�M� _�q������uS �q    �@sM��P6��K@��! aT`M��M�IO���m�I��2�OK _O�Py��� �E��bPO{WE" 7��x EQ�1E � y#s%Ȳ$DSBo�GGNA�b� C�P�2�BS232S�$� �iP��xc�I3CE<@%�PE`2�� @IT��P�OPB�7 1�FLOW�T�Ra@2��U$�CU8N��`�AUXT��2�>��ERFAC3İ�UU���SCHN��% t<_9��EЎA$FREEOFROMЦ�A�P8X q�UPD"YbfA�PT.�pEEX04����!�FA%b��5��RV�aG� _&  C�E�"- 1�AL�  �+��jc'��D�  2&� �S\PcP(
O  �$7P�%�Rh�2SP��T�`AXU���DSP���@�W���:`$��RNP�%�@�����K��_MIR������MT��A�P���P"�qD�QSaYz������QPG7�BRKH���ƅ A;XI�  ^���i���1 ����BS�OC���N��DU�MMY16�1$�SV�DE��I�FSPD_OVR7�9� D����OR$��֠N"`��F_����@OV��SF�RUN��"F0����ӳUF"@G�TOd�L�CH�"�%RECOV��9@�@W�`&�Ӑ�H��:`_0� � @�RTINVE\��8AOFS��CK�KbFWD������X1B��TR�a�B �FD� ��1= B1pBL� �6� A1L�V��Kb����#0��@+<�AM:��00��j��_M@ ~�@h���T$X`x �>�T$HBK���F���A�����PPA�
��	�������DVC_DB �3@pA�A"��X1`�X3`��S�@�`�0��Uꣳ�h�CABPP
R�S #���c�B�@���GUB'CPU�"��S�P�` R��11)ARŲ~�!$HW_CGp l�11� F&A1Ԡ@~8p�$UNITr��l e ATTRI8r@y"��CYC5B��CA��FLTR_2_FI�������2bP��CHK_n��SCT��F_e'cF_o,�"�*FS�Jj"CHA�Q�'918Is�82RSD���0�1���_Tg�`�� i�EM�NPM"f�T&2 8p&2- ޫ6DIAGpERAOILACNTBMwУLO@�Q��7��P�S��� � ��P�RBSZ`�`BCt4&�	��FUN5s��RIN�PZaߠ�07Dh�RAH@���`� `C�@�`C�Q�?CBLCURuH�DaA�K�!�H�HDAp�0aA�H�C�ELD�������C��jA�1�CT�IBUu�8p$C�E_RIA�QJ�AF P��>S�`DU�T2�0C��};OyI0DF_LC�XH���k�LMLF�a�HRDYO���RG�@HZ0��ߠ�@�UMULSE�P�']3iB$J��J�����FAN_AL�M�dbWRNeHGARD��ƽ�P��Bk@2aN�r�J�_}�AUJ R+4�TO_SBR��~b����je 6?A�cMPINF��{!�d�A�c7REG�NV��ɣjZ�D��NFLW%6r$M�@� ��fd� �0 h'uCM43NF�!�ON	 e!�e#�(b*r3F�3 ��	 ���q)5�$��$Y�r����u�_��p*$ ��/�EG@����qAR��i���2�3�u�@�<�AXE��ROBn��RED��WR��2c�_���SY`��qt� ?�SI�WRI���vE STհ�ӭ d�J��Eg!���t8��D^a��B����9�3.� OTO�a����ARY��ǂ�1������FIE���$LwINK�QGTH�M�T_������s30���XYZ��8�!*�OFF���)��ˀB��,B�l������m�FI@� ��C@Iû�,B��_J$�F�����S`4����3-!$1�w0Ƚ��R��C��,�DU����3�P�3TURB`XS.�Ձ�bXX�� ݗFL�d���p�L�0���34���� W1)�K��M��5�5%B'��ORQ�6��fC㘴��0B�O;�D�,����ќ�a�OVE��rM �����s2��s2��r1����0���0�g /�AN =!�2�DQ�q���q� }R�*��6����s��LV���ER��jA	�2!E��.�C��A���0��XE�2Ӈ�A��AAX��F��A�N!� SŴ1_��Q_Ɇ�^ʬ� ^ʴ�^��0^ʙ�^ʷ�^�1&�^ƒP[ɒPk� �P{ɒP�ɒP�ɒP�� �P�ɒP�ɒP������x� �R>�DEBU=#$8ADc�2����
�CAB�7����V� <" 
��i�q�� -!��%��׆��׬��� �����1�י��׷�JTp��DR�m�LAB��qݥ9 FGRO� 4ݒ=l� B_�1� u���}��`����ޥ��qa��AND���� ���qa� �Eq���1��A@�� �NT8$`��c�VEL�1���m��1u���QP��m�NA[w�(�CN1� ���3줙�  �SE�RVEc�p+ $�@@d@��!��P�O
�� _�0T �!�󗱬p, w $TRQ�b�
(� -DR2�,+"P�0_ .� l"@!�&ERR���"I� q���~TOQ����L�p]�e���0G��%�����|	 �@ / ,��/I -��RA� �2. d�&��"  0�p$`&��2tPM��OC�A�8 1  pC�OUNT�� ���SFZN_C;FG2 4B �f�"T�:#��Ӝ��Z��`�s3 ���M:0�R�qC@��/�:0�FA1P��?V�X�����r����� �P:b�pHE�Lpe4 }5��B_BAS�c�RSR�f @�SH�!QY 1�Y 2|*U3|*4|*5|*6|*e7|*8�L!RO�����NL�q �AqB���0Z ACK��[INT_uUS`8�Pta9_PU�>b%ROU��PH@�h9#�u`w�9�TPFWD_KAR��ar RE���PP��A�QUE�i&��	�f�>`QaI`��9#�j38r��f�SEME��6t��PA�STY43SO�0�DI'1�`p���18�rQ_TM�c�MANRQXF�E�ND�$KEY?SWITCHj31�:A�4HE	�BEA�TM�3PE�pLEP����HU~3F�4�2S?DDO_HOeMBPO:a0EF���PRr��*�v�uC��@O�Qo �OV_�Mϒ��Eq�OCM����7� �8%HK��q5 D��g�U�j�2M�p�4R��FwORC�cWAR����P8%OM�p G6 @�Ԣ�v`U|�EP�p1�V'p�T3�VY4����S#O�0�L�R7��hUNLiOE0hdEDVa�  �S�@d8� <pAQ9�l1M�SUPG�UaCALC_PLANccM1��AYS1�1:b>�9 � X`��P �q;a�թ�w��2��j�M$P�㣒�fXyt$��rSC�M�p m�q ���aq��0�t5YzZzEU�Q�b�� T!�Hr�pPv�p��SNPX_AS�f: 0g ADD|��$SIZ%a�$VA��MU/LTIP�"ns�P�A�Q; � A$T9op�B���rS���j!C~ �vFRIF��2S�0�YT�pN=F[DODBUX�B�0�u&�!���CMtA��������������|Z ��< � �pƛTEg�����$SKGL��T��X�&{𷃥㰀��STMT<e�ЃPSEG�2���BW���SHOW�؅�1BAN�`TP�O���gᣥ�������, V�_G�= ��$PC���O�kFB�QP\�SP�01A&0^���VDG���>� �cA00�����P���P��P�P���P��5��6��U7��8��9��A�� b`���P��w᧖S`��!F����h���1��v�Th�י1�1�1��U1�1�1%�12�U1?�1L�1Y�1f�U2��2��2��2ʙU2י2�2�2��U2�2�2%�22�U2?�2L�2Y�2f�U3��3��3��3ʙ3י3�3���Ȫ�3�3%�32�3�߹3L�3Y�3f�4���4��4��4ʙ4�י4�4�4��4��4�4%�42�4�߹4L�4Y�4f�5���5��5��5ʙ5�י5�5�5��5��5�5%�52�5�߹5L�5Y�5f�6���6��6��6ʙ6�י6��6�6��6��6(�6%�62�6�߹6L�6Y�6f�7���7��7��7ʙ7�י7��7�7��7��7(�7%�72�7*߹7L�7Y�7f�OR�V�`_UPD��?s �c 
9`�V���@ x �$TOR�1T�  ��cOP �, ZQ_7RE^��� J���SsC�A��_�U�p� 7 YS�LOA"A �  �u$�v��w�@���@<��bVALUv10�6�F�ID_YL[C:HI5I�R?$FILE_X3e�u4$�C�SAVΔ�B hM �E_BLCK�3�ȁ�D_CPU��p� �p5hzQPY��R3�R C � �PW��� 	�!LAށSR�#.!'$RUN�`G@%$D!�'$�@G%e!$e!'%H`R03$� '$�QT2Pa�_LI�RD  ]� G_O�2�0�P_EDI�R�pTo2SPD�#E�"�i0ȁ�p	��D�CS9@G)F � 
$JPC71Tq�� S:C;C9�$MDL7$�5P>9TC�`@7UF�@?8S� ?8COBDu �@ �"|�L�G�PE;;� 9:;�OQTABUI_��!L�HGb�% �FB3G$�3A��sR�LLB_AV�AI�B?��3�!��I� $� SEL� N�Ẽ�@RG_D N���Ta���3SC�P�J �1/AB�PT��R�1w@_M]`L�Kc \M f/QL_�R�FMj��PGi�U9R��6��PS_�P�\� �p�EE7B�TwBC2�eL ����``�`b$�!FT��P'T�`
�TDC�g�� BPLp�sNU;WT�H��qhTgtWR��2$�pERVE�.S�T;S�Tw�R_A�CkP MX -$�Q�`.S�T;S�P�U@�`IC�`LOW&�GF1�QR2g�`��p�S�ERTI�A�d^0iP�PEkD�EUe�LACEM&zCC#c�V�BrppTf�edg�aTCV�l�adgTRQ�l�e�j@|�Scu��edcu�J7�_ 4
�J!��Se@qde�Q2�0���1��PRcuPJKlvVK@<�~qcQ~qw�spJ0�l�q�sJJ�sJJ�sAAL�s�p�s�p�vd���r5sS�`N1�l �p�k�`5dXA_́�IR_QCF�BN{ `M GROU (��bh�NPC0sD�?REQUIR�R� GEBU�C�Q�6g0 2Mz��Pd�Q�SGUO�@�)A�PPR0C7@� 
u$� N��CLO� �ǉS^U܉Se>@BC��@A�"P �$PM�]P�`�`sR�_MGa!�C���+��0�@�,�BRK*�NOL�D*�SHORTM!O�!m�Z��JWA�SP�tp`�sp`�sp`�s�p`�sp`�A��7��8�sQ�B�PTQ� m��R.Q�cQ�PATH�*� �*���X&���P�NT�|@A�"p��� �INF�RUC4`a��C�`KUM��Y
`�)p ��>�Q��cP���p���PAYLOAh�J;2L& R_Am@ꥁL �����+�R_F2LSHR�T/�LO���0���>���ACRL0z�p�y��ޤsRH5b$H�+���FLEX��:��JVR P��_�._�_�_QJ�US :�_�Vd`0ǀG��_tQd`�_�_lF1G��ũ�o0oBoTofoxo��E�o�o�o�o �o�o�o ����w z3lt����3EWF�^zT!��X�'qju ��uu~�W؁�� �p�u�u�u�u���t��RJ(�T �P`5�G�Y�� ' AT��l�pEL0�_B��s��J�Sz�JEW�CTR7B`NA��d�HAND_VB��Q��TUO@`4+�`TSW� �P�V� $$M��e G�AV�Qs�De�oAA���@�	$�A5�G�A�U�Ad�� 6��G�D*U�Dd�PD�G/ -CSTI�5V�5Ng�DYF ��+�x��� �P&�G�&�A��lw�o�Q�k�P������ʕ0ӕܕ��DX�T�W 7 �� ���3%�?!ASYM$T��m�T�V�o�A�t�_SH�~��� ���$����Ưد�J񬢐�#39"���_VI��`8�q0V_UNIrS�4��.�Jmu�2��2A��4 X��4�6a�pt��������&E_�������E���CH( Xc ̱���TOc�PP�VsSvD�US�RU�P�����z@�D�A}@_5�U��P�EyA�a��RPROG_N�A��$�$LAsST���CANs��ISz@XYZ_SP�u�DW]R@Ͱ,VS�V@�E1QENc��DC�UR�H�P��HR_�T��YtQ9S��d��O�T �9�tQ?�Z ��I�!A�D���Q���#��S����P3�vP �[ � MEB�O��R#B�!T�PPT0F@1�a��A̰� h1a%iT0�� $DUM�MY1��$PSm_��RF��  1��lfװFLA*�Y�P�bc$GLB_TI �U�e`ձ�PLIF(!\����g`OW�P��e�VOL#qb �a_	2��[d2�[`����b�P�cZ`TC���$BAUDv��cS�T��B�2g`ARI{TY0sD_WAIt�AIyCJ2�OU�6�ZqyyTLAN1S�`�{S�SZc��BUF_�r�fиx��PyyCHK_�@CkES��� JO`�E�aA�x�bUBYT�����r�.��.� ��aA��M���8����Q] Xʰ��֚�ST����SB=R@M21_@��T$SV_ER�bL����CL�`��A1��O�BpPGLh0EW~(!^ 4 $a�$Uq$�q$AW�9�A�@R��t%ՁUم_ "���D$GI��}=$ف ^҄��(!` L�.��"}�$F�"E6�NEA9R��B$F}�йTQ��J�@R� a�$J�OINTa�)� d�ӃMSET(!b E +�Ec�2�^�Se��PJ�_�(!c� � ��U�?���L?OCK_FO@� ޏPBGLV��GL6'�TE�@XM���'EMP��:�K��b��$U�؂a�2_���q�`<� �q�^��CE/�?���_ $KARb�M�STPDRA܀�����VECX�����IU�q�av�HE�TO�OL���V��RENǠIS3��6�ᦢACH̐m b^QOINe[d3���IdB��`@$RAIL_�BOXEa���R�OB�@D�?���HOWWAR0Aa�i`-�ROLMtb��$��*���T��`����O_�FU�!��HTML58QS�� e�"Հ�(!d��N@�@��(!e��������B�
8Ӄ}p(!f t��m��^a��t��B�POJ��AIPE�N����O����q��AORDED�m �z�XT`��A)��pPP��O�P g D �`OB���������Uc�`��� ��SYS��ADR��pP`|U@^  h ,"�N�f$A��EԼ�EnRVWVA�Qi � �@ق�U�PR�B�$ED�I�Ad�VSHWR2U�z���IS�Uq��pND�P7���G�H�EAD�! @���!fi�KEUqO`CP)P���JMP��L�UC��TRACE�TUj���IL�S��C��NE���T�ICK!MKQ��Q��HNr�k Q@���HWC��PHV�F��`STYeB+�LAO�a�S��[�C�l3��
�@�F%$A��D=:��S�!$�1�p� a�e�q�ePv HVS3QU��#LO�b_1�TERC`���T=S?�m 5���@R�m@3���ܡ�O`�	c IZ�d�A�e@ha�qtb}�hA}pP~rN��_DO�B�X�p9SSQ�SAXI�q��!v�bS�U�@TL��ƞREQ_ܠ��E�T���`�CY%��FdY'��Af\!\d�9x�P ЂSR$$nl-�w �@����c
�uV
Qh(�A���dC`�A��	�Y���D��p�E"�	CC�C��/�/�/	4�F�SSC�` o h5�DSmడ[`3SP�@�AT� 
R���L��XbADD�R�s$Hp� IF<�Ch�_2CH���pqO����- �TUk��Ir p��CU�CpnQV��I�Rq��4���c��
K�
p�^ ���Pr \z��D����|,K� P�"C�N��*CƮ��!�TXSCREE��qs�Pp@�INA˃<�4�D������`t Tᫀ�b�����O Y6���º�U4h�R�R�������R1�T����UE��u ��j �qz`Ś��RSML��U����V�1tPS_��6\��1�9G\���C��2@4� 2��0Ov�R��&F�AMTN_FL*�`Q��W� � �BBL_/�9WB`�Pw ����B5O ��BLE"�Cxg�R"�DRIGHt�RD��!CKGR�B`�ET���G�AWIDTHs���RB��a��r�UI��EYհRx d�ʰ�����`y�BACKЍ�tb>U���PFO܉�QWLAB�?(��PI��$UR�m�~P��P�PHy1 y 8 $�PCT_��,"�R�PRUp@�s5�da���QO%!Jt�zV�ȇ�pU�@r�SR ���LUM�S�� ERVJ�рP�P��T{ � " GE�Rh� �¯ГLPAeE��)�^g�lh�lh�ki5
ik6ik7ikpP`� Z�x����$u1��p��Q zQUS=Rل| <z��P1U2�a#2�FOO 2�PRI*m9�[�@p�TRIPK�m�oUNDO��})���Yp��y���Pi����p ~�Rp�qG ��T���-!&�rOS2��vR��2�s�CA�����rH`�F�h�UIaCA�����3Ib_�sOFFTA�D@���Ob��r�5�L�t��GU��Ps������+Q�SUB`� ��E/_EXE��Veуs�WO� �#���w��WAl�p΁zfP
 V_DB�H�9!pT�pO�V☖����3OR/�5�RAU@6�TK���y__���� |j ��OWNj�34$GSRC�0`���DA�<��_MPFI����ESP��T�$0��c��g�{n�z�E!G� `%�ۂ34J�n��COP��$`��p_���/�+�6���CT�Cہ�ہ���DCS��P�4�COMp�@�;��O`�=��b�K�^�/�VT�qU'���Y٤Z���2���@p�w#SB�����2�\0˰_��M8��%!]�DIC#��sAY�3G�PEE�@T�QS�VR1���eQL�� a��P�D  ��f�z��f�> ����6�QA�t�b# �~L2SHADOW���#ʱ_UNSCA�d�׳OWD�˰DG�DE#LEGAC�)�q'C�VC\ C>��� v����だm�RF07���7�d`C2`7�DRIVo���ϠC�A]�(��` ���MY_UBY�d?Ĳ��s��1�� $0�����_ఆ����L��BM�A$n�DEY	�EXp@,C�/�MU��X��,���0US����;p_R@"1�0p#�2�G�PACIN*���RG��c�y�:�y��sy�C/�RE�R"!�qq�y�D@� L 
!�G�P�"��Tp�	R�pD@�&P�Px1Q���	.���RE��SMWq�_Ar��+�{�Oq�AA/�3�h�EZ�U���� ��p�HK���P�J��_/�Q0{�EA�N��ۀ2�2�: �MwRCVCA� �:`GORG��Q�dR	��8L�����REFoG�� ���!�+`	�p��������<���q�_ ����r��� S�`C���Ú����@D� ���0�!��#q�š�O�U����?� ��Վ2�J@0� 1�*p����0 �UL�@��CO̷0)��� NT �[i�Z�Qf�af% L飏��Q���a�VIAچ�� �ÀHD7 6P�$JO�`oB��$Z_UPo��2Z_LOW��$�QxiBn��1$EP �s�y�� 1!f ���0æ4� 5��PA�A �C7ACH&�LO�w@�ВaB���Cn�%I#F^��Tm��N��$HO2�32{��Uÿ2O�@���R`o��=a��ƐVP��<X@A"_SIZ&�K$�Z$�F(�G'���CM]Pk*FAIo�G���AD�)/�MR1E���"P'GP�0����9�ASYNBUFǧRTD�%�$P!��COLE_2D_D4�5W�sw�~�U��QO��%ECCU��VEM��v]2�VIRC�!5�#�2��!_>�*&�pWp��AuG	9R�XYZ@�3�W���8��4+Q2z0T"��IM�16��2`�GRABB��q��;�LERD�C ;�F_D��F�f50MH�PE�R�0�������JRLAS��@��[_GEb�� �H൑~23�ET@����"���b��I�D��ҙ6m�BG_LEVnQ{�PK|Л6\q���GI�@N\P4� l��A��!g�dr�IS� �NRT��Lʁc�Ų��#a��c"!D�qDE����Xа(�X���0��2��
d��pzZ���d�c*���D4q�k�2puT��U&�� $�ITPr9p[Q��Փ�V�VSF$�d� a fp/�f�UR��5 R`MZu�dr���ADJ`C�� ZD�Vf� D�XAL�� � 4 PERI�KB$MSG_Q�3$Q!o% 
���p'��dr:g�q�Q� �XVR\t�̆B�pT_\��R��/ZABC"����Sr̚��
	�`�aAC�TVS' � �� $|u�0�cCgTIV�Q!IOu�s&D�IT�x�D�Vϐ
x�P��4�!���pPS����� �#��!���q!L�STD�!�  �_ST�tp�aq�;CHx�� L-�@���u�Ɛ*���P G�NA#�C�!q�_gFUN�� 	vp�IPu��HR�$�L���XZMPCF"��`bƀ�rX��ف��LNK��
C�Ł�0#�� �$ !��ބCMCM�k�C8�C"����P~{q $J8�2�D6!>�O�H�i�T��i�2�����M���UX�1݅UXE1Ѡ��1 C���Y���������˗7�FTFG>�������Z��� P�k�����YD'@_ � 8n�R� �Uӱ$HEIGHd�:h?(! 'v��z���� �c Gd��p$B% x� E��SHIF��hRVn�F�`�HpC� 3�(�8H`O� ѡ�C��+%D	�"��CE�pV���SP�HERs� � �,! M�c�u�	�$�POWERFL �4P|����|�p�RyG�`���������A� E ��?�p���pd���NSb ����?�  �Bz|� l�  <k@�|��%�涀�˃����ŵ�� �2ӷ�� 	H���l&���>ߪ��A |��t]$��*��/�� **:���p�ϥ�d�͘���������ɘ��|�����5� ������%ߟ�I�[� ��ߑ��������� ��w�!�3�a�W�i��� ���������O���� 9�/�A���e�w����� ��'����� =O}s���� ���k'UK ]������C/ ��-/#/5/�/Y/k/ �/�/�/?�/�/?�/ ?�?1?C?q?g?y?�? �?�?�?�?�?_O	OO�IO?OQO�� 	  �O�O�O_�E��3_����O`_�O�_�_÷PR�EF Ӻ�p��p
��IORITCY a|����p�����pSPL`z����WUqT�VqÈ�ODU~������_?�O�G��Gx��R��,fH�IBqOy�|kTO?ENT 1��yP?(!AF_t�`��o�g!tcp|�o}!ud�o~)~!icm��0bXY̳�k ;�|�)� �����p����u� �����N�5�r� Y�������̏�����	*/c̳ӹ���E��W�|�>�M#�FB��/��4���|��,��7�A��,  ��P����%�|�
'���Z��h�z������|��ENHA?NCE 	#�7��A9�d�����  �,f�T
�_�S��=��PORTe�rb��@�U��_C?ARTREP�Pr|>brSKSTAg�koSLGS�`�k�����@Unothing���� ��Ϳ>�P�b�To��TEMP ?i�sϨE/�_a_seibanm_��i_ �����0��T�?�x� cߜ߇ߙ��߽����� ��>�)�N�t�_�� ������������ :�%�^�I���m����� ������ ��$H 3lWi���� ���D/h S�w���uϪ��VERSI�P=g�  disa�ble��SAV�E ?j	2670H705�	�k/!�m//*��/ 	�(%b�O�+�/�Se?6?H?Z?l?�z:%<�/�?4�*'_�j` 1�kX ��0ubuE�?OqG�PURGE��Bp`�ncq�WF<@�a�TӒ*fW��`]Daa�WRUP�_DELAY �z�f�B_HOT %?e'b��OnE�R_NORMAL��HGb�O%_�GSEM�I_*_i_�QQSKKIP�3.��3x� �_��_�_�_�]?eo +goKo]ooo5o�o�o �o�o�o�o�o�o5 GYi�}�� �����1�C�U� �y�g���������я�����-�?�7%�$�RACFG ،[ќ�3�]�_P/ARAM�Q3y��Sw @И@`�G��42C۠��2���CbFB�B]�B�TIF���J]�CV�TMOU����]�]�DCR�3�Y� ��Q+��ۘBόB��e@��@?B�;��й_q��on�����;e�m����KZ;�=g�;�4�<<�૯f@�����  �5�G�Y�k�}��������ſ׿���xURD�IO_TYPE � �V�5��EDP�ROT_a�&�>��4BHbCE�ސSǆQ2c� ��B�ꐪϸ�� �ϐ����&�ݹ�W� V_~�o����߱��� ������A�O�m�r� ��9��������� �����=�_�d���� ������������� 'I�Nm��� ������#E Ji+k��� ���//4/F// g//�/y/�/�/�/�/ �/	?+/0?O/?c?Q? �?u?�?�?�?�?�??�;?,O��S�INT �2�I����1G;� jO|K��鯤O�f�0 �O�K�?�O �?___N_<_r_X_ �_�_�_�_�_�_�_�_ &ooJo8ono�ofo�o �o�o�o�o�o�o" F4j|b��� ������B�O��EFPOS1 1�"�  x O��o×O����ݏ� ����Ϗ0��T��x� ���7���ҟm����� ���>�P����7��� ����W��{����� :�կ^���������� S�e��� ��$Ͽ�H� �l��iϢ�=���a� �υ�� ߻����h� Sߌ�'߰�K���o��� 
��.���R���v�� #�5�o�������� ��<���9�r����1� ��U�����������8 #\����?� �u��"�FX �?���_� �/�	/B/�f// �/%/�/�/[/m/�/? �/,?�/P?�/t??q? �?E?�?i?�?�?O(O �?�?OpO[O�O/O�O SO�OwO�O_�O6_�O Z_�O~_�_+_=_w_�_ �_�_�_ o�_Do�_Aoxzocf�2 1r� o.oho�o�o
o. �oR�oO�#�G �k�����N� 9�r����1���U��� �������8�ӏ\��� 	��U�����ڟu��� ��"����X��|�� ��;�į_�q������ 	�B�ݯf����%��� ��[���ϣ�,�ǿ ٿ�%φ�qϪ�E��� i��ύ���(���L��� p�ߔ�/�A�Sߍ��� ����6���Z���W� ��+��O���s���� �����V�A�z���� 9���]��������� @��d��#]� ��}�*�' `���C�g y��&//J/�n/ 	/�/-/�/�/c/�/�/ ?�/4?�/�/�/-?�? y?�?M?�?q?�?�?�? 0O�?TO�?xOO�O�o�d3 1�oIO[O �O_�O7_=O[_�O_ _|_�_P_�_t_�_�_ !o�_�_�_o{ofo�o :o�o^o�o�o�o�o A�oe �$6H �����+��O� �L��� ���D�͏h� 񏌏�����K�6�o� 
���.���R���퟈� ���5�ПY����� R�����ׯr������ ���U��y����8� ��\�n�������?� ڿc�����"τϽ�X� ��|�ߠ�)������� "߃�nߧ�B���f��� ����%���I���m�� ��,�>�P������� ��3���W���T���(� ��L���p��������� ��S>w�6� Z����=� a� Z��� z/�'/�$/]/���//�/@/�/�O�D4 1�Ov/�/�/@? +?d?j/�?#?�?G?�? �?}?O�?*O�?NO�? �?OGO�O�O�OgO�O �O_�O_J_�On_	_ �_-_�_Q_c_u_�_o �_4o�_Xo�_|ooyo �oMo�oqo�o�o�o �o�oxc�7� [����>�� b����!�3�E���� ˏ���(�ÏL��I� �����A�ʟe�� �����H�3�l���� +���O���ꯅ���� 2�ͯV����O��� ��Կo�����Ϸ�� R��v�Ϛ�5Ͼ�Y� k�}Ϸ���<���`� �τ�߁ߺ�U���y� ��&��������� k��?���c������ "���F���j����)� ;�M���������0 ��T��Q�%�I��m��/�$5 1�/���mX� ��P�t�/� 3/�W/�{//(/:/ t/�/�/�/�/?�/A? �/>?w??�?6?�?Z? �?~?�?�?�?=O(OaO �?�O O�ODO�O�OzO _�O'_�OK_�O�O
_ D_�_�_�_d_�_�_o �_oGo�_koo�o*o �oNo`oro�o�o1 �oU�oyv�J �n������ �u�`���4���X�� |�ޏ���;�֏_��� ���0�B�|�ݟȟ� ��%���I��F��� ��>�ǯb�믆����� �E�0�i����(��� L���翂�Ϧ�/�ʿ S�� ��LϭϘ��� l��ϐ�ߴ��O��� s�ߗ�2߻�V�h�z� ��� �9���]��߁� �~��R���v����x#�	6 1& ��������������� }���<��`�� ��CUg� �&�J�n	k �?�c��/� ��	/j/U/�/)/�/ M/�/q/�/?�/0?�/ T?�/x??%?7?q?�? �?�?�?O�?>O�?;O tOO�O3O�OWO�O{O �O�O�O:_%_^_�O�_ _�_A_�_�_w_ o�_ $o�_Ho�_�_oAo�o �o�oao�o�o�o D�oh�'�K ]o�
��.��R� �v��s���G�Џk� 􏏏���ŏ׏�r� ]���1���U�ޟy�۟ ���8�ӟ\������ -�?�y�گů����"� ��F��C�|����;� Ŀ_�迃������B� -�f�ϊ�%Ϯ�Iϫ� ���ߣ�,���P�6�H�7 1S���� I��߲�������3� ��0�i���(��L� ��p�����/��S� ��w����6�����l� ������=������ 6���V�z � 9�]�� �@Rd���#/ �G/�k//h/�/</ �/`/�/�/?�/�/�/ ?g?R?�?&?�?J?�? n?�?	O�?-O�?QO�? uOO"O4OnO�O�O�O �O_�O;_�O8_q__ �_0_�_T_�_x_�_�_ �_7o"o[o�_oo�o >o�o�oto�o�o!�o E�o�o>��� ^�����A�� e� ���$���H�Z�l� ����+�ƏO��s� �p���D�͟h�񟌟 ���ԟ�o�Z��� .���R�ۯv�د����5�ЯY���}�c�u�8 1��*�<�v��� ߿��<�׿`���]� ��1Ϻ�U���y�ߝ� ������\�G߀�ߤ� ?���c����ߙ�"�� F���j���)�c��� ��������0���-� f����%���I���m� �����,P��t �3��i�� �:���3� �S�w /�� 6/�Z/�~//�/=/ O/a/�/�/�/ ?�/D? �/h??e?�?9?�?]? �?�?
O�?�?�?OdO OO�O#O�OGO�OkO�O _�O*_�ON_�Or__ _1_k_�_�_�_�_o �_8o�_5ono	o�o-o �oQo�ouo�o�o�o4 X�o|�;� �q����B�� ��;�������[�� �����>�ُb������!�������MAS�K 1 ��������ΗXNO  �ݟ���MOTE�  ���S�_CFOG !Z���N������PL_RAN�GV�N������OW_ER "��Ϡ���SM_DRYP�RG %���%�W��եTART �#Ǯ�UME_�PRO���q���_�EXEC_ENB�  ����GSP�DJ�������T3DB����RMп���IA_OPTIOYN��������NGVERS���`�řI_A�IRPUR�� pR�+���ÛMT_֐�T X���ΐOB�OT_ISOLC�����������N�AME8��H�ĚOB_CATEG��ϣ,��S�[�.�O�RD_NUM ?�Ǩ��H?705  N�����ߺ�ΐPC_TI�MEOUT�� x�ΐS232s�1$���� LT�EACH PEN�DAN��o���)���V�T�Ma�intenanc�e ConsN��&�M�"B�P�No Use6�r�8����������̒��NPQO$��Ҏ�"���/CH_LM�Q����	a�,�!UD�1:��.�RՐVA3ILw��粥*�_SR  t� ����5�R_INT7VAL���� ����V_DATA_GRP 2'����� D��P �������	��� ���B0R Tf������ /�/>/,/b/P/�/ t/�/�/�/�/�/?�/ (??L?:?p?^?�?�? �?�?�?�?�?O O"O $O6OlOZO�O~O�O�O �O�O�O_�O2_ _V_ D_z_h_�_�_�_�_�_ �_�_o
o@o.oPovo�do�o��$SAF�_DO_PULS�W�[�S���i�SCA�N�������SC�à(
�����
S�S�
������q�q�qN� �L^ p���5���� ��$��+�"�r2M�qX�dM�h�rJ�	t/� @��@������ʋ|��� r �ք��_ @N�T ��'�9�K�X�?T D��X��� ������ɟ۟���� #�5�G�Y�k�}�����x��䅎������Ǧ  "�;G�oR� ���p�"�
�u��D�i���q$q�  � ���uq%�\� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z����珈������ ������g�;�D�V� h�z���������������(�Ӣ0�r�i�y� ��$�7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/?r�+?=?O?a? s?�?�?�?�?�?8��? OO'O9OKO]OoO�O ��$�r�O�O�O�O 	__-_?_Q_c_u_�_ �Y�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4@FXj|�c�路 g�������0� B�T�f�x���������ҏ������:�.Ҧ��y�3�	��	123456�78��h!B!�� \��p0����Ο�� ���(�:�@��c� u���������ϯ�� ��)�;�M�_�q��� ��R���ɿۿ���� #�5�G�Y�k�}Ϗϡ� �����ϖ�����1� C�U�g�yߋߝ߯��� ������	��-���Q� c�u��������� ����)�;�M�_�q� ��B���������� %7I[m� �������! 3EWi{��� ����////� S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?D/�?�?�?�?�? OO'O9OKO]OoO�O@�O�O�O�O�O*��� �O	_�E�?5_G_Y_�yCz  A��z_   ��x2�r� }��)�
�W�  	�*�2�O�_�_ o$o"l�#\��_ho zo�o�o�o�o�o�o�o 
.@Rdv� ���Mo���� *�<�N�`�r������� ��̏ޏ����&�8��J��X #P$P�Q�R<�u� k��Q  ������S�P����Q�Qt  ЌPÙ۟�P(� `�,b����]�PFl��$SCR_GRP� 1*+�4� � ��,a �U	 v��~������d���%����ɯ���h]���P�D1� D�7n��3��Fl
C�RX-10iA/�L 234567W890�Pd� r���Pd�L ��,aC
1o��������[ ¶~�+fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@�R�d�t�?��H�~����m��ϴ����������,a��1���U�T[�G�imXhuP,��?B�  BƠߞ��Ԛ�A�P��  @�1`�՚�@����� ?���H��������F@ F�` A�I�@�m�X��|�� �������������`:�%�7�I�[�B�i� ��������������� -Q<u`��@En�ٯ���W�P�"+f@_�5��1`4b���x����ͣ�O�,dA����$���Fa�,a �#!"/4/E-!�Z(f/x/G/ (�P�!(� �/�/�/��/�/?#9b�����S7س�M�ECLV�L  ,a���ݲ�Q@f1L_D?EFAULTn4b1_�1`�3?HOTSTR�=���2MIPOWER�Fm0pU�5�4W7FDO�6 �5L��ERVENT 1�+u1u1�3 L!�DUM_EIP�#?5H�j!AF�_INE�0SO,d!'FT)O�NIO�O9!���O ��O�O�!RPC_MAIN�O�H��O>_S'VIS_�I�-_�_?!OPCUf�_�Wy_�_!TMP�PPU�_<Id�_�"o!
PMON_�PROXY#o?Fe ono�R<o8Mf]o�o�!RDM_SR�V�o<Ig�o!�R��"=Hh�oR!%
PM�o9LiA��!RLSYNC̟�y8��!gROS(O��4��6�!
CE�PMT'COM7�?Fk%���{!	K�CONS���>Glq�Ώ!K�WOASRC�o?Fm��v�!K�USB��=Hn	�f�!STM�0��;JoU����O�֟�c����CICE�_KL ?%K� (%SVCPGRG1��G�1�2G�DL�6�3o�t�6�4��D��6�5��į6�6��6�7��6���W�R�9_�d�3��� 6�9���6�a�ܿ6��� �6���,�6�ٯT�6� �|�6�)���6�Q��� 6�y���^����^�ʿ D�^��l�^�ϔ�^� Bϼ�^�j���^���� ^���4�^���\�^�
� �2���6��/� ���V��<�'�`�K� ��o����������� ��&J5nY� ������� 4F1jU�y� ����/�0// T/?/x/c/�/�/�/�/ �/�/�/??>?)?P?�t?_?�?
�_DEV� I�M{C:�84���4?GRP 2/E�0�+�bx 	�/ 
 ,@�?O ��ODO+OhOOOaO�O �O�O�O�O�O�O__ @_R_9_v_]_�_�_O �_�_�_o�_*ooNo `oGo�oko�o�o�o�o �o�o&8\�_ Q�I����� ��4�F�-�j�Q��� ����ď���Ϗ�� uB�T�;�x�_����� ��ҟ����ݟ�,�� P�7�t���m�����ί �7����(�:�!�^� E�����{�����ܿÿ տ���6��Z�l�S� ��篅���}������  ��D�+�h�z�aߞ� �����߻������� �R��v��o��� ��������*��N� `�G���k��������� ��k�8��\n U�y����� �	F-jQ� ������/ /B/T/;/x/_/�/�/ �/�/�/�/?�/,??�P?7?I?�?�3d ��6	t?�?�?�?�?O�?)O8K%�8O]O����vA"AvE�O �G~O�O�O�O�O�O
Y JO/_rI�O\_J_�_n_ �_�_�_�__o@_�_ 4o"oXoFo|ojo�o�_ o�oo�o�o0 TBx�o��oh� d���,��P�� w��@�����Ώ��ޏ ��(�j�O������ p�����ʟ��ڟ �B� '�f��Z�H�~�l��� ��Ư������د��  �V�D�z�h����ſ �������
��R� @�vϸ���ܿf��Ͼ� �������Nߐ�u� ��>ߨߖ��ߺ�����  �V�|�M��&��n� ��������.��R� ��F���V�|�j����� �����*���B 0Rxf���� ���>,N t���d��� �//:/|a/s/*/ L/&/�/�/�/�/�/? T/9?x/?l?Z?|?~? �?�?�?�?,?OP?�? DO2OhOVOxOzO�O�O O�O(O�O_
_@_._ d_R_t_�O�O�_ _�_ �_�_oo<o*o`o�_ �o�_Po�oLo�o�o�o 8zo_�o(� �������R 7�v �j�X���|��� ���*��N�؏B� 0�f�T���x�����՟ 矞������>�,�b� P���ȟ���v��ί ���:�(�^����� įN�����ܿʿ��  �6�x�]Ϝ�&ϐ�~� �Ϣ�������>�d�5� t��h�Vߌ�z߰ߞ� �����:���.���>� d�R��v������� �����*��:�`�N� �������t����� ��&6\����� L������" dI[4|� ����<!/`� T/B/d/f/x/�/�/�/ /�/8/�/,??P?>? `?b?t?�?�/�??�? O�?(OOLO:O\O�? �?�O�?�O�O�O _�O $__H_�Oo_�O8_�_ 4_�_�_�_�_�_ ob_ Go�_ozoho�o�o�o �o�o�o:o^o�oR @vd���� �6�*��N�<�r� `������Ϗ������ ��&��J�8�n����� ԏ^�ȟ��؟ڟ�"� �F���m���6����� į��ԯ֯��`�E� ���x�f��������� п&�L��\���P�>� t�bϘφϼ�����"� ��ߨ�&�L�:�p�^� ���ϻ��τ������  �"�H�6�l�ߓ��� \������������ D���k���4������� ������
L�1C�� ��d����� $	H�<*LN `����� � //8/&/H/J/\/�/ ��/��/�/�/?�/ 4?"?D?�/�/�?�/j? �?�?�?�?O�?0Or? WO�? O�OO�O�O�O �O�O_JO/_nO�Ob_ P_�_t_�_�_�_�_"_ oF_�_:o(o^oLo�o po�o�o�_�oo�o  6$ZH~�o� �n�j���2�  �V��}��F����� ��ԏ
���.�p�U� �����v��������� П�H�-�l���`�N� ��r��������4�� D�ޯ8�&�\�J���n� ���˿
�������� 4�"�X�F�|Ͼ���� l���������
�0�� Tߖ�{ߺ�D߮ߜ��� �������,�n�S�� ��t�������� 4��+������L��� p����������0��� $46H~l� ������  02Dz���j ����/
/,/� �y/�R/�/�/�/�/ �/�/?Z/??~/?r? ?�?�?�?�?�?�?2? OV?�?JO8OnO\O~O �O�O�O
O�O.O�O"_ _F_4_j_X_z_�_�O �__�_�_�_ooBo 0ofo�_�o�oVoxoRo �o�o�o>�oe �o.������ ��X=�|�p�^� �����������0�� T�ޏH�6�l�Z���~� ������,�Ɵ �� D�2�h�V���Ο��� |��x����
�@�.� d�����ʯT������ п���<�~�cϢ� ,ϖτϺϨ������� �V�;�z��n�\ߒ� �߶ߤ�������� ����4�j�X��|�� ����������� 0�f�T��������z� ������,b �����R���� �j�a�: ������ /B '/f�Z/�j/�/~/ �/�/�//�/>/�/2?  ?V?D?f?�?z?�?�/ �??�?
O�?.OORO @ObO�O�?�O�?xO�O �O_�O*__N_�Ou_ �_>_`_:_�_�_�_o��_&oh_Mo�_�Q�$�SERV_MAI�L  �U�`�~rhOUTPUT�h_�P@vd�RV 20f  �` (a\o�ovd�SAVE�l�iTO�P10 21�i d �_HZl ~������� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d�v������� ��П�����*�<��euYPscFZ�N_CFG 2e�c�T�a�e~|�GRP 23���q ,B   �AƠ�QD;� B}Ǡ�  B4�S�RB21�fH7ELL�4ev��`�o��/�>�%RSR>�?�Q���u� ����ҿ������,� �P�;�t�_ϘϪϼ�?�  �¼ϰ������� �P��&�'�ސW��2Pd��g��HKw 15�� ,� �߫ߥ��������� @�;�M�_���������������OMM� 6��?��FT?OV_ENB�d�a�u�OW_REG�_UI_�tbIMI_OFWDL*�7.��ɥ��WAIT\� `ٞ����`���d��wTIM�������VA�`����_UNcIT[�*yLCy�WTRY��uv`ME�8���aw�rdt ��9� ����h�<���X�Pڠ6p`?� � ��o+=1`VL�l�f�MON_ALIA�S ?e.��`heGo������ /)/;/M/�q/�/�/ �/�/d/�/�/??%? �/I?[?m??�?<?�? �?�?�?�?�?!O3OEO WOO{O�O�O�O�OnO �O�O__/_�OS_e_ w_�_�_F_�_�_�_�_ �_o+o=oOoaoo�o �o�o�o�oxo�o '9�o]o��> ������#�5� G�Y�k��������ŏ ׏������1�C�� g�y�����H���ӟ� ��	���-�?�Q�c�u�  �������ϯᯌ�� �)�;��L�q����� ��R�˿ݿ��Ͼ� 7�I�[�m��*ϣϵ� �����ϖ��!�3�E� ��i�{ߍߟ߱�\��� ��������A�S�e� w��4�������� ���+�=�O���s��� ������f����� '��K]o��> �����#5 GY}�����l�$SMON_�DEFPROG �&����� &*S?YSTEM*����RECALL �?}� ( �}/[/m//�/�/�/ I/�/�/�/?"?4? �/X?j?|?�?�?�?E? �?�?�?OO0O�?TO fOxO�O�O�OAO�O�O �O__,_�OP_b_t_ �_�_�_=_�_�_�_o o(o�_Lo^opo�o�o �o9o�o�o�o $ 6�oZl~��� G���� �2�� V�h�z�������C�ԏ ���
��.���R�d� v�������?�П��� ��*���N�`�r��� ����;�̯ޯ��� &���J�\�n������� ��I�ڿ����"�4� ǿX�j�|ώϠϲ�Eπ��������0���*�copy mc:�diocfgsv�.io md:=�>192.168�.56.1:17�447߆ߘߪ߽�5�K�frs:ord�erfil.da�t virt:\�temp\b�36�372���#�5� ;}-��*.d������ߊ�����
xy�zrate 11 V�h�z���/��������������������8����mpback��}�#5� }/K�dbS�*������������3x��:\T� f� �"4��4�a ��| ����� ��c~/!/3/F� j��/�/�/�Wi �??/?B�/�/x��?�?�?�tpdisc 0k?�0h?�z?OO/O�tpconn 0 �? �?�?�O�O�O@J�3SO eOwO__,_��Z/ ��_�_�_=/O/j_s/�oo(o7k�$SN�PX_ASG 2�:���Va�  0DQ�%�7o~o  ?��GfPARAM �;Ve`a �U	lkP>TDP>X~�d� ��I`�OFT_KB_CFG  CS\eFc�OPIN_SIMW  Vk�b+�=OYsI`RVNO�RDY_DO  ��eukrQST_P_DSB~�b|�>kSR <Vi � &�j�>W�>TW`I`TOP_?ON_ERRxGb~�PTN Ve�P��D:�RING_PRM'���rVCNT_GP� 2=Ve�ac`x 	���DP��я�����BgVD�RP 1>�i�`�Vq؏ 0�B�T�f�x������� ��ҟ�����,�>� e�b�t���������ί ���+�(�:�L�^� p���������ʿ��  ��$�6�H�Z�l�~� �Ϸϴ����������  �2�D�V�}�zߌߞ� ����������
��C� @�R�d�v����� ����	���*�<�N� `�r������������� ��&8J\n �������� "4[Xj|� ������!// 0/B/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?t?�?�?�?�?�?��?�?O�PRG_�COUNT�f�P�)IENBe�+EM�UC�dbO_UPD �1?�{T  
 ODR�O�O�O�O�O_ _A_<_N_`_�_�_�_ �_�_�_�_�_oo&o 8oao\ono�o�o�o�o �o�o�o�o94F X�|����� ����0�Y�T�f� x������������� �1�,�>�P�y�t��� ������Ο��	��� (�Q�L�^�p������� ���ܯ� �)�$�6� H�q�l�~�������ƿ ؿ���� �I�D�V��"L_INFO 1=@�E�@��	 yϽϨ������?=ք?����>G�q=�>�����´�� �Y�o�� D  ��  D	� �4  6(�l��~�-@YSDEBU)G:@�@�o�d�I��SP_PASS:E�B?��LOG �A���A  ro�i�v�  �A�o�UD1:\x��}���_MPC�ݐ�Ek�}�A&�� ��AK�SAV B���IAK��*�i��1�SVB�TEM_TIME 1C���@ 0o�zEzE�2�%���MEMBK'  �EA��x�����X|�@g� @��n���� ������h�9
�� K�@�as� �J߻���nà@Rdv� ����
Le�/ /(/:/L/^/p/�/�/ �/�/�/�/�/ ??$?06?H?Z?��SKV�[��EAj��?�?�?��=Bo�4]��Oo� � 
�
:O.@R�O��O�O}N�o�� ��OBi�p�O_'_9_-L2�Y_�_�_�_�_�_o�$�_�_� o'o9oKo]ooo�o�o �o�o�o�o�o�o#�5GYk_?T1SVGUNSPD!��'����p2MO�DE_LIM �D��Ҋt2�p�q�E�݉uABUI_?DCS H}5��!�0�G�n��D���|-�X�>���*���� 
��e��iđ��r�i������uEDIT I���xSCRN �J���rS�G �K�.�(�0߅SK_OPTION�и^����_DI��ENB  -�����BC2_GRP 2L�����&AMP�C�ʓ�|BCCF2/�N���� =��`�>�W�B�g� ��x�����կ����� ���S�>�w�b��� ������Ͽ����� =�(�a�Lυϗ�Ň�� ��������v��
�/� U�@�yߧ��`�iМ� �߰�����
���.�� >�@�R��v����� �������*��N�<� r�`������������� ��̀4FX�� |j������ �B0fTv x�����/� ,//</b/P/�/t/�/ �/�/�/�/�/�/(?? L?d?v?�?�?�?6? �?�?�?O O6OHOZO (O~OlO�O�O�O�O�O �O�O __D_2_h_V_ �_z_�_�_�_�_�_
o �_.oo>o@oRo�ovo �ob?�o�o�o�o <*Lr`��� �����&��6� 8�J���n�����ȏ�� �ڏ��"��F�4�j� X���|��������֟ ��o$�6�T�f�x��� ������ү������ �>�,�b�P���t��� �����ο��(�� L�:�\ς�pϦϔ��� �������� ��H�6� l�"��ߖߴ�����V� �����2� �V�h�z� H������������ ��
�@�.�d�R���v� ������������* N<^`r�� �����&8� \Jl����� ���"//F/4/V/ X/j/�/�/�/�/�/�/ ?�/?B?0?f?T?�? x?�?�?�?�?�?O�? ,O�DOVOtO�O�OO �O�O�O�O�O_ V4P��$TBCSG_�GRP 2O U��  ��4Q 
 ?�  __q_[_�__�_�_��_�_�_o%k8R?SQ~F\d�HTa�?4Q	 HA��}�#e>���>$a��\#eAT�̓A WR�o�hdjma�OG�?Lfg�bp�o�n�ffhf���ȼb4P|j��o*}@���Rhf�ff>�#33pa#e<qB�o+D=xrRp�qUy�rt~��H�y rIpTv�pBȺt~	xf	x (�;���f���N�`�Ю�ˏڋ����	�V3.00WR	�crxlڃ	*@��3R~t��HH�ư� \�.�]�  cC.�����8Q+J2?SRF]�����CFG T UePQ SPܚ��9r�1��1�W� e�	Pe���v�����ӯ ��������Q�<� u�`���������Ϳ� ޿��;�&�_�Jσ� nπϹϤ������� WRq@�0�B���u�`� �߫ߖ��ߺ������ )�;�M��q�\��� ����4Q _���O �� �J�8�n�\������� ����������4" XFhj|��� ���.TB xf��nO��� �//>/,/b/P/�/ t/�/�/�/�/�/�/�/ ?:?(?^?p?�?�?N? �?�?�?�?�?�? O6O $OZOHO~OlO�O�O�O �O�O�O�O __D_2_ T_V_h_�_�_�_�_�_ �_
o�_o@o�Xojo |o&o�o�o�o�o�o �o*N`r�B �������&� �6�\�J���n����� ȏ��؏ڏ�"��F� 4�j�X���|���ğ�� �֟���0��@�B� T���x�����ү䯎o ���̯ʯP�>�t�b� ������������� Կ&�L�:�p�^ϔϦ� ���τ������ �"� H�6�l�Zߐ�~ߴߢ� ���������2� �V� D�z�h�������� �����
�,�.�@�v� ������\������� <*`N�� ��x��� 8J\(��� �����/4/"/ X/F/|/j/�/�/�/�/ �/�/�/??B?0?f? T?v?�?�?�?�?�?�? OO��2ODO�� O�O tO�O�O�O�O�O_�O (_:_L_
__�_p_�_ �_�_�_�_ o�_$oo 4o6oHo~olo�o�o�o �o�o�o�o D2 hV�z���� �
��.��R�@�b� ��v���&OXO֏菒� ����N�<�r�`��� ����̟ޟ🮟�� $�&�8�n�������^� ȯ���گ��� �"� 4�j�X���|�����ֿ Ŀ����0��T�B� x�fψϊϜ������� ����>�P���h�z� ��6߼ߪ��������� �:�(�^�p���R��������� ���  9&�*� *�>��*��$TBJOP_GRP 2U����  ?���C*�i	V�]�Wd������X � *��� ��, � ����*� @&�?���	 �A���~��C�  DD������>v�>\�? ��aG�:��o��;ߴ�AT������A�@<��MX����>���\)?����8Q�����L���>�0 &�;iG.��Ap< � F�A�ff�v��� ):VMՂ.�� S>o*�@w��R�Cр	���������f�f�:�6/�?��33�B    ��/�������>):�S����� �/�/@��H@�%&/�/��=� �<#�
*��v�;7/�ڪ!?���4B�3?'?2	��2? hZ?D?R?�?�?�?F? �?�?�?�?OAOO�?�`OzOdOrO�O�O*�C�*���A��	V�3.00{�crxl��*P��%��%c5Z F�� JZH F6�� F^ F��� F�f F�� G� G�5 G<
 G^�] G� G����G�*�G��S G�; G���ERDu�\E[�� E� F�( F-� FU�` F}  F��N F� F��� Fͺ F��� F�V G�� Gz G?a 9ѷ�Q�L�HefJ4�o,b�*�0c1���OH�E�D_TCH XXd�+X2S�&�&�d$'X�o�o*�1�F�TESTPARS  ��cV��HRpABLE ;1Yd� N`*�H�����g$j�g�h��h)�1��g	�h
��h�hHu*��h��h�h%vRDI0n�GYk}��u	�O�#�-�?�Q�Hc�u�)rS�l� �z 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z���I���m� Fwͩ��ȏڏ쏘������x)r��NUoM  ��n���2� Ep�)r_CFG Z���I���@V�IMEB�F_TTqD��e�޶VER������޳R 1[8{ �8�o*�%�Q� ��د  9�K�]�o� �ϓϥϷ��������� �#�5�G�Y�k�}��� �߳����������� 1���E�W�i�{��� ������������/� A�S�e�w��������� ������+=OR�_���@��`�LIF \��	D`����DR�](FP
�!p�!p�� d� ��MI_�CHAN� � ~DBGLVL���fETHER�AD ?u���0`1�_}�R�OUT�!�j!���SNMA�SKY�j255.%S///A/S��`OOLOFS_�DIp�COR�QCTRL ]8{��1o�-T�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OL�/6O%OZOcPE_�DETAI7�*P�GL_CONFI�G c�������/cell/$�CID$/grp1^O�O�O�O
__|���G_Y_k_}_�_�_ 0_�_�_�_�_oo�_ CoUogoyo�o�o,o>o �o�o�o	-�oQ cu���:�� ���)���_�q� ��������׮}N�� ��%�7�I�a�KOq�P��M�����ʟܟ�  �G�$�6�H�Z�l�~� �����Ưد���� ��2�D�V�h�z���� ��¿Կ���
ϙ�.� @�R�d�vψϚ�)Ͼ� �������ߧ�<�N� `�r߄ߖ�%ߺ����� ����&��J�\�n� ����3��������� �"���F�X�j�|���������@�Us�er View ��I}}1234567890�����+=Ex �e����2��B����@��`r��3� Oas����x4>//'/9/K/]/�~/x5��/�/��/�/�/?p/2?x6 �/k?}?�?�?�?�?$?�?x7Z?O1OCOUO gOyO�?�Ox8O�O �O�O	__-_�ON_TR� lCamera���O�_�_ �_�_�_�_˂E�_o )o;n��Uogoyo�o�o�o�)  mV�	�_�o #5GY o}� ��o������F_�mV=�k�}��� ����ŏl����X� 1�C�U�g�y���2�D� �"�ן�����1� ؏U�g�y�ğ������ ӯ�����D��k��E� W�i�{�����F�ÿտ �2���/�A�S�e� �nUY9���������� ��	߰�-�?�Qߜ�u� �ߙ߽߫���v�D�I f��-�?�Q�c�u�� ����������� )�;���D��I����� ����������) t�M_q���N�`�93��0 B��Sx�1��@���//�J	oU0�U/g/y/�/�/�/ V�/�/�/�?-??? Q?c?u?/./tPv[? �?�?�?OO(O�/LO ^OpO�?�O�O�O�O�O �O�?oU�k�O:_L_^_ p_�_�_;O�_�_�_'_  oo$o6oHoZo_;% N��_�o�o�o�o�o  �_$6H�ol~� ���moe��]� $�6�H�Z�l����� ���؏���� �2� �e&�ɏ~������� Ɵ؟���� �k�D� V�h�z�����E�e�� 5����� �2�D�� h�z���ׯ��¿Կ�x��
ϱ�  �� 9�K�]�oρϓϥϷ����������    ��5�G�Y�k�}ߏ� �߳����������� 1�C�U�g�y���� ��������	��-�?� Q�c�u����������� ����);M_�q�  
��( � �-�( 	 ������� #35G}k����
� � Y�
//./��R/d/v/ �/�/�/����/�/�/ A/?0?B?T?f?x?�/ �?�?�??�?�?OO ,O>O�?bOtO�O�?�O �O�O�O�O_KO]O:_ L_^_�O�_�_�_�_�_ �_#_ oo$ok_HoZo lo~o�o�o�_�o�o�o 1o 2DVh�o �o���	��
� �.�@��d�v���� ����Џ���M�*� <�N���r��������� ̟�%���&�m�J� \�n��������ȯگ �3��"�4�F�X�j� ����������ֿ��� ��0�w���f�xϊ� ѿ�����������O� ,�>�Pߗ�t߆ߘߪ� ���������]�:�L�^�p����߻@� ������������ ��"frh�:\tpgl\r�obots\cr�x!�10ia_l.xml��D�V�h� z�������������������0BTf x�������� �,>Pbt� �������/ (/:/L/^/p/�/�/�/ �/�/�/��/?$?6? H?Z?l?~?�?�?�?�? �?�/�?O O2ODOVO hOzO�O�O�O�O�O�? �O
__._@_R_d_v_ �_�_�_�_�_�O�_o o*o<oNo`oro�o�o��o�o�o�n �6�� ���<< 	� ?��k!�o ;iOq��� ������%�S� 9�k���o�����я�����(�$TPG�L_OUTPUT� f������ �&�8�J� \�n���������ȟڟ ����"�4�F�X�j��|�������į�p��ր2345678901�����1� C�K����r������� ��̿d�п��&�8�J��}T�|ώϠϲ� ��\�n�����0�B� T���bߊߜ߮����� j�����,�>�P��� �߆��������x� ���(�:�L�^���l� ����������t��� $6HZlz� ������ 2 DVh ��� ����/./@/R/ d/v//�/�/�/�/�/��/�/ۂ $$��ί<7*?\?N?�? r?�?�?�?�?�?�?O O4O&OXOJO|OnO�O �O�O�O�O�O_�O0_"_T_}�an_�_�_�_�_�_�]@�_o	z ( 	 V_ Do2ohoVo�ozo�o�o �o�o�o
�o.R @vd����� ����(�*�<�r��`���ܦ�  <<I_ˏݏ��� ����:�L�֪��}� ��)���ş������� k��C�ݟ/�y���e� ������������-� ?��c�u�ӯ]����� W���Ϳ��)χ��� _�q��yϧρϓ��� ��M��%߿��[�5� Gߑߣ�߫���s��� �!���E�W��?�� ��9���������i� ��A�S���w���c�u� ���/�����= )s�����U ���'9�! o	[����� K�#/5/�Y/k/E/ w/�/�/�/�/�/�/ ?�/?U?g?�/�?�? 7?�?�?�?�?	OO���)WGL1.X�ML�_PM�$TP�OFF_LIM ����P����^FN_SVf@  ��TxJP_MOoN g��zD��P�P2ZISTRTCHK h���xFk_aBVTCO�MPAT�HQ|FVWVAR i�M�:X�D �O �R_�P�BbA_D�EFPROG �%�I%�PAU�LP�_WL_DIS�PLAYm@�N�RI�NST_MSK � �\ �ZIN�USER_�TLC�Kl�[QUICK�MEN:o�TSCR�EY`��Rtpsc�Tat`yi4xB�`_�iSTZxI�RACE_CFGW j�I:T�@�	[T
?��hHNL 2k�Z���aA[ gR-?Qcu����z�eITEM� 2l{ �%�$1234567�890 ��  =�<
�0�B�J�  !P�X�dP���[S ���"���X�
�|� ��W���r�֏����.� �0�B�\�f�����6� \�n�ҟ�������� >���"���.����� ίR����Ŀֿ:�� ^�p�9ϔ�Tϸ�xϊ� ��d���H��l� �>�Pߴ�\������� v� ������h�(�� �߰�4�L��ߦ��� ��@�R��v�6���Z� l���������*��� N��� ���������� ��X���J
 n���b�� ��"4F�/| </N/�Z/���// �/0/�/?f/?�/�/ e?�/�?�/�?�?�?,? �?P?b?t?�?�?DOjO |O�?�OOO(O�O�O ^O_0_�O<_�O�O�_ �O�__�_�_H_�_l_(~_Go�dS�bm�oLj��  �rLjq �a�o�Y
 �o��o�o�o{jUD1�:\|��^aR_�GRP 1n�{� 	 @�P Rd{N�r����~��p���q+�x�O�:�?�  j� |�f����������ҏ ����>�,�b�P���`t���������	e����\cSCB 2ohk U�R�d� v���������Я�Rl�UTORIAL �phk�o-�WgV_�CONFIG �qhm�a�o�o��<�O�UTPUT r<hi}�����ܿ � ��$�6�H�Z�l� ~ϐϢϴ�z�ɿ����  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������� �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/��/�/?? 0?B?T?f?x?�?�?�? �?�/�?�?OO,O>O PObOtO�O�O�O�O�? �O�O__(_:_L_^_ p_�_�_�_�_�_f�x� ǿoo,o>oPoboto �o�o�o�o�o�o�O (:L^p�� �����o ��$� 6�H�Z�l�~������� Ə؏��� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я�� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� ���������������X���# ��N�_r���� ���&8J ��n������ ��/"/4/F/X/i |/�/�/�/�/�/�/�/ ??0?B?T?e/x?�? �?�?�?�?�?�?OO ,O>OPOa?tO�O�O�O �O�O�O�O__(_:_ L_^_oO�_�_�_�_�_ �_�_ oo$o6oHoZo k_~o�o�o�o�o�o�o �o 2DVgoz �������
� �.�@�R�d�u���� ����Џ����*� <�N�`�q��������� ̟ޟ���&�8�J��\�k��$TX_S�CREEN 1s�% �}�k�����ӯ���	���Z��I�[�m� ������,�ٿ��� �!�3Ϫ�W�ο{ύ� �ϱ�����L���p�� /�A�S�e�w��� ߭� ���������~�+�� O�a�s���� ��� D�����'�9�K��� �������������R� ��v�#5GYk}�����$UALR�M_MSG ?����� �n�� �	:-^Qc ������ /��SEV  ��2&�ECFG �u����  }n�@�  Ab!�   B�n�
 /u����/�/�/�/ �/�/??%?7?I?W7~>!GRP 2vH+w 0n�	 /��?� I_BBL_NOTE wH*�T��l�u���w�T �2DE�FPRO� %� (%�Ow�	OBO -OfOQO�OuO�O�O�O��O�O_�O,_�<FK�EYDATA 1yx���0p W'n� U?�_�_�00_�_�_�U,(7_o n��_7oo[oBoo�o xo�o�o�o�o�o�o 3E,iP��� �������A�p^��Q�x������� ��ҏu�f�����1� C�U��y��������� ӟb���	��-�?�Q� c�򟇯������ϯ� p���)�;�M�_�� ��������˿ݿ�~� �%�7�I�[�m����� �ϵ�������z��!� 3�E�W�i�{�
ߟ߱� �������߈��/�A� S�e�w������� �������+�=�O�a� s���\����������� 
�'9K]o� �"����� �5GYk}� �����//� C/U/g/y/�/�/,/�/ �/�/�/	??�/??Q? c?u?�?�?�?:?�?�? �?OO)O�?MO_OqO �O�O�O6O�O�O�O_ _%_7_�O[_m__�_ �_�_D_�_�_�_o!o 3o�_Woio{o�o�o�o��o���k�������o}�o8J$v,6�{.�� �������/� �S�:�w���p����� я�ʏ��+��O� a�H���l�������ߟ ���'�9�Ho]�o� ��������ɯX���� �#�5�G�֯k�}��� ����ſT������ 1�C�U��yϋϝϯ� ����b���	��-�?� Q���u߇ߙ߽߫��� ��p���)�;�M�_� �߃��������l� ��%�7�I�[�m��� ������������z� !3EWi���� �����П/ ASew~��� ���/�+/=/O/ a/s/�//�/�/�/�/ �/?�/'?9?K?]?o? �?�?"?�?�?�?�?�? O�?5OGOYOkO}O�O O�O�O�O�O�O__ �OC_U_g_y_�_�_,_ �_�_�_�_	oo�_?o Qocouo�o�o�o:o�o �o�o)�oM_ q���6������%�7�9�}����b�@t���^�������,�� 돞����3�E�,�i� P�������ß����� ����A�S�:�w�^� ������ѯ����ܯ� +�
O�a�s������� �Ϳ߿���'�9� ȿ]�oρϓϥϷ�F� �������#�5���Y� k�}ߏߡ߳���T��� ����1�C���g�y� ������P�����	� �-�?�Q���u����� ������^���) ;M��q���� ��l%7I [������ h�/!/3/E/W/i/ @��/�/�/�/�/�/� ??/?A?S?e?w?? �?�?�?�?�?�?�?O +O=OOOaOsOO�O�O �O�O�O�O_�O'_9_ K_]_o_�__�_�_�_ �_�_�_�_#o5oGoYo ko}o�oo�o�o�o�o �o�o1CUgy ������	� ��?�Q�c�u����� (���Ϗ������ ;�M�_�q�������~ ����~ ���ҟ���Ο�*��,�[���f��� ����ٯ�������3� �W�i�P���t���ÿ ���ο��/�A�(� e�Lωϛ�z/������ ����(�=�O�a�s� �ߗߩ�8�������� �'��K�]�o��� ��4����������#� 5���Y�k�}������� B�������1�� Ugy����P ��	-?�c u����L�� //)/;/M/�q/�/ �/�/�/�/Z/�/?? %?7?I?�/m??�?�? �?�?�?���?O!O3O EOWO^?{O�O�O�O�O �O�OvO__/_A_S_ e_�O�_�_�_�_�_�_ r_oo+o=oOoaoso o�o�o�o�o�o�o�o '9K]o�o� �������#� 5�G�Y�k�}������ ŏ׏������1�C� U�g�y��������ӟ ���	���-�?�Q�c� u��������ϯ��h���0���0���B�T�f�>�����t�,��˿~� �ֿ�%��I�0�m� �fϣϊ��������� ��!�3��W�>�{�b� �߱ߘ��߼�����? /�A�S�e�w��� ������������=� O�a�s�����&����� ������9K] o���4��� �#�GYk} ��0����/ /1/�U/g/y/�/�/ �/>/�/�/�/	??-? �/Q?c?u?�?�?�?�? L?�?�?OO)O;O�? _OqO�O�O�O�OHO�O �O__%_7_I_ �m_ _�_�_�_�_�O�_�_ o!o3oEoWo�_{o�o �o�o�o�odo�o /AS�ow��� ���r��+�=� O�a����������͏ ߏn���'�9�K�]� o���������ɟ۟� |��#�5�G�Y�k��� ������ůׯ����� �1�C�U�g�y���� ����ӿ������-�@?�Q�c�uχ�^P����^P���������ͮ���
���, ��;���_�F߃ߕ�|� �ߠ����������7� I�0�m�T������ �������!��E�,� i�{�Z_���������� ���/ASew ������ �+=Oas� �����//� 9/K/]/o/�/�/"/�/ �/�/�/�/?�/5?G? Y?k?}?�?�?0?�?�? �?�?OO�?COUOgO yO�O�O,O�O�O�O�O 	__-_�OQ_c_u_�_ �_�_:_�_�_�_oo )o�_Mo_oqo�o�o�o �o���o�o%7 >o[m���� V���!�3�E�� i�{�������ÏR�� ����/�A�S��w� ��������џ`���� �+�=�O�ޟs����� ����ͯ߯n���'� 9�K�]�쯁������� ɿۿj����#�5�G� Y�k����ϡϳ����� ��x���1�C�U�g� �ϋߝ߯�����������`����`���"�4�F��h�z�T�,f���^���� �����)��M�_�F� ��j����������� ��7[B� x�����o! 3EWixߍ�� �����///A/ S/e/w//�/�/�/�/ �/�/�/?+?=?O?a? s?�??�?�?�?�?�? O�?'O9OKO]OoO�O O�O�O�O�O�O�O_ �O5_G_Y_k_}_�__ �_�_�_�_�_o�_1o CoUogoyo�o�o,o�o �o�o�o	�o?Q cu��(��� ���)� M�_�q� �������ˏݏ�� �%�7�Ə[�m���� ����D�ٟ����!� 3�W�i�{������� ïR������/�A� Яe�w���������N� �����+�=�O�޿ sυϗϩϻ���\��� ��'�9�K���o߁� �ߥ߷�����j���� #�5�G�Y���}��� ������f�����1��C�U�g�>�i��>>�������� ����������,� �?&cu\�� �����) M4q�j��� ��/�%//I/[/ :�/�/�/�/�/�/�� �/?!?3?E?W?i?�/ �?�?�?�?�?�?v?O O/OAOSOeO�?�O�O �O�O�O�O�O�O_+_ =_O_a_s__�_�_�_ �_�_�_�_o'o9oKo ]ooo�oo�o�o�o�o �o�o�o#5GYk }������ ��1�C�U�g�y��� �����ӏ���	��� -�?�Q�c�u�����p/ ��ϟ�����;� M�_�q�������6�˯ ݯ���%���I�[� m������2�ǿٿ� ���!�3�¿W�i�{� �ϟϱ�@�������� �/߾�S�e�w߉ߛ� �߿�N�������+� =���a�s����� J�������'�9�K� ��o�����������X� ����#5G��k�}���������������&�HZ4,F/�>/���� �	/�-/?/&/c/J/ �/�/�/�/�/�/�/�/ ?�/;?"?_?q?X?�? |?�?�?���?OO%O 7OIOXmOO�O�O�O �O�OhO�O_!_3_E_ W_�O{_�_�_�_�_�_ d_�_oo/oAoSoeo �_�o�o�o�o�o�oro +=Oa�o� �������� '�9�K�]�o������ ��ɏۏ�|��#�5� G�Y�k�}������ş ן������1�C�U� g�y��������ӯ� ��	��?-�?�Q�c�u� ��������Ͽ��� Ϧ�;�M�_�qσϕ� $Ϲ��������ߢ� 7�I�[�m�ߑߣ�2� ���������!��E� W�i�{���.����� ������/���S�e� w�������<������� +��Oas� ���J�� '9�]o��� �F���/#/5/�G/�$UI_IN�USER  ����h!��  H/L/_�MENHIST �1yh% � ( u ���)/SOFTP�ART/GENL�INK?curr�ent=menu�page,1133,1�/�/??�	(�/�/5�/{?�?�?�?���?�?�?�?O "O4O�?XOjO|O�O�O �OAO�O�O�O__0_ �OA_f_x_�_�_�_�_ O_�_�_oo,o>o�_�boto�o�o�o�o�m� \a�!\o�o/A SVow����� `���+�=�O�� ���������͏ߏn� ��'�9�K�]�쏁� ������ɟ۟j�|�� #�5�G�Y�k������� ��ůׯ��o�o�1� C�U�g�y�|������� ӿ������-�?�Q� c�uχ�ϫϽ����� ��ߔ�)�;�M�_�q� ��ߧ߹�������� ��7�I�[�m���  ������������� �E�W�i�{������� ����������A Sew���<� ��+�Oa s���8��� //'/9/�]/o/�/ �/�/�/F/�/�/�/? #?5? �2�k?}?�?�? �?�?�/�?�?OO1O CO�?�?yO�O�O�O�O �ObO�O	__-_?_Q_ �Ou_�_�_�_�_�_^_ p_oo)o;oMo_o�_ �o�o�o�o�o�olo�%7I[F?���$UI_PANE�DATA 1{�����q�  	�}  �ttp://12�7.0�p1:30�80/frh/j�cgtp/fle�xdev.stm�?_width=�0m���  )�  rim�9�  �pP�b�t������� �����Ǐ��(�:� !�^�E�����{������ܟ�՟�I6� X14�G�L�^�p��� ������ʯ=�ܯ �� $�6�H�Z���~�e��� ����ؿ����� �2� �V�=�zό�sϰ�#��Ɠs�����)� ;�Mߠ�q�䯕ߧ߹� ������V��%��I� 0�m��f������ ������!��E�W��� �ύ�����������:� ~�/ASew� �����  =$asZ�~ ����d�v�'/9/ K/]/o/�/��/�/* �/�/�/?#?5?�/Y? @?}?�?v?�?�?�?�? �?O�?1OCO*OgONO �O�/�/�O�O�O	_ _-_�OQ_�/u_�_�_ �_�_�_6_�_o�_)o oMo_oFo�ojo�o�o �o�o�o�o%7�O �Om���� �^_�!�3�E�W�i� {������Ï����� ����A�S�:�w�^� ������џDV�� +�=�O�a�������
� ��ͯ߯���|�9�  �]�o�V���z���ɿ ���Կ�#�
�G�.�k�ޟ�}�|ϵ����������)��4ߧ� #�`�r߄ߖߨߺ�!� ���������8��\� C���y������������������$U�I_POSTYP�E  ��?� 	 �s��B�QUICKME/N  Q�`�v��D�RESTORE� 1|��?  ����!��������mA Sew�,��� ���+=Oa n����� //�9/K/]/o/�/ �/6/�/�/�/�/�/� ??0?�/k?}?�?�? �?V?�?�?�?OO�? COUOgOyO�O6?@O�O �O.O�O	__-_?_Q_ �Ou_�_�_�_�_`_�_ �_oo)o�O6oHoZo �_�o�o�o�o�o�o %7I[�o������SCRE���?��uw1sc��u2�U3�4�5�6��7�8��sTAT�M�� ����:�UGSER�p��rT�p��ks���4��5*��6��7��8��B��NDO_CFG �}Q�����B�PD�E���N�one��v�_IN_FO 2~��)���0%�D���2� s�V�������͟ߟ ��'�9��]�o�R����z��OFFSEOT �Q�-��� hs��p�����G� >�P�}�t���Я��׿ ο����C�:�L�@^Ϩ����͘���
�����av��WORK �!�����.��@ߢ�u�UFRAM�E  ���R�TOL_ABRT8�����ENB�ߣ�?GRP 1�����Cz  A�� ����*�<�N�`�r��֐�U�����?MSK  �)����N��%!��%xz����_EVN��b���+�ׂ3�«�
 h�UE�V��!td:\�event_usger\�u�C7z�d��jpF��n�SPs��x�spotwe{ld��!C6��������!���G |'��5kY�� ���>�� �1�Ug��� /��	/^/M/�/-/ ?/�/c/�/�/�/�/$?��/H?�/:J�W�3�����8C?�?�? �?�?�?�?O+OO OOaO<O�O�OrO�O�O �O�O_�O'_9__]_�o_J_�_�_�_�$V�ALD_CPC {2�« �_�_� w��qd�@R�*o_oqo��hsNbd�j�`��i�da{�o av�_�ooo3BoW i{�o�o�o�o��o �PA�0�e�w� �������� �(�=�L�a�s�
��� ����ʏ�����$� ޟH�:�o��������� ڟ؟����� �2�G� V�k�}�������¯ԯ �����.��R�S� yϋϚ���������� 	��*�<�Q�`�u߇� �ϨϺ��������� &�8�M�\�q���� ����n������"�4� F�[�j��������� �������!0�B�W f�{���������� �,>teT ������� /+/:La/p�/�/ ./�����//'? 6/H/?l/^?�?�?�/ �/�/�/�/?#O�?D? V?kOz?�O�O�?�?�? �?�?_O1_@ORO9_ vOw_�_�_�O�O�O_ �__-o<_N_`_uo�_ �o�o�_�_�_�_o &o;Jo\oq�o�� ��o�o�o� �"7� FXj������� ����!�0�E�T� f�{�������ßҏ� ���
�,�A�P�b��� ��x�����Ο���� �(�*�O�^�p����� ����R�ܯ� ��Ϳ 6�K�Z�l�&ϐ��Ϸ� ��ؿ���"� �2�G� ��h�zϏߞϳ����� ����
��1�@�U�d� v�]�ߛ��������� �,��<�Q�`�r�� ������������� &�;J�_n������ ��������$ F[j|���� ���0E/T i/x��/��/�/�/ �//,/.?P/e?t/ �/�/�?�?�?�?�/? ?(?:?L?NOsO�?�? �O�?�O�OvO OO$O 6O�OZOo_~O�OJ_�O �_�_�_�O_ _F_D_�V[�$VARS_�CONFIG ��Pxa�  FP]S��\lCMR_GRPw 2�xk h�a	`�`  %�1: SC130EF2 *�o�`]TəVU�P�h`�5�_Pa?�  A�@%pp*`�Vn 	No9xCVXdv��a��<uA�%p�q�_R��_R B���#� _Q'��H��l�;��� {�����؏ÏՏ�e� �D�/�A�z�-������ddIA_WORKW �xeܐ�Pf,		�Qxe��>�G�P ���Y�ǑRTSYNCS_ET  xi�xa�-�WINURL 3?=�`������������ȯگSI?ONTMOU9�]S�d� ��_C�FG �S۳�S۵P�`� FR:\��\�DATA\� ��� MC3�L�OG@�   U�D13�EXd�_Q'� B@ ����x�e_ſx�ɿ��VW � n?6  ���VV���l�q  =�C��?�]T<�y�Y�TRAIN���N� 
gp?�CȞ���TK���b�xk (g�����_����� ����U�C�y�g߁���ߝ߯������_GuE��xk�`_P��
�P�RꋰRE���xe*�`hLEXr�xl`1-e��VMPHASE � xec�ecR�TD_FILTE�R 2�xk �u�0����0�B� T�f�x�����VW���� ���� $6HZ�l_iSHIFTM�ENU 1�xk
 <�\%����������= &sJ\��������'/�	�LIVE/SNA��c%vsfli�v��9/��� �7�U�`\"menu r/w//�/�/����Y�]��MO��y�Y�5`h`ZD4�V��_Q<��0��$WA�ITDINEND���a2p6OK  !�i�<���?S�?�9wTIM�����<Gw?M�?*K�?
J�?x
J�?�8RELE���:G6p3���r1_ACCTO 9Hܑ�8_<�7 �ԙ�%�/:_<af�BRDIS�`�N��$XVR���y��$ZABCv�b1�S; ,��
j�I�2B_ZmI1�@VSPT �y�\�eG�
�*�/�o�*!o7o�WDCS?CHG �ԛ(���P\g@�PIPL2�S?i��o�o��o�ZMPCF_G' 1��ii�0'¯S�;Ms�S��i��p�'��g��e2޸�  ?�Gó;�.I��� D�  ��p	�r1��p�۞�� ���
�Z�~��N��Ï�>��4  6(�֏�ӈ*�� �*�@�N�x������*���D/@�1+�0 ��ן�Tp���o�_CYLIND��ݢ { Х� ,(  *=�N�G�`:�w�^����� ȟ ѯ���7����<�#� 5�r�����������޿ y�_����8�ύ�n�Ȁ�㜻ã wQ �5�����Sǟ��Ϡ(�ٻ�X�זr�A���SPHERE 2���ҿ��"� �������P�c�>�P� ̿t���ߪ����� '���]�o�L���p� W�i������������PZZ�F �6