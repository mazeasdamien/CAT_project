��   ��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����CCSCB_�GRP_T  � � $COM�PMATEXP � 9RIX �  0$IN7NER��P0D_�OFFSETS�hCMPAzCO}FsFS_TYCSBFRAMES � Y IT_T�OL�RANGE_� �r�FTRATIOS�h_H_LIM�D �L�FSOOFST1�
2�����$$CL�ASS  �S��3����(VERSION0o<XKD?IRTUAL0B�' 3 Q� �<  0 -��S��� ���  a����&�H��ٸ����� ���/��� ��B�,��4 @�=  ��D �W!o%k!C�  T%3 1 �� BpI'Z/�/�-