��   �c�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����DCSS_C�PC_T 4 �$COMMEN�T $EN�ABLE  �$MODJGRP�_NUMKL\�  $UFR�M\] _VTX �M �   $�Y�Z1K $Z�2�STOP_T�YPKDSBIO�IDXKENBL_CALMD��USE_PRED�IC? �ELAY�_TIMJSPEED_CTRLKOVR_LIM? *p D� �L�0�UT�OOi��O���&S. ǰ 8J\TC �u
!���\�� jY0 � � �CHG�_SIZ�$A�P!�E�DIS"�]$!�C_+{#�s%O#J�p 	]$J d#� �&s"�"{#�)�$��'�_SEEX�PAN#N�iG�STAT/ D�FP_BASE_ $0K$4�!� .6_V7>H�73hJ- � q}�\AXS\3UP�LW�7������d4r �< w?�?�?��?�?��// *%EL�EM/ T �&B.2NO�G]@%C�NHA�DF#� $/DATA)�6e�0  PJ�@ _2 
&P5' �� 1U*n   _VSiSZbR�j0jR(�VyT(�R|%S{TROBOT�X��SARo�U�V$�CUR_��R DS�ETU4"	 �$d P_MGN��INP_ASS e#�PB!� `CiH�7�7`e�.fXc1�C�ONFIG_CH�K`E_PO* }dS/HRST�gM^#/e�OTHERRBTF�j_G]�R�dTv ��ku�dVALD_�7h�e�4�FT1r
�0R HLHt� 0  �lt<NerRFYhH~t�5�1� ��9W�_A$R�JTwSPH/ (@G%Q�Q�Q3?wwBOX/ 8�@ F!�F!�G �r��s� DTUIRi@ � ,�F�pER�%@2 $�p �l�_Sf��uUIZN/ '0 IF(@�p&��Z_�0�_�0?wu0  @�QWyv	�*��~
�$$C�L`  ����!���Q��Q�V�ERSION��  XK~2�IRTUAL��0�' 2 ?�Q  (������&@^����P�����ϟ��������d<�9�Cz   P�8���a��������� ׯ�����.�@� R�d�f����������� �Կ	��*�<�N�`� r����ϫϺ�̿��� �߮�8�J�\�n�)� �ϧ߶��ς������ %�4�F�X�~�|ߎߣ� .����������!�0� B�T�f�x������� �������/>�P� b���v��������� �+:L^p �������  /'/9/HZl/�/ ��/����//#? 5?D/V/h/z/�/�?�/ �?�/�/�?
?O1OCO R?d?v?�?�O�?�O�? �?O	_�O-_?_NO`O rO�O�O�O�_�_�O�O o_)o;o�_\_n_�_ �_Mo�_�o�_�_�oo 7IXojo|o�o�o �o�R�o�o�3� E�Tfx����� Տ��ݏ��A�S� b�t���������џ�� ���(�=�O�^�p� ��������ʟ߯� � �$�9�K�]�l�~��� 6���Ưۿ����#� 2�G�Y�h�z������� ��Կ����
��.�C� U�g�vψϚϬϮ��� �����<�-��Q�c� r߄ߖߨߺ������� ��)�8�M�_���� ����q�������� ��4�&[m|����� �������v3 BWix���� ���/>?/ e/w/�����/� �///(/=?L/a?s? �/�/�/�/�/�?�/O ?$?9OH?]OoO�O�? �?�?ZO�O�?�OO O 2OG_VOk_}_�O�O�O �O�O�_�Oo_._Co R_goyo�o�_�_�_�_ �o�_	o*o`oQ@ u��o�o�o�o�o�o ��&8M�\q��� ��������� "�4��X�J������ಏď�����$D�CSS_CSC �25��?Q  P�;� ��Z���~�A�����w� د������ ��D�V� �z�=���a�¿��� �����߿@��d�'� ��KϬϾρ��ϥ�� ��*���N��r߄�G� ��k��ߏ��߳��&� ��J��n�1��U���y�������GR�P 2� ����	�s�^����� ����������'�� 7]H�l��� ����5 2 kV�z���� ��/
///U/@/y/ d/�/�/�/�/�/�/	? �/-??*?c?N?�?r? �?�?�?�?�?�?OO 'OMO8OqO\O�O�O�O �O�O�O_�O%__"_ [_F__�_�_n_�_�_ �_�_o�_oEo0oio��_GSTAT �2�E��<� 6�? �����5=��k�A����)�d�a5��M�� �D58o�G?�NC˃V�X`�<�f}m�>��%��>�4���$?�  �a��`4��Z����e�>t��=�H�?xj!�u���u)>wl��yC)��A� �VD,=� ziI��=>�?y ����9�`�����t�v���ܠ>k��P�&tg3=6�k�?y.�p��p���q>���}N��<Cz�D,���B��D,�9 y?|q�>��=�.�����?�p�Cy����`���z�`��D1��`yD���z�o�o�l�� \�n��P�������Џ ����jp������z !�O�5�G�i�k�}��� ͟��՟������ ŏ{�������ï���� ����O�5�c�-�k� Q�c����������Ͽ ����9�g�i�� ��ۯ���������'� �/�]��Eߓߥ�?� ���ߵ��������G� Y�3�}��i�{���� �������1�C��/� y�o߁߯���[����� ����-?cuO ������� )5_9K�� ����w�/%/� I/[/5/c/�/k/}/�/ �/�/�/?�/?E?? 1?{?�?g?�?�?�?�? �?��?/OAO�?eOwO QOcO�O�O�O�O�O�O _+___a_;_M_�_ �_�_�_�_�_�_oO OKo]o�_io�omoo �o�o�o�o�oG !3}�i��� ����1�C�9oG� y��e���������� я��-���c�u�O� ��������៻�͟� )��M�_�9�g���O� }�˯ݯw������ I�#�5����k���ǿ ������׿�3�E�� i�{�U�gϱϧ����� �ϓ��/�	��e�w� Qߛ߭߇߹��߽��� �+��O�a�;�m�� q������������� �K�]�7�����m��� ����������5G !O}Wi��� ���1��g y������ �/-//Q/c/=/O/ �/s/�/�/�/�/?? �/?M?CU�?�?/? �?�?�?�?OO�?7O IO#OUOOYOkO�O�O �O�O�O�O	_3___ i_{_q?_�_K_�_�_ �_�_o/o	o7oeo?o Qo�o�o�o�o�o�o�o �oOa;�� q���_���� 9�K�%�7���[�m��� ɏ�����ُ�5�� !�k�}�W��������� ����1�˟=�g� A�S�������ӯ寿� �����Q�c�=��� ��s���Ͽ������ ��M��9σϕ�o� ���ϥ��������7� I�#�m��Y߇ߵߏ� ��������!�3��;� i�#�Q���K����� �������	�S�e�?� ����u��������� ��=O);�{� ���g��� 9K%o�[�� �����#/5// A/k/E/W/�/�/��/ �/�/�/?1??U?g? A?o?�?w?�?�?�?�? 	OO�?#OQO+O=O�O �OsO�O�O�O�O_�/ �O;_M_�Oq_�_]_o_ �_�_�_�_o�_%o7o o#omoGoYo�o�o�o �o�o�o�o!_)_W iu�y��� ����)�S�-�?� ����u���я��ݏ� ��=�O�ES���� q���͟����ݟ� 9��%�o���[����� �����ǯٯ#�5���Y�k�a��$DCS�S_JPC 2�`�Q (G DQ�����ʴ Կذ����ʿܿ1� � �$�y�Hχ�l��ϐ� �ϴ�	�����,�Q� � 2߇�V�h�z��ߞ��� �����;�
�_�.�@� ��d�v��������� %���I��m�<�N��� ��������������3 W&{J�n� ������A O4�X�|�� ��/��O//0/ B/�/f/�/�/�/�/? �/'?�/?]?,?>?P? �?t?�?�?�?�?O�? 5OOOXO}OLO^O�O �O�O�O�O�O_�OC_ _g_6_�_Z_l_�_�_��_�_	o�_o4c��S
����Louo&o�o�`ddo�o�o�o�o	 �o-�oQu<� `r������ ;��_�&���J���n� ˏ��ُ���ڏ��� �m�4���X���|�ٟ ����ğ!��E��� 0�y���f�ï��篮� �ү/���S��w�>� ��b������������ �=��a�(υ�Lϩ� p��ϔ��ϸ�����%� K��o�6ߓ�Z߷�~� �ߢ�����#���1�� k�2�D�V�h������ �����1���U��y� @���d�v��������� ��?c*�N �r����� �q8�\� ���/�%/�Fd�MODEL 2�Skx�o(
 �<o$c (  o&�(�/�/�/�/ �/�/�/�/??d?;? M?�?q?�?�?�?�?�? O�?ONO%O7OIO[O mOO�_�Oy/�O�O&_ �O_\_3_E_W_�_{_ �_�_�_�_o�_�_o Xo/oAo�oeowo�o�o �o�o�o�o�O�O�O /����� ����P�'�9�K� ]�o���Ώ�����ۏ ����#�5���Y�k� ��Se��������� ��1�C���g�y�Ư ������ӯ���D�� -�z�Q�c�u������� ��Ͽ�.�ɟ۟	�� ���qσ��ϧϹ�� ����<��%�7߄�[� mߺߑߣ��������� 8��!�n�E�W��?� Q�cϑ��y�����F� �/�|�S�e�w����� ��������0+ =Oa����� ����>��� ]o������ ��/#/p/G/Y/�/ }/�/�/�/�/�/$?�/ ?Z?1?C?U?+�?O }?�?�?�?�?2O	OO hO?OQOcO�O�O�O�O �O�O_�O__d_;_ M_�_q_�_�_�_�_�_ �?*o�?�_oroIo[o �oo�o�o�o�o�o& �o\3EWi{ �������� �/�A�o��;oi�{� 菿�я�����+� =�O���s���ҟ���� ͟ߟ��P�'�9��� ]�o������������ ��߯�^�5�G���k� }���ܿ��ſ���� H��1�Cϐ�g�y��� �ϯ���������D�� -���'�U�g���O� ���������R�)�;� ��_�q������ ����<��%�7�I�[� m����������ߝ��� ��J��3EWi{ ������� /|Se��� ����0///f/ A/S/�/;/�/�/ ?�/�/>??'?t?K? ]?o?�?�?�?�?�?�? (O�?O#OpOGOYO�O }O�O�Ow/�/�/�O�O �O_1_~_U_g_�_�_ �_�_�_�_�_2o	oo ho?oQocouo�o�o�o �o�o�o�Ov _?Q'���� �*���%�7�I�[� �����ޏ��Ǐُ� ���\�3�E���i�{����Җ�$DCSS�_PSTAT ������Q    l�� � (&��K�2�o����  ������$�˟į֯���� �����'���SETUP 	N�Bȶ��� X�r���������ۿ��g��T1SC �2
K����Cz��#�5�G� �CP [R�D$�Dl �Ϥ�^�����ϻ�� "�4�F�X�j�|ߎߠ� ������������0� B�T�f�x������ ��������,�>�P� b�t������������� ��(:L^p ����~����� �-�Qcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �__/_BS_e_w_ F_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o���� �����#�5�G� Y�k�}�������ŏ׏ �����1� _U�g� y��_����������� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W� i�{�J��߱�ğ���� �����/�A�S�e�w� ������������ �+�=�O�a�s����� ����������' 9K]o���� ����#5G Yk}������ ���/1/C//g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_�!o3oEoX/ io{o�o\o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� ok�}��o^���ů�� �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ����������%�7��I�[�m����$D�CSS_TCPM�AP  ������Q W@ ������������������	��
������������W�  �������������R��⡋�����U��������U ��!��"��#��U$��%��&��'��U(��)��*��+��U,��-��.��/��U0��1��2��3��U4��5��6��7��U8��9��:��;��U<��=��>��?���@��UIRO 2]������� ����0BTf x�������,1��U�� y������� 	//-/?/Q/c/u/�/ �/�/6�/Z�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O �/[O�/O�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_NO�_���UIZN 2.��	 �����(o :oLoR�%ozo�o�oao �o�o�o�o
.�o RdvE���� ����*�<�N�`� #�����e���̏ޏ�� ���&�8��\�n��� C�����ȟ������ ӟ4�F�X�'�|����� c�u�֯请���0���_��UFRM R�������w��� ������ѿ����� +�=�O�a�sυϗϩ� ����������'�9�K�\�r��\߄ߖ� qߺ��ߧ������&� 8��\�n�I���� ����������4�F� ]�o�|���-������� ������0Tf A��w���� �>Pg�t� %������/ (//L/^/9/o/�/�/ �/�/�/�/ ??�/6? H?_l?~??�?�?�? �?�?�?�? O2OOVO hOCO�O�OyO�O�O�O �O
_�O._@_W?d_v_ _�_�_�_�_�_�_�_ o*ooNo`o;o�o�o qo�o�o�o�o�o& 8O_!n��� �����"��F� X�3�|���i���ď�� ���Տ�0�B�Yf� x��������ҟ䟿� ����>�P�+�t��� a�����ί����߯ (�:�@�