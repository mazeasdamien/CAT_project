��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ���ADV_IN� �0   � OPE�N� CRO ?%$CLOS� $��AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�o#IN_;OU�FAC� g�INTERCEP�fBI�IZ@����ALRM_R�ECO>""AL]M�"ENB���&sON�!� MDG/� 0 $DEBUG1A�"d�$�3AO� _"��!_�IF� � �$ENABL@�t#� P dt#UE5K�%1MA�s �"�
�� OG�f J0CU�RR_u1P $�3L�IN@�1z4$t$AcUSOK4� OD2�$SEV_AND�_NOA 3PPI�NFOEQ/  �L �0p1�5�1_ H �749�EQUIP 3�@NAM0��,B_OVR�$VERSI� ��!PCOUPLE] � 	 $�!PP�1CES0�2eG � OC> �1
� � $SOF�T�T_ID�2TOTAL_EQ 0��1�@N" �@U SCPI
 �0^�EX�3�CRE -DdBSIGJ@dOvK�@�PK_FI90�	$THKY"WP�ANE�D � D_UMMY1dIT�1TU4QQNU�A�Rx1R� � _$TIT91�  ��� �Td�T0�ThP��T5�V6�V7�V8
�V9�W0�W�WOQ�UP�WgQ�U�W1�W1�W�1�W1�W2�R�S�BN_CF�!@$<!J� ; ;2��1_CMNT�?$FLAGS]��CHEK"$�b_�OPTJB� � EL�LSETUP 7 `@HO8@9 �PR�1%�c#�aR'EPR�hu0D+�@���b{uHM9 M�N�B;1 UTO�BJ U�0� 49DEVIC&�STI/@�� �@�b3�4pB�d�"VA�L�#ISP_UN9I�tp_DOcv7�yFR_F�@|%u1�3��A0s�C_W�A�t,q�zOFF_�T@N�DEL�L�w0dq�1�Vr?^q�#S?�o`Q"U1�t#*�QTB��A��MO� �E 	� [M�����wREV�BIL����XI� v�R � !D�`��_$NOc`M� |��0��ɂ/#ǆ�� ԅ���!X�@D�ed p E R�D_E��h�$F�SSB6�`KBD�_SE�uAG� G
�2Q"_��2b�� V!�k5p`(��C� 0q�_ED� � �# t2�$!S�p-D�%$� �#�B�ʀ_OK1��0] P_C� ʑ0t��U ^�`LACI�!�a��Y�� �qCOMM� # $D
� ��@����J_\R�*�BIGALLOW�G (Ku2-B�@VAR���!�AB ��BL�@� � ,�K�q���`S�p�@M�_O]˥��C?CFS_UT��0 �"�A�Cp'��+pX�G��b�0 4� I'MCM ��#S�p��9���i �_�"t�  ��M�1 h�$�IMPEE_F �s��s��� t��F��D_�����D��)F����_����0 T@L��L��DI�s@G�� ��P�$Ix�'�� �CFed7 X@GRU@�z�Mb�NFLI�<\Ì@UIRE�i4<2� SWITn$`0k_N�`S 2CF�0=M� �#u�D��!��v`����`%J�tV��[ E��.�p�`�ʗELBOF� �շ�p`0 ���3����� F�2T�`�A`�rq1J1��z _To!��p���g���G� �>r0WARNM�p#t�C�v`�ç` � CO�R-UrFLTR^��TRAT9 T%p>� $ACCVq���� ��r$ORIX�_&�RT��S<���0CHG�0I����TW��A�I'�T��!D��� ��202�a1��HDR�2��2�2J; S�᪭�3��4��5��6*��7��8��9 1m�x׀
 �2 @� TRQ�$vf��'�1�<�_U<�G� {COec  <� �P�b�t�53>B_�LL�EC��!~�MULTI�4�"u�Q;2�CHILD��;1���@T� "'�S�TY92	r��=��)�2���EN��ec# |r056$J ���`���uTOt���E^	EXTt�����2��22"(M����$`@D	��`&��p����� %�"��`%�ak�� ���s!���&'�E��Au��Mw�9 �%� ��TR�� ' L@U#9 ��z�At�$JOB��x��P�TRIG��( dp������^'#j�~�x�pO�R�) t$�F�L�
RNG%Q@�TBAΰ �v&r�*`1�t(��0 �x!�0�+Pd�p�%�Q!��*�Ё͐U��q�!�;2J��_R��>�C<J��8&<J D`5C�F9���x"�@J�?�Pq_p�7p+ \@�RO"pF�0��IT�s�0NOM��>Ҹ4Ps�2�� @U<PPg�*��P8,|Pn��0b�P�9�͗ RA����l�?C�� �
$T\ͰtMD3�0T���pU�`�΀+AH,lr>�T1�JE�1\� J���PQ��\Q��hQC�YNT�P��PDB�GD̰�0-���P�U6$$Po�|�u�AqX����TAI�s7BUF,�tp�C�1�. ����F�`PIV|�-@PvWMuX�M�Y�@�VFvWSI�MQSTO�q$7KEE�SPA��  @?B�B>C�B�A��/�`=��MARG�u2��FACq�>�SLEW*1!0����
�6�2MCW$0'����pJB�Ї�qDE�Cj�e�s�V%w1 Ħ�CHNR�;MPs�$G_@�g�D�_�@s��1_FP�5�@TC�fFӓC@�Й���qC��+�VK��*��"*�JRx���SoEGFR$`IOh!v�0STN�LIN>�csPVZ�ذ�Ц@�D2����r 2��hr�r�� P��3` +^?���եq�`��q�|`�����t��|aSCIZ#�!� �T�0_@%�I��qRS� *s��2y{�Ip{�pTp�LF�@�`��CRC����CCTѲ�Ipڈp�a���b��MIN���a1순���D<iC �C/���!uc���4�Ln j�EVj���F��_!uF��N����|a(��=h?KNLA�C{2�AVSCAB�@A��2�@�4�  cSF�$�;��Ir �3�a�05��	D-Oo%g��,�,m����ޟ�2R>C�6� n����sυ�U��R�0HA;NC��$LG��ɑ6DQ$t�NDɖ��AR۰N��aqg�����X�ME��^�Y�[PfS�RAg�X�AZ��蟸��rEOB�FCT ��A��`�2�!Sh`0ADI��O��y�" y�n!�������~#C�qG3�!��BMPmt�@�Y�3�afAES�$�����W_;�BA�S#XYZWPR$��*�m!��	VQU�87  ƀI�@d���8\�p_C�:T���#��� Rs_L
 � 9 ����C�/�(zJ�LB�$�3�D��5��FORC�b�_A�V;�MOM*�q�SaԫBP`Ր�y�HBP��ɀE�F����AYLwOAD&$ER�t&3�2�Xrp�!��R_FD�� :� T`I�Y3��Ed�&��Ct��MS�PU
$(kpD���9 �b�;�B�	E�VId�
�!_7IDX2$����B@X�X<&�SYn5� �_H�0�e�<��ALARM(��2W�rt�_�0�= h�@Pnq�`M<\qJ@$PL`A&�M#�$�`��� 8Ѡ	���V�]�0��1U��PM{�U��>�T[ITu�
%�!�[q�BZ_;���? ŔB pQk��6NO?_HEADE^az� �}ѯ��`􂳃���d@F�ق�t4���@���@��uCIRTRH�`��ڈL��D�CB@64�RJ��p�[Q����A�2>���ORĭr��O����T`UN3_OO�Ҁ$���P�T�����I�VaCzx�� PXWOY�z��B�$SKA�DR��DBT�TRL��C��րfpbD�s��~�DJj4 _��DQ}��PL�qwbWA���WcD�A��A=�2��UMMY9��1�0��`DB����D�;[QPR���`9�qD�Z���E OжY1$�a$8���L)F!/_c��R�0GG/Y$C�1Hf/~���PENEA@�Tf�I�/��%�R�ECOR`"JH� @ �E$L�#F$#PR���+jp���nq�_D$�qPROSS]�
���R�r�|` u�$TRIG�96PAUS73ltE�TURN72�MR�:�U 0Ł0EW�$��SIGNALA�QR$LA�З5�1�G$PD�H$�Pİ�AI�0�A�C�4�C��DO�D�2��!�6GO_AWAY2MOZq�Z��W DCS��CSCBg�K Իa#���WERI�0Nn�T�`$�����FCBPL�@QBGAGE���P���ED|BD�wA[CD�OF��q[F0�FoC��MP�MAB0XoC�$FRCIN��2Dk��@���$NE�@�F�DL8�� L� ����=��Rw�_��}P� OVR10����lҠ�$ESC�_�`uDSBIO����pTe�E�VIB�� `s��Z��V���pSSW��$�V	L��:�Lk��X����`��bQ����USC�PⓂA=�	Q��MP1�%e&S*`�(bt`'c5۳ESUd��-cWg &SWg?cWd����Wd��xWd.���AUTO$�0Ya҃�ac�SB���� -d��&SwB[��GB�f�$VOLT�g ��  �GAOD�!�q���@:�OR�QҀKra�$DH_THE&0�Rgpx� qtnwALPHnt��o��w0 Vp]�$�.�Ra�[��s�5�`r�HCQ#BUD�S� F1	M��sV
��;���Lb�tk���BRT#HR��L��T`�Z�
�Vɖ��SDE  �1��2�� ����������kѯ� aәTt0V�ꆸ�������̈Я�-�"�N�~��sS2����INHB��ILTG0ɡ�T ?��3$�w��E��PqQ�xQ�TqPe��0Y�AF}�O�ນ�� ڗ��qPڳē����bPܙ���PL?���3���TMOU��ēS� ��� ��s�/�S18���O�Aܙ��I����C�DIƑ˩o�STI��գ�O:ҋ�,0���AN��Qg�S��+r�#x$�����bw�_����PRA�P�`vC����MC�NeQe�����VECRS��r�oPIw�AFPåǲШ۷G.��DN��G>�����F��2�Ƿ�M�7�F*��_�MN�D̠,�����d�{ƭa����O�B���U˱z���DI���#���3�����A���w�Fx���3��ON�5��Q��VA�L�CR[�_SI�Z��b���n�REQ��Rb��]2b���CHq�΂�ڃ�Ռ�����:�n�S_U��X��.wWFLG���wU/$CV�iMGP�QδFLXP�923R楘u���EAL�P-�C(	��+rT��W��� �R�c���NDM�S7� ��K>S�P_9M'0h�STWv������AL�P���Q����U���U�IA�G,�o��d�U�-�T"A-`� ���A��@���H`��Q`��6��Pq_D&��1s��.@�P�F�>2�T�� ?7 1A>М�#�#L��?�_=i @@>LD��c���0�FRI�0 `Ѐ��1}��IV\1�*�^1�UP`��a��C�CLW��
`L=S &-c&&S�C.w� � L���!����d�QB$w�҇��$w�����
�P�5RSM����V0h � �r��d^2AW�a_T�Rp}�8@NS_P�EA����< ��$�SAVG�8�6G]%���CAR �`�!�$���"CRa���$ d�#E�@��"STDă��!Fpo��'QOaF��%��"RC���&RC۠�(F�2A�R`#7���%, gMA�Q_�a��
QQ��al2J��u4Ib�r7I�R �9wQ�7�8M/��!uCpR�  �p:�2F<�SDN�a�   W2QM P $Mi��s$c A�$C�cm�9���4�AT�0CY_� N LS!IG�1x'yB��y@@H2�Y�NO����SDwEVI�@ O@�$�RBT:VSaP�3�CuT�DBY|��A	W`3CHNDG�DAP H@GR%P�HE iXL�U��PVS�Fx2� CL1p� Q6ROp��F9B�\]�FEN�@��S��ChAR d��@DOd�PMC�Sb�P薇P�R��HOOTSWz42�DMpGELE�1/e�9C8`�RS T�@���r�� hf��`OL�GH�A�Fk�Fs������C�A@T � �$MDLUb 2S@�E���q�6�q�	0�i�c�e�cJ��	�uݢ�#~5t+w�PT�O��� �byU�TS�LAVS� U  ��INP �	V��t�yA_;�ENUAwV $R�PC_�q
�2 1bL�wpp�R�p�SHO+� W  ���A�a�q�2�r�v��u�vS_CF� ?X` ,f��r�OG gE��%D�h���pC�Iߣi�M�A��D�x AY?�W�� p�NTV	�D�V�E�0@�SKI��T��`g?Ň2�� JZs�! Cꆻ��f��_SV� �`XCL�U��H���ONLd��'�Y�T��OT:e�HI_V,11 AP7PLY��HI4`;��U�_ML�� $VRFY8�	�U�=M{IOC_I���"J 1"��߃O�@X��LSw"`@$DUMMY4���ڑ�C=d L_TP���8kC��^1CNFf��@�E��@T�y� D_#�UQ_��ݥ�YPCP���=�� ������aD���� Y �+�
0RT_;P��uNOCCb Z�r�TE���=�פr�TG�@[ D��P_BAe`Lkc�!��_���H��u�� �\�pAb=cARG�I�!$���`[ �Md_SGNA]� ��`U��IGN��Տ��� ��V�������ANNUN���&�˳�EU�J'�ATCH��J��8�d�rA^ <@g������:c$Va��`����qqEF] }I�� _ @@�FͲITb�	$TOTi �C�O�cͶ @EM�@NI�aQ`tB��c���A>����DAY@CLOA�D�D\�n����q��[EF7�XI�Ra���K���O%��a��ADJ_R�!@b"��>�H2�"[�
 Hc�%��`a͠MPI�J��D�A��?�Ac 0��х�� �ђZ�ϡ�Ui ���CTRL� Yp �d��TRA8 ?3I?DLE_PW  ��h���Q��V�GV_���`c �o�;Q@?e� 1$��6`<cTAC-3��P�LQH�Z�Rz\ A-u6:ɰSW;�A \���"J��`b�K�;OH�(OPP; �#�IRO� �"BRK��#AB ���� ���� _ ���F���`�d͠, j@S�RQDMW��MS�P6X�'�z��IFECAL,�� 10^tN��V―�豊�V�(0��C)P
��N� Yb� !gFLA_#�OVL ��HE���"SUPCPO��ޑ\�L�pH��&2X�$Y-
Z-
W-
��/��0�GR�XZ�q�$Y2&�CO�PJ�SA�X2 R��*r�!��:��"�RyI�0)�f `�@/CACHE��c؛�0�s0LAZ SU7FFI, C��q\���6o�NaM�SW�g 8�K�EYIMAG#TM�@S��n
2j�r|!�bOCVIE���~�h �aBGLx����`�?� 	qqԚ��i��!`STπ!�����������EMAI��`N��`A�PZ�FA�U� �j�"�q�a��U�3��� }�?k< $I#�U�S�� �IT'�BU!F`��DNB���'SUBu$�DC_���8J"��"SAV�%�"�k������';��P��$�UORD��UP_pu �%��8OTT��1_B`��8@LMl�F4���C7AX@Cv���XXu 	��#_G��
�P'YN_���l6���UD�E��M����T��F� caC�D]I`BEDT)@C���~�m�rI�G�!c�&���l`��-�P��F�ZP n (�pSV� )d\�ρ���QA~��o� �����>"$3C_R�IAK��kB��hD{pRf8gE.(ADSP~KBP�`�IIM�#�C�Aa�A��U�G���iCM! IP��KC��� ��DTH� �S�B*�T̤�CHS�3�CBSC��� ��V�dYVSP��#[T_DrcCONV�Grc[T� �Fu 	F�ቐd�C�0j1���SC5�e]CMER|;dAFBCMP;cv@ETBc p\�FU DUi ��+�~�CD�I%P70�2#9�EO���qWӏ�SQ��QǀSU���MSS�1ju�4`�T�aAa��A�1r�� "�з��4$Z!O@s���l�U6�&�2�eP���eCNc�l�x�l�l�iGROU�Wd)��S c�MN�k Nu�eNu�eNpR|b|�i��cH�pi��z
 �0CYC���s�w�c�6�zDEL�_D��RO�a���qVf���v{�O�2���1��t���:R�ua�.#��&��AL� �1sˢI1¡�J0�PB���G��ER^�T�Gbt �,!@��5��aGI1L~cR1s 
HO������1u��������R�P����Cڠ	�<����DMA��J0��0vH *	�L U�1#J�Q��V
�[�7A z���z��z��z�Ѩz�Fz�7w�8w�9Pw���y���1��1��U1��1��1Ě1њU1ޚ1�2��2�����2��2��2��2�Ě2њ2ޚ2�3J��3��3����3��U3��3Ě3њ3ޚe3�4���2XTF��1w6�.(�0�f�0�U�0ŷ�e��FDR�5�xTU VE���?1���SR��REr�F���OVM~Cz)�A2�TROV2ɳDT� R�MXa�I�N2���Q�2�IND�p�r�
���0�0�0G@u1��[�G`��{�D_֎[�RIV�P��G�EAR~AIOr�K"N�0�y�p�5`�@�a�Z_MCM�� �����UR�Ryxǀ��!? ���p?nЋ�?n�ER�v�=a�!�P���zI:�PXqB�R�I0%�`�#ETUP?2_ { ���##TDPR�%TBp��p����3���BAC�2G| T��"�4)�:�%	`^B��p�IFI��� Mc���.��PT��!FLUI�} � ��K UR�c!���B�1SP�x E�EMP�p�2$���S^�?x��J8ق0
3VRT���0_x$SHO��Lq�6 ASScP=1��PӴBG_���������FOR�C3"f�d~)"F%UY�1�2\�2
A���h� p� |��N�AV�a��������S!"��$VI�SI��#�SCM4S�E����:0E�V�O���$���M����$��I��@��FMR2��� �5`�r�@ �� �2�I�9 F�"��_���LIMI�T_1�dC_LM�������DGCLFl����DY�LD����5�����ģ� �����u	 T�sFS0Ed� P���QC�0$EX_QhQ1i0�P�aQ53�5��GoQ��g� ����RSW�%�ON�PX�EBUG���'�GRBp�@U��SBK)qO1L� ��POY 
)�(�P��M��OXta`�SM��E�"me�����`_E �� 
@����TER�MZ%�c&��ORI��1_ �c' �SM�epO��_ �c%�����`�(��)UP�>� �� -����b���q#� ����G�*� ELTO0Q�p�0�PFIrc�1�Y��P�$�$�$U;FR�$��1�L0e� OTY7�PT�4q�k3NST�pP�AT�q4PTH	J�a`EG`*C�p1ART� !5� y2�$2REL�:)ASHCFTR1�1�8_��QR�Pc�& � $�'@�� ��s�1 @�I�0�U�R G�P�AYLO�@�qDYN_k���.b�1|��'PERV��RA��H ��g7�p�2�J�E-��J�RC���ASY�MFLTR�1WJ*7����E�ӱ1�I��aUT�pbA�5��F�5P�PlC�Q1FO5R�pM�I!���W��/&�0F0�qr� H��Ed� �m2XN���5`OC1!>?�$OP�����c�����bRE�PR.3�1a���3e��R�5e�X�1>(�e$PWR��_���@R_�S�4��et�$3UD��N�Q72 ����$H'�!^�`ADDR�fHL!�G�2�a�a�ae��R���U�� H��SSC����e-��e���eƪ�SEE���HS{CD��� $����P_�_ B!rP􍀌���HTTPu_��HU�� (��OBJ��b(�$��fLEx3Us��� � ���ะ_��T?#�rS�P��z�sKRN�LgHIT܇ 5��P���P�r������PL��PSS<�ҴJ�QUERY_FL�A 1�qB_WEBwSOC���HW��1U���`6PIN'CPU���Oh��q�����d���d�������IHMI_ED^� T �RH�;?$��FAV� d�~Ł�IOLN
◓ 8��R�@�$SLiR$INoPUT_($
`���P�� %ـS�LA� �����5�1��C��BmQI�O6pF_AS7��$L%�}w%�A��\b.1�����T@HYķ�����g�wUOP4� `y� ґ�f�¤�������`PCC
`����#��>�QIP_ME��7� Xy�IP�`�U�_NET�9����Rĳs�)��DSaP(�Op=��BG`��T���M�A��� �l�:CTAjB�pAF TI�-U��Y ޥ��0PSݦBUY IDI�rF ��P��a��� �y0�,�����Ҥ�NQ�Y R���IRCA�i� ך ěy0�CY�`EA�����񘼀�CC����R�0�A�7Q�DAY_���NTVA����$��5 ����SCAd@��CL@����.��𵁛8��Y��2e�o�N_�PC P�q��ⱶ��,�N� ���
�xr���:p�~N� 2� ؀��(ᵁ����xr۠�LABy1��Y ��U�NIR��Ë IT!Y듭��ed�R#�5����R_URLގ��$AL0 EN���ҭ� ;�T��T�_U��ABKY_z��2DISԐ�A�C�Jg����P�!$���E��g�R���"� A�/���J����FLs��7 Ȁ����
�UJR� ���F{0G��E7⬙�J7 O R$J8I�7��R�d�7��E�8{�H�A7PHIQS��=DeJ7J8B���L_KE*�  ��K��LM[� o� <X�XRl��u���WATCH_�VA��o@D�tvFIELc��cy�`��4� � o1Vx@��-�CT[�9�m�q�L�GH��� $~��LG_SIZ�t��z�2y�p�y�FD��Ix���+!��w�\  ����v��S���2�� p�������\ ���A�0_gCM]3NzU
RFQ\vv�d9(u�"B��@2�p����I���+ �\ ��v�R�S���0  �ZIgPDUƣE�LN=�
��ސ�p�z6� ��f�>sD�PLMC7DAUiEAFp���TuGH�R�q|��BOO�a��3 C��I�IT+��̦`��RE���SC�R� �s��DI��S�F0�`RGIO"$D������T("�t|�S��s{�W$|�X��J{GM^'MNCH;�&|�FN��a&K�'u�ƅ)UF�(1@�(FW�D�(HL�)STP��*V�(%Г(��(RES9HIP�+��C[T@�# R��&p:'^9U=q��$9'�H%C𜓚"Gw)�0PO�7�*��#�W}$���)EX��TUI�%I���Ï�����rCO#C� *�$	S��	)��B@�;NOFANA|��Q�
�AI|�t:��ED�CS��c�C�c�BO��HO�GS���B�HS�H(IGN�����p�!O���DDEV<7LL�� �-���i�(�;�T�$���2�p���	��#A����(�`�{�Y��PO+S1�U2�U3�Q��8�2�@�Ш ��{�PtD����&q)���0�d��VSTӐR�Yl�\@ ` �$E.fC.k�p<p�=fPf�?��4�ѩ LRТ� ��x�c�p���<�Fp�dY�@!�_ � ��7Lpx&���c�MC7�� ��CLD�PӐ��TRQLI0#ѽ�ytFL��,r��5s8�D�5wːLqD5ut5uORG���91HrCRESERAV���t���t�� �c~�� � 	u095t5u��PTp���	xq�t�vRCLMC�������q��M��k�������$DEBUGMA�S��ް��?U8$T�@��Ee�g����MFRQՔ� �� j�HRS_KRU��a��A���k5FREQ� �y$/@x�OVER�С�n��V#�P�!EFI�%�a��g�I9���t� \R�ԁ�d�$U�P��?��p�PS�P��	�߃C��͢a��U|\�l�?( 	ha�MISC� d�@�QRQ��	��TB � Ȗ0A՘�AX����ؗ�EXGCESj�	᫒M��
\�������԰Q���SC�P � H��̔_��Ƙǰ]�����KHԳK�J� �m�B_K�FLIC��dB�QUIREG3MO��O˫3�q��ML�`MGմ @�`��T���a#NDU�]��>���k�G�Df��INAsUT���RSM>�a��@N)b]3-��p�5�PSTL\�� �4X�LOC�VRI�%��UEXɶANG�uBu�R�ODA��ŷ�������MF O����Y�b@�e4��2k�SUP�fTAw�FX��IGG� � ��p�c ���cQ6�dD�%�b|� !`��!`��|��3w�ZW�a�TI��P;� M���[�� t��MD
��I�)֟@����HݰM��DIA�����W,!�wQ�1*�D�)��O���n]�� 0�CU��VP��p��O!_V��ѻ ���S�LX�5������P��h0N���P��KES2���-$B� �����ND2����2_{TX�dXTRA�C�?�/��M�|q�`�Pv��XҰ�Pt �SBq`�USWCS��T��	���PULYS��A�NSޔ��<R��JOIN��H��~`j�=��b��b�����P=��$��b$���TA����S���hS�HS�E��SCF�b��J��R��PLQ�o ���LO�b�н.���^����8�������0�RR}2��� 1��zeA�q d$��IIΐ+�G�A2+�/� �PRI�N�<$R S�W0"�a/�ABC�D_J%�¡u���_J3�
�1S�Pܠe�u�P��3P��р`u��J/�(��r�qO8QIF��CSKP"z{�{�J���QL28LBҰ_AZ�r��~ELQ��OC�MPೕ�T���RT�����1�+���P�1��>@�Z�ScMG0��=�JG�`�SCL�͵SPH�_�@��%V�u� RTER`  �< A_�@G1"�A0�@c��\$DI�
"�23UDF  �ǀ~ LW�(VEL�qIN�b)@� _BL�@u��$G�q�$�'��'�%`<�� ECH<ZR/�TSA_`� K���E}`<����H5�Bu��1}`_�� �)5D2d%��A4bI��N9t&R�DH�tA���ÀP$V `�#>A$��łV�$Q��R}�����H �$B�ELvᵆ<!_AC�CE�!c��7/��0I�RC_] ��pNyTT��S$PS�rL� d�/Es��F {�@F
��9gGCgG36B���_�Q�2�@p�A���1_MGăcDD�A]"łFW�`����3�EC�2�HDE>�KPPABN>G��SPEE�B�Q%_p�B�QY�Y��11$U�SE_��,`Pk�C�TReTYP�0�q P�YN��Ae�V�)хQM���ѷ��@O8� YA�TINCo�ڱ��B�DՒ�WG֑ENC����u�.A�2Ӕ+@/INPOQ�I6Be���$NT�#�%NT�23_�"łIcLO� ł_`��I�_�if�� _�k�? �` ej�C<400fMOSI�A���ОA䃔�PERCGH  �c��B" �g ��c��lb=������oUu@�@	A6B(uL eT	~�1eT�ljgv΂fTRK@%�AY ��"sY��q6B�u�s۰p�]��RU�MOMq�ՒY�MP�^��Ca�s�CJR��DUF ��BS_BCKLSH_C6B)����f����St�H��RR��QDCLALM-d\��pm0���CHK���GLRTY���d��pY��)Üd_UM]��ԉC��A!�=PLMT� _L�0��9��E�.� ��#E )�#H� =��Q3po�xPC�axHW�頿E�ׅCMCE��@�GC�N_,ND�Ζ�S	F�1�iVoR��g<!p��6B���CATގSH)�,�DfY���f��7A���܀PALބ�R_P݅�s_� �v���s����JG�T]���Y�����TORQUaP��c�yPOU��b��P%�_W�u�t��1D�P�3C��3C�IK�IY�I�3F�6�����@VC�00RQ�t���1���@ӿ��ȳJRaK�����UpDB �M��UpMC� DL�1BrGRVJ�Cĭ3Cĳ3$�H_��"�j@�q�COS~˱~�LN���µ�ĭ0���@��u����̓��Z���f$�MY��؊��|��>�THET0reNK23�3hҧ3��[CBm�CB�3C! AS� ��u��ѭ3���m�SB�3��x�GT	S$=QC������x�����$DU��@Kw�B�%(��%QqA_��a��x�{�K���b(��\�A`Չ��8p�{�{�LPH~�g�Aeg�Sµ��������@g������֚�V��QV��0��V��V��UV��V��V	�V�V%�H��������G�T����H��H��H	�UH�H%�O��O��OV	��O��O��O���O��O	�O�O�Fg���	������SPBALANC�E_-�LE��H_`�SP!1��A��|A��PFULCE`lTl��.:1���UTO_����T13T2��22N���2 9`�!�qnL�=B�3��qTXpOv 
A4�I�NSEG�2�aREqV��`aDIF�ufS91�8't"1�6`COB.!t�M��w2��9`��,�LCHWA�RRCBAB�� �@�#�`-ФQ 5�X�q�PR��&��2�� �
�""��1eROB�͠CR6B5������C�1_��T �� x $W�EIGH�P`$Ȝ�?3àI�Qg`IF�YQ�@LAG�Rq�S��R �RBILx5O1D�p�`V2ST�0V2P!t�W0�11�&1/0��30
�P�2�QA � 2řd[6DEB�Ug3L_@�2�M'MY9&E Nz�D�`$D_A�a$��0��O� ��DO_@A.1� <B0�6�m�Q�IB�2�0N-cdH_p`�P �2O�� �/� %��T`"a���T/!�4)@TICYKh3| T11@%�C� ��@N͠�XC͠R�?��Q�"�E�"�E8@P�ROMP�SE~� $IR��Q��8R;pZRMAI)��Q4�R4U_r02S; t�q�PR8�COD�3sFU�Pd6ID_[��vU R!G_SU;FFu� l3�Q;Q�BDO�G �E�0�FGRr3�"�T�C �T�"�U�"�Uׁ�T8D��0�B0Hb _FIv�19*cORD�13 50�236V�+b|�Q1@$ZDT}U�s0�1;E�4 *:!L_NAmA�@�b>�EDEF_I�h�b �F�d�E�2�F�4�F�c�E�e�FISP��PAKp�Ds�C�d��44בi��2D�"�It��3D�O#OBLOCKEz��S�O�O�Gq�R�PUM�U�b�T �c�T�e�T!r�R�s�U �c�T�d�R�6�q�S � ���U�b�U�c�S�Z��X�@P` t�@qDe�)@W�x���s 1�TE�<D�( }l1LOMB_���ɇ0V2VIS;�I�TYV2A��O�3A�_FRI��a SIq�QR�@��@R�3�3V2W��W��4����_e��QEAS^3�Rϡ��_�[p:R��4�5�6_3ORMULA_Iz����THR^2 �EGtg�30f��<8�5COEFF_O�A�	 ��A��GR�^3S�g0BCAnO/C$���]3 1�0GRP� � � $�p4�YBX�@TM~w��`�u�B�s��bCER, qTttsd�0�  ��LL�TSpS~�_SAVNt�ߐ���0�8 ���0� ��SE;TUsMEA*P�P౰W0�1+b/0� �3 h��  @ڐ@o�l�o�cqz��b�@$cqq`tP�G��R�� Q\p*q[p��>�:c NPREC>at���ASK_$|��� PB11_USER����{ ���VEL���{ 0��$Ō!I]`��MT�ACFG��� � �@@ O�"NO�RE-0l@o�V�SIb.1�d��6�"UXK��fP!��DE�� �$KEY_�3>�$JOG��0SV������!��}��SW�"�a\aS�ՐT�|�GI���| ^�� 4 h��'d2�!XYZc���3�1�_ERR#��! 8Ԡ�AfPV�d���1����$BUF��X��!0�MORn|�� HB0CUd� lA�!��GQ\aB�,"!aO$� ���aП���?�G~�� ?� $SIՐ����VO��T�0OB�JE_��ADJU<)B��ELAY���%�DR�OU.`=ղ�\�Q0b=��T�p��0���;BDIR�����; I�"0DYNHW�#���T��"R����@�0�"�OPWO�RK���,%@S�YSBUy�SO!P��ޑ�U�; 1P�pN�<�PA�t�X>�"��OP�PUd!�0�`!��l�IM�AGw�B0y�2IM�Õ�INe�d��?RGOVRD��-��o�Pq��0��J�(Os���"L�pBa���>o�PMC_Ee`�ъ�1Ny M A�21��2U���SL_���� � $OVSAL�ǫ�?q�`��2�" -�_��k�P��k@�Pu���2�C� ��`�Ź���_ZE�R�D��$G�ƀA�>���� @h*���%O~PRI��� 
JP8+��T=!/�L��ح�T� ަ0ATUS��TRGC_T���sB�� }fs�9s�1Re`���� DFAm����L����"��0a� ޱ��X�Ew{�����C0vUP��+p	qCPXP�j�43 ^��PG\���$SUBe�%�q�e9JMPWAI�T z}%LO��F<�A�RCVFBQ�@�x"�!R�� �x"AC�C� R&�B�'IG�NR_PL9DB�TB�0Pqy!BW�bP�$w�Uy@�%IG�T�PI��TNLND�&2R��rL�NP���PEED \HADOW�06�w���E[q4jO!�`SP]DV!� LbAz�p�`�07�3UNIr�ȡ�0"!R��LY�Z`� o��PH_P�K��e�RETR#IE9{�q����0v'PFI"�� �G`��0D 2�g�D�BGLV�#LOGgSIZ��EqKT�!�U��VDD�#$0_T�G�MՐCݱ��|@�eMRvC}�3�CHEsCK0���PO��V!�k�I��LE,(!��PArpT�2K��W��@P2V!� ?h $ARIBiR� c�a/�O�P8�ӐATT��2�IF|@0z�Aq4S�3UX����2LI2V!� $<g���ITCHx"[�-W �AS9�wS�LLBV!�� /$BA�DYs���BAM!���Y9F�PJ5��Q��R6�V>�Q_KNOW�Cb��U��AD�XV��0�D�+iPAYLOAt��Ic_��Rg��RgZOcL�q��PL�CL_�� !@7��b�QB��d���fF�iC֠�js��d��I�hRؠ�g�ҢdBd����J��q_J�a:#���AND��Ĳ`.t�b�aL!q�PL0?AL_ �P�0P���QրC��DNc�E���J3CpWv�{ TPPDCK�������P�_ALPHgs�sBE��gy|� �K�1�� �s ���HoD_1Oj52ydDP�AR�*���;�&���TIA4�U�5U�6��MOM���a���n���{�Y�B� ADa���n���{�PUB��R��҅n��҅{���2�Wp��W �/  PMsbT�� /wR���?� e$PI��81���TgJ��niJ�I
V�Id�Ir��[��3!��>!��r�Ӫ�U3HIG�SU3�% �4얎4�%� ���"�����!
��!�%SAMP���^��_��%�P4s ю���[  	ӝ�3 ���0���&��C�����^��Sp��H&0	�IN�SpB��� �뤕"��6��6�V�/GAMM�SyI�F� ETْ��;�D�tvA�
$ZpIBR!�62IT�$HIِ_����C�˶E��ظAҾ���LWͽ�
̀��7���rЖ,0�qC��%CHK��" �~I_A����� Rr�Rqܥ�Ǚ��ԥ�|��Ws �$�x� 1���I7R�CH_D�!� R1N{��#�LE��ǒ�!,��x���90MS�WFL�$�SCR�((100��R@��3 ]B��ç��a����َ0ޤ�PI3A9�ME�THO����%��AXH�XX0԰62�ERI��^�3��R$�0$u	��pF{�_����?ⲣ1�L�L8�_�a�OOP����8wᲡ��APP:���F���@{���أR	T�V�OBp�0T���0�;��� 1�I���� ��r���RA�@MeGA1P�SSV-�w�P_@CURg��;�GRO[0S_�SA�Q��Y�#NO�pC!"�tY�� Zolox�������!b��,��&�DO�1A���A ����Х��A���A"�0WS�c P�Q}M)�� � �ãYLH�qܧ��S rZ�]B�o�����Ĕ�q_�C1��M_W���g���c�M� �`Vq�$Ap�x1o�3"�PMJ�,�� �'A� 9�!YWi:�$�LWQ |ai�tg�tg�tg{t� �N`���S��JSpX�0O�sRqZ���P� *�� ���M��������������pX��� ��@LNK�P:�q_~R� |�q#( Y����&n��&{�Y�Z� �'�&t��Q���0'�"J0���0}`�$PQ��PMON_QU�c� � 8�@Q�COU��%PQTH��HO�^0HYSf:PES�R^0UEI0tO��@O|T�  �0�PGõz�RUN_TO�%�0ْ.�'� PE`�5C��A�<�INDE�ROGGRAnP� 2g��NE_NO�4�5I�T��0�0INFO�1� �Q�:A����AB� (��SLEQݖFAѕ�F@�6uPOSy�T�� 4�@ENAB|��0PTION.S%0ERVE���G���wFGCF�A� @bR0J$Rq�2����R�H�O�G "�EwDIT�1� �vR�K�ޓʱE�sNU0W*XAUTu�-UCOPY�ِN\����MѱNXP\[qƯPRUT9� _RN��@OUC�$G��2�T� �$$CL<`� ����Q0M0 �P�S�@n�X�PX�QVIRTU��_�P�A� _WRK 2� e�@ ?0  �5�QMorYhJo|m |lA	�`�m�o0`��o�o�f�e�l}�a`I[ct'`BS��*� 1�Y� <7��� ����&�8�J�\� n���������ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T�f�x����� ����ү�����,� >�P�b�t���������vsrCC��LMT� v���s  dѴ�INڿ�дPRE/_EXE��)����0jP��za'`DVʽ�S�@e)�%�select_macro����k�|��qtIOCNVVB��� ��P��US�ňw���0V 1.4kP $$p��a�|�`?���0>� P�b�t߆ߘߪ߼��� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������� ��$�ѰLARM�RECOV �^�����LMDG� �Ь�LM_IF ���d  YST-�040 Oper�ation mo�de AUTO �S��ed P) �hang�(L:3)������)�;��M�_�q��, 
� ���#�>TE�LEOP ǘLI�NE 0ǑقAB�ORTEDǘJO�INT 100 1%�����$����@�$�A��AT	Aǒؑ3��גؒ��  clear�𪯼�ί��NGTO�L  @� 	 �A |���ѰP�PINFO �� f�L�^�p����  ������k� ��ۿſ�����5��`Y�C�iϏ�%���ٯ ����������'�9��K�]�o߁ߓߙ�PP�LICATION� ?t�����Han�dlingToo�lǖ 
V9.?40P/17���
883ǀ����sF0�	�549���������7DF5x�О�ǓNone���FRA�� �69��_ACT7IVE1�  �� ��  ��ڀMOD���������CHG�APONL�� ��OUPL[�1	��� >�B�T�f����CUREQ 1]
��  Tp�p�p�	��������l� ������������i�3l�p�3��^H��A��t
HTTHKY �FXv|�� *<N`��� �����//&/ 8/J/\/�/�/�/�/�/ �/�/�/�/?"?4?F? X?�?|?�?�?�?�?�? �?�?OO0OBOTO�O xO�O�O�O�O�O�O�O __,_>_P_�_t_�_ �_�_�_�_�_�_oo (o:oLo�opo�o�o�o �o�o�o�o $6 H�l~���� ���� �2�D��� h�z�������ԏ� ��
��.�@���d�v�`����������TO������DO_CLE�AN���E�NM ; �� p���९��ɯۯv�DSP�DRYRL���HI��o�@��G�Y�k�}� ������ſ׿����ϻ�MAX��,�����=�X,�<�9�<�>��PLUGG,�-�\9���PRC��Bm�Eq�6�(ϗ�O�¼��SEGF�K ���� �m��G�Y�k�p}ߏ�����LAP$� 7ޡ������+�=� O�a�s����� �TOTAL_ƈ� �_USENU$�1�� ������RGD�ISPMMC�2d�C�O�@@�1��O"�D��-�_S�TRING 1~��
�M���S��
��_ITwEM1��  n�� �������� $6 HZl~��������I/�O SIGNAL���Tryou�t Mode���InpNSimu�lated��O�ut`OVE�RR!� = 10�0��In cy�clT��Pro?g Aborj���JStatus���	Heartb�eat��MH �Faul��Aler�!/!/3/E/�W/i/{/�/�/�/ (���(����/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4OFO�/WORИ�~A �/XO�O�O�O�O�O _ _$_6_H_Z_l_~_�_��_�_�_�_�_�^PO���"`�KoEoWo io{o�o�o�o�o�o�o �o/ASew8��bDEV%n�p 9o����#�5�G� Y�k�}�������ŏ׏������1�C�PALT�-j��OD��� ����ȟڟ����"� 4�F�X�j�|�������8į֯X�GRIB��� ����6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�z�����R�-��&��������� �"�4�F�X�j�|ߎ� �߲�������������PREGn�W��� 0�~���������� ��� �2�D�V�h�z����������$�$A�RG_~@D ?	������  	]$$	[]��$:	��SBN_?CONFIG��XWqRCI�I_SAVE  �$zm��TCE�LLSETUP �
%  OM�E_IO$$%MOV_H� ���REP��#��UT�OBACK� �	tFRA:\D� .D�z �'`�D�w�� �s  �25/11/29� 20:26:16D�;D���#//h��C/j/|/�/�/�/�/D�X/�/? ?(?:?L?�/p?�?�? �?�?�?�?g? OO$O 6OHOZO�?~O�O�O�Op�O�O�O���  c�_F_\ATBCKCTL.TM��)_;_M___q_8IN�Im��j~CMESSAG� �Qz| �[ODE_D� �j�XO�p�_@�PAUS6` !�� , 	��; :oHg,		2oloVo�ozo�o�o �o�o�o�o 
D.�Pz}d`TSK � mw}_CUP3DT�P�Wd�p�V�XWZD_ENB8�Tf
�vSTA�U��u��XISX UN�T 2�vwy �� 	 ����J �Ѽ� V�'��� %��D�R����T���M��l��K���_m�����z�I���;�f)���x`t�:���s������4�METV��2@��y PQ��BEc�A�_y�BߤBWl��B-��B�x���?;��>����?)"�?���W?���@ K��5�SCRDCFoG 1Yw ��� � ���%�7�I�pD�Q�	ܟ������ϯ� �Z��~�;�M�_�q��������6���FGR`9��p�_ԳPNA� �	FѶ_E�D�P1��� 
� �%-PED�T-¿ R�v���AE�<�GE�D�;�9/�>���  ����2�����B� � ���{�����j�����3��#� �G�Y���G� �ߠ�6�����4�W������Zݨ��Z�l������5K��ߘ� �Y�t���&�8���\���6��d��Y�@@����(��7� S0wY�w��f���8����{�IZ��C/��2/�B��9{/��//LZ݀�/?V/h/�/�/��CR���?�?Tn?�?� ?2?�?V?԰!�NO�_DEL�ҲGE?_UNUSE޿д�IGALLOW �1�   (�*SYSTE�M*��	$SERV_GR[�@`7REG�E$�C����@NUM�J�C�M�PMU?@��L�AYK���P�MPAL�PUCY'C10 N3^P!^YSULSU_�M5R�a�CLo_�TBO�XORI�ECUR�_�P�MPMCNmVV�P10I^>�PT4DLI�p�_��I	*PROGR�A�DPG_M1I!^Ko]`AL+ejo�Te]`B�o�N$�FLUI_RES�U9W�o�O�o�dMR�N�@�<�?�;M _q������ ���%�7�I�[�m� �������Ǐُ�����!�3�E�W�2BLA�L_OUT ��K���WD_AB�OR:PcO��ITR_RTN  �$��빸�NONST�O�� lHCC�FS_UTIL ��̷CC_A�UXAXIS 3$� h}�j�|������ƽCE_RIgA_I`@�נ���FCFG �$�/�#��_�LIM�B2+�� �� � 	��B�\���$� 
Ԡ�V�)�Z���/�����[�����.R���!$�����L��(
5������PA�`GP 1H�����A�PS�e�w�6�CC� �C7��J��]��p�������� C�����������������é�̩�ձ�ߪ���������;L���PCk�������U�������������ɱ���������� D� D�!�!�!�!� m��&?��HE@�ONFIpC�G�_P�P1H� +EH��ߟ߱�����������C�KPAU�S�Q1H�ף  IR�S�H�A��e�� ������������� E�+�i�{�a����A?Iץ�MؐNFoO 1���� �3��$4�A��Y���[���2#�@"���Nl,�*�����B����C�_��0C�+�r�|�2���Pb�O� �� ��LLECT�_�!�����E�N+`�ʒ���ND�E�#�/��1234567890�"�A��$/ҵHw��#)j� �<i{��;��/ ��/`/+/=/O/�/ s/�/�/�/�/�/�/8? ??'?�?K?]?o?�?��?�?�?O�?��$ο ��IOG &��"S�`�O�O�O�O`GTR�2'DM(��^�?�N�N�(oM Z��_�MOR)q3)H�� 7ىU3��Y�_�_�_�_ �_�[bR�kQ*H�C�?<�<Ѡ<cz�K(Fd���P,��;ϒo�o�o˿�o�o(œh�UY@E�o�S �sj]a�PDB.����4cpmidbag3��Рs:��>�uqpz��v  ���>x��}`.��}�`��|�<�CmgP���t��~f�������@ud1�:�?��XqDEFg -��zC)*��cO�buf.txAtJ��|K�[`�/DM=��>���R�A6��MCiR20_{RC�d���hS21����G���CzA�d4��EI�jC%�e�C6� G/X"DO[oF]��H�j�F� �F�TWJ��i�G�JI؂��LڒYJ4�JN�N���mKE�NMSo��������f23FDLD�	>z�!� Y2��}��yc
�@�x9� C�Ĵ�  D4G�E����  E%q��F�� E�p��u�F�P E���fF3H ?��GM��Ъ>5�>�33��?��xn9�q@�Q5�����RpA?a��=�L��<#�QU��@,�Cϒ���RS�MOFST +xi�����P_T1Ɠ�4DMA =ք�M?ODE 5dm�@c��	Q�M;���%��?���<�M>��Ͷ�/TESTc�2i�`�ER�6�O�K�CN�QAB���n� 8��\�n�CdB���C�pp�����p:;d�QS ��ՠ ������4�I7R>���>B8m5�$�RT_c�PRO/G %j%��d�|1�h@NUSER���x�KEY_TBL�  e�����	�
�� !�"#$%&'()�*+,-./(:�;<=>?@AB�Cc�GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������>���͓���������������������������������耇��������������������4A8�LCK��F�y��OSTAT��2�X��_ALM�����_AUTO_DO��E�FDR 3�:i�2h&q[~��� BUO�SYST-322� Auto st�atus che�ck time out ���i�$TELEO8|�i� ��)q�A�ʜ@Ĭ������?�ڛ�MsB�õ��?*?���?Mf=�o�TR��-����D.�B����C���B�yN�*p�4�N�4�J5Hj5H���>�i�BJ�d�B�F��pZ��[~�b bt����5/��M*F�B�G�A+$����@R��J�}�BQ�H����������2�>��@�@����&��CBxHCKH<B��6>Tbt���/��[��+���g?/$/�?��'lS�!���rA��7�A��y��x��&��BC��!@��?�1�?+*���0��0&����@ڒ�?���Ba��5�&o-�tO�tD�:O���/�/?��u�US�O�O�Oi�$ �O_:�c@m� _J_p ��N_8_�_�_V_�_�_ �_�]�Oo)o;o�OLo qo_�o�o�_�o�o�o �o�o�oFXo ��No���o�� ��@�N�$�b�x� ����n������ A��b�\�z�|�n��� ����ʟ���(�֏O� a�s������T�ʯį ��֯����2�H� ~���>���ɿۿ��� ϼ�2�,�J�L�>�x� ��\Ϛϰ����Ϧ�� 1�C��T�y�$Ϛߔ� �ϴߦ��������� N�`�߇���V߼� ���������H� V�,�j�������v��� ��$I��jd ���v����� 0��Wi{&� �\�����/ &/�:/P/�/�/F�/ �/�/��/?�:?4? R/T?F?�?�?d?�?�? �? O�/'O9OKO�/\O �O,?�O�O�?�O�O�O �O�O
_ _V_h_O�_ �_�_^O�_�_�O
oo "_$ooPo^o4oro�o �o�o~_�o	�_, Q�_rl�o�~� ����&�8��o_� q���.����dڏԏ ��� �.��B�X� ����N�ǟٟ럖��� !�̏B�<�Z�\�N��� ��l����������/� A�S���d���4����� ¯Ŀ�����Կ�(� ^�p���ϩϻ�f��� �Ϝ���*�,��X� f�<�zߐ����߆��� �#���4�Y��z�t� �ߔ����������� .�@���g�y���6�� ��l�����������( 6J`��V�� ����)��JD bdV��t�� �/�7/I/[/l/ �/<�/�/��/�/�/ ?�/?0?f?x?&/�? �?�?n/�?�?�/OO 2?4O&O`OnODO�O�O �O�O�?__+_�?<_ a_O�_|_�O�_�_�_ �_�_�_ o6oHo�Ooo �o�o>_�o�ot_�o�o o�o0>Rh ��^o����o� 1��oR�L�jl�^��� ��|���Џ���?� Q�c��t���D����� ҏԟƟ ���"�8� n���.�����˯v�ܯ ���"��:�<�.�h� v�L�����ֿ迖�� !�3�ޯD�i���τ� ���ϖ����ϴ���� >�P���w߉ߛ�FϬ� ��|�����
����8� F��Z�p���f��� ������9���Z�T� r�t�f�����������  ��GYk�| �L������� �*@v�6� ��~�	/�*/$/ BD/6/p/~/T/�/�/ �/�/�?)?;?�L? q?/�?�?�/�?�?�? �?�?�?OFOXO?O �O�ON?�O�O�?�O�O O__@_N_$_b_x_ �_�_nO�_�_o�Oo Ao�Obo\oz_|ono�o �o�o�o�o(�_O aso��To�� �o�����2�H� ~���>��ɏۏ�� ��2�,�J�L�>�x� ��\����������� 1�C��T�y�$����� ��������į�� N�`��������V��� ῌ�������H� V�,�jπ϶���v��� �߾�$�I���j�d� �τ�v߰߾ߔ����� �0���W�i�{�&ߌ� ��\������������ &���:�P�����F�� ����������:4 R�TF��d�� � ��'9K��\ �,������ ��
/ /V/h/�/ �/�/^�/�/�
?? "/$??P?^?4?r?�? �?�?~/�?	OO�/,O QO�/rOlO�?�O~O�O �O�O�O�O&_8_�?__ q_�_.O�_�_dO�_�_ �O�_�_ o.ooBoXo��otc�$CR_F�DR_CFG };re�Q?
UD1:�W�Pu�PJ�d  �`��\�bHIST 3�<rf  �` � ?�R@�tAtB�bC��PYpDtEtI�tg�Ppotw��_��bINDT_�EN6p�T��q�bT1_DO  �U�u�s�T2��wVAR �2=�gp h�q  -�Mt��t�R��4�����m[��RZ�`S�TOP��rTRL?_DELETNp�t� ��_SCRE�EN re�r_kcsc�rUw��MMENU 1>~��  <�\%�_��T��R��S /�U���e�w�ğ���� ��џ�	�B��+�x� O�a�����������ͯ ߯,���b�9�K�q� ������࿷�ɿ�� ��%�^�5�Gϔ�k�}� �ϡϳ��������H� �1�~�U�gߍ��ߝ� ��������2�	��A� z�Q�c������� ����.���d�;�M� ��q�������������YӃ_MANUA�L{��rZCD�a�?�y�rG ����R�f"
�"
?�|(��PdTGR�P 2@�y�cB� � s��~� �$DBCO�p�RIG���v�G_�ERRLOG 	A��Q�I[m� �NUMLI�M�s��u
�P�XWORK 1B�8���//��}DBTB_�� CC%���S"�� �aDB_AWA�Y��QGCP Ϋr=�ןm"_AQL�F�_�Yz�����p�vk  1D>� , 
��/0"�/%?/(_M�pq�w,@�=5ONTImM����t�_6�)
�0�'MOT�NENFpF�;RECORD 2J�� �-?�SG�O��1�?"x"!O3OEO WO�8_O�O�?�OO�O �O�O�O�O(_�OL_�O p_�_�_�_A_�_9_�_ ]_o$o6oHo�_lo�_ �o�_�o�o�o�oYo }o2�oVhz��o ��C�
��.� �R��K�������� Џ?��ߏ�*����� +�b�t�㏘�����Ο =�O�����:�%��� p�ߟ񟦯��O�ǯ� ]������H�Z��� ������#�5��������i"TOLERE�NCv$Bȿ"� L���� CSS_CCSCB 2K�	\0"?"{ϰ� ����7��
����@�@R�d�3߈ߚ�"�x� ��������'�9�K� ]�o��������� �����#�5�G�Y�k� }��������������� 1CUgy��� �����Y�R�LL]�La��m1T#2 C�C��F�^W A�C�pC���#�0� 	 3A���B���?�  �$�����\0袰�0��B��`#s�K/]/o/��
�/�/�/s/�/��/�K{�0L�e�>5�1�r��9Kr�Ȧ��/��/`?;�@��O?�?�?�?Ȏ0AF��?{F�A OO�7�1���9M	AB
AZOdBAE@�9$O�O�O�Oi:P�н`�@0�DJC^A� @��
�X-.
[#_   M?�>O�ڴ�q_�_ �_�_:W�A<o�:[<ǲ/o�/�_�+oPoboto�eACH�C�V�WB$�Dz�cD�`�a=/�o�oo��oW�a.+!��2 =t,y�J?�.s�s� js�w�yj���� ���Q�Qs�@`� �$�����A����B މ�o��'�9��_]� o�N���r���ɟ۟_��B�ʄ��YZ>`��>��A��zB��@��6>V�y��X0� Z�l�~����`_ м¯���
���̯9� ,�]�o��� �H����� ٿ뿊��ƿ3�E�W� iϬ���$ϱ����� � �����/�A�S߶�w� V�h߭ߌ��S���ߐ�_�f	��H�?� Q�~�u������� �����D��-�g� q�������������
 @7Icm�8�߾�  ��� ��)M@qd v������� //I/P�m/�v/�/ �/�/�/�/�/�/?3? *?<?i?`?r?�?^/�? �?�?�?�?O/O&O8O JO\O�O�O�O�O�O�O|�O�g	  Q��P�s ��PC4p*p�pp6U6P\C9p/p�� ]V^PM]�6P�:P�>P�VJ_+�^P�bP�fP�VLr]v���p Q
k� ��_oo�id1Q&oNo ;o_co�oˏUUA   �o�k1Q@�  �o�k�b�]�����p( �� 1��6�01C���C�cPfL��?#��c>�{��2�`�cP�@@�d�,�r�`B�cP>�s�q;C��p����b�t�<�o?�PH?�)S�B�tq0�q�p�r�`B���eDIC�&�Q�4( �o�z�UU�:��9���@���>V�^Ϲ�/Q�-R@�`���W�c��Bg�)�by��`ځ`  ?�p����U�[?����}t��$���$DC�SS_CLLB2� 2M���p�P�^?�NSTC�Y 2N��?�  ��� ����ʟ؟���� � 2�D�Z�h�z��������¯ԯ��SA�DEV�ICE 2O��!�$��4&V�h��� ����˿¿Կ���
� 7�.�[�R�ϑϣϵ������4(A�HNDG�D P��*�Cz|�A�LS 2Q��_�Q�c�u߇ߙ߫������?�PARAM RP��1�`�&տRBT 2T��/ 8�P<C�'pG �qi�l��sF@"�R��(qI�X���0�pB CW  ��B\x�N��`Z��&���%��)���X�@j��p����zq�����B �(s,�F�p��V��q���b��B ��4&c �S�e�l�4+�����H1~�����D�C�$Z|��b���A,� �4�u@�X@��^@w���]�B���B�cP%���C4�C3�:^C4��n��� ��p8�-B�{B��A����� l��C��C3�JC4jC3��yn�+�3 Dff 2�A PB W4+@:�]o�W�� ���/�/P/'/ 9/K/]/o/�/�/�/�/ ?�/�/�/?#?5?�? Y?k?�?�?�o�?�?O �?6O!OZOlOWO�O�E s�?�?�?�O�O_�O �OL_#_5_G_Y_k_}_ �_�_�_ o�_�_�_o o1o~oUogo�o�o�o �o�owO D/A ze����O�o�o 
��o��R�)�;��� _�q����������ݏ �<��%�r�I�[�m� �������ǟٟ&�8� �\�G���k������� گů�����F�� /�A�S�e�w�Ŀ���� ��ѿ�����+�x� O�aϮυϗϩϻ��� ��,���b�t�ﯘ� �߼ߧ��������� :��C�U߂�Y�k�� ����������6�� �l�C�U�g�y����� ������ ��	- ?Q������ �@+dvQ� ������� *///%/r/I/[/�/ /�/�/�/�/�/&?�/ ?\?3?E?�?i?{?�? �?U�?�?"O4OOXO CO|OgO�O{��?�O �?�O�O0___f_=_ O_a_s_�_�_�_�_�_ o�_oo'o9oKo�o oo�o�o�o�o�o�O :%^I�������H�$DCS�S_SLAVE �U���	����z_4D�  	��AR_MENU V	� �j�|�������ď��BY�� ��~?�S�HOW 2W	� � �b�aG�Q� X�v���������П֏���� @�:�d�a� s����������߯� �*�$�N�K�]�o��� ����̯ɿۿ��� 8�5�G�Y�k�}Ϗ϶� ����������"��1� C�U�g�yߠϝ߯��� �����	��-�?�Q� c��s��������� ����)�;�M�t��� �������������� %7Ip�m�� ��������! 3ZWi���J ����//DA/ S/e/��/��/�/�/ �/�/?./+?=?O?v/ p?�/�?�?�?�?�?�? ?O'O9O`?ZO�?�O �O�O�O�O�OO�O_ #_JOD_nOk_}_�_�_ �_�_�O�_�_o4_.o X_Uogoyo�o�o�o�_ �o�o�ooBo?Q cu���o:��~�CFG X)��3�3q5p��FRA:\!�L�+�%04d.CS�V|	p}� ��qA g�CHo�z@v�	����3q�����́܏� ���4��JP����q�p1� �RC_�OUT Y���C��_C_�FSI ?i� .����� ��͟�����>�9� K�]���������ίɯ ۯ���#�5�^�Y� k�}�������ſ�� ���6�1�C�U�~�y� �ϝ����������	� �-�V�Q�c�uߞߙ� �߽��������.�)� ;�M�v�q����� �������%�N�I� [�m������������� ����&!3Eni {������� FASe�� ������// +/=/f/a/s/�/�/�/ �/�/�/�/??>?9? K?]?�?�?�?�?�?�? �?�?OO#O5O^OYO kO}O�O�O�O�O�O�O �O_6_1_C_U_~_y_ �_�_�_�_�_�_o	o o-oVoQocouo�o�o �o�o�o�o�o.) ;Mvq���� �����%�N�I� [�m���������ޏُ ���&�!�3�E�n�i� {�������ß՟���� ��F�A�S�e����� ����֯ѯ����� +�=�f�a�s������� ��Ϳ�����>�9� K�]φρϓϥ����� ������#�5�^�Y� k�}ߦߡ߳������� ���6�1�C�U�~�y� ������������	� �-�V�Q�c�u����� ����������.) ;Mvq���� ��%NI [m������ ��&/!/3/E/n/i/ {/�/�/�/�/�/�/�/�3�$DCS_C�_FSO ?����71 P ??T? }?x?�?�?�?�?�?�? OOO,OUOPObOtO �O�O�O�O�O�O�O_ -_(_:_L_u_p_�_�_ �_�_�_�_o oo$o MoHoZolo�o�o�o�o �o�o�o�o% 2D mhz����� ��
��E�@�R�d� ��������ՏЏ�� ��*�<�e�`�r��� ������̟����� =�8�J�\�������?_C_RPI4>F? �������3?�&��o����� >SLү@ d������%�7�`� [�m�Ϩϣϵ����� �����8�3�E�W߀� {ߍߟ���������� ��/�X�S�e�w�� �����������0� +�=�O�x�s������� ������'P K]o����� ���(#5Gp k}�����Q�� �/6/1/C/U/~/y/ �/�/�/�/�/�/?	? ?-?V?Q?c?u?�?�? �?�?�?�?�?O.O)O ;OMOvOqO�O�O�O�O �O�O___%_N_I_ [_m_�_�_�_�_�_�_ �_�_&o!o3oEonoio {o�o�o�o�o�o�o�o FASe�������>�NOC�ODE ZU���?�PRE_CHK \U���pA �p�< ��pU�]�o�U� 	 <Q����� ���ۏ�Ǐ�#��� �Y�k�E�����{�ş ן��ß����C�U� /�y�����s���ӯm� ��	���?��+�u� ��a�������ɿ�Ϳ ߿)�;��_�q�K�}� �ϝ������ω���%� ���[�m�Gߑߣ�}� ���߳����!���E� W�1�c��g�y����� ���������A�S�-� w���c����������� ��+=asM _������ '�]o	�� ����/#/� G/Y/3/e/�/i/{/�/ �/�/�/?�/?C?9 Ky?�?%?�?�?�?�? �?	O�?-O?OOKOuO OOaO�O�O�O�O�O�O �O)_____q_K_�_ �_a?�_�_�_�_o%o �_Io[o5oGo�o�o}o �o�o�o�o�o�oE W1{�g���_ ����/�A��M� w�Q�c���������� Ϗ�+���a�s�M� ��������ߟ��� '���3�]�7�I����� �ɯۯ������� G�Y�3�}���i���ſ ��������1�C��� +�yϋ�eϯ��ϛ��� ������-�?��c�u� Oߙ߫߅ߗ������� �)��M�_�U�G�� ��A����������� ��I�[�5����k��� ����������3E Q{q���] ����/Ae wQ������ �/+//7/a/;/M/ �/�/�/�/�/��/? '??K?]?7?�?�?m? ?�?�?�?�?O�?5O GO!O3O}O�OiO�O�O �O�O�O�/�O1_C_�O g_y_S_�_�_�_�_�_ �_�_o-oo9oco=o Oo�o�o�o�o�o�o�o __M_�ok� o������� �I�#�5����k��� Ǐ��ӏ��׏�3�E� �i�{�5c���ß�� ���ӟ�/�	��e� w�Q�������ѯ㯽� ϯ�+��O�a�;��� �����Ϳ߿y��� �!�K�%�7ρϓ�m� ���ϣ���������5� G�!�k�}�W߉߳ߩ� �����ߕ��1��� g�y�S������� �����-��Q�c�=� o���s��������� ����M_9�� o����� 7I#mYk� �����!/3/) /i/{//�/�/�/�/ �/�/�/?/?	?S?e? ??q?�?u?�?�?�?�? OO�?%OOOE/W/�O �O1O�O�O�O�O__ �O9_K_%_W_�_[_m_ �_�_�_�_�_�_o5o o!oko}oWo�o�omO �o�o�o�o1U gAS����� �	����Q�c�=� ����s���Ϗ�o��� ���;�M�'�Y���]� o���˟����۟� 7��#�m��Y����� �������!�3�ͯ ?�i�C�U�������տ �������	�S�e� ?ωϛ�uϧ��ϫϽ�������$DC�S_SGN ]�	�E��-����01-DEC�-25 19:2�0 ��29-�NOVV�20:2�7_�x�x� /[}�t��q�т��xҚك�JѨ�E���Þ� ������  1�HOW �^	�� x�/�VERS�ION =�V4.5.2���EFLOGIC �1_���  	�����C��R�%��PROG_ENB  ��:�{�s�ULSE  X����%�_ACCL{IM������d��WRSTJN�T��E��-�EM�O|�zя�$���IN�IT `2�����OPT_SL �?		�	�
 	�R575��]�7�4b�6c�7c�50��1���C���@�TO  L���� �V�DEX��d�E�x�PATHw A=�A\�k}��HCP_CLNTID ?�:� D�ռ���IAG_GRP� 2e	�����z�	 @��  
ff?a�G���B�  2��/�8[I�@c�ς!�7�@�z�@^��@
�!��m�p2m15 89�01234567�����  �?��?�=q�?��
?޸R�?�Q�?���?�����(��?�z���x�@o�  A_�Ap ,!7A�88_�;B4�� ��L��x�
�@�@���\@~�R@�xQ�@q�@�j�H@c�
@�\��@U�@Mp��//'$��; �O)H��@C�t >d 9��@4��/\)@)� #�t {@���/�/�/�/�/P'?�/��?���_ �?}p�?u�?n{?s ?\�Q�? ?2?D?|V?h8�
=?��鎌0w5�z�H�?p�h��?^�R�?�?�?�?�?h8���t0���,@�?��0�;@ &O8OJO\OnOP'�$_ �_Y_k_�O?_�_�_ �_�_�_s_�_�_1oCo !ogoyoo�o��Bj"�� �2{1�@"?�Ś�f�t0�d"5!{�
u4V��u@"�B3t�A>u��?�@[q��@`,=q��=b��=��E1>�J�>��n�>��H"<w�o �z�s�q���� �x�C�@<w(�Uz� 4i�� ����A@x�?*�o��m*�P�b� ��tn���2���Ώ��x���i>J��&��bN2�"��GI�N��o@�@v���0y����@ffr9!l ��33����(��"C�� �ƒI�CH�)�C.dBت "8"����'��� "~�A?�&"K����pf�B��@�p��������p��?5���3�|Y=�y�2��/�6�B���65=���6
�*�~�`C���B���C�_�xВ������D3��N�T������0C+�r�|�2�G#�����ȿ ���׿����?,��<�o��CT_CONFIG f���|�eg�Y��STBF_TTS��
����О�t}���1�MAU�������MSW_CF���g�  # ��O�CVIEW��h!�-���s߅ߗ� �߻��ߟ�a����� ,�>�P���t���� ����]�����(�:� L�^������������ ��k� $6HZ ��~������ y 2DVh��������v�R%C�i���!��� /S/B/w/f/�/�/�/���SBL_FAULT j*6��!GPMSK���'���TDIAG k���-�������UD1: 67�89012345 I2��=1�Ǥ�P\υ? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�Od696���r
t?�O|ƟTRECP"?4:
 B44_[7��s?p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�O�O��O�o7�UMP_O/PTIO=��.�a�TR����)uP�ME��Y_TE�MP  È�+3BC�gp�B�Qt�UNI����gq�Y�N_BRK l�L�7�EDITOR��a�a@�r_
PEN�T 1m) � ,&TELE�O[p���&SET_WCp,��l>�pPSNAP^PX�>?�MTPG�pW� i��/��IĦ��ʏ� ��=�$�a�H����� ~�����ߟ�؟��� 9� �2�o�V���z��� ɯ���ԯ�#�
�G��DɴpMGDI_S�TAzuV�gq�uNC�_INFO 1n<!��b���X����������n�1o!� C��o����
�d�oU�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫���  u����
��*�B�*� P�b�t������� ������(�:�L�^� p���������2����� ��9�CUgy �������	 -?Qcu�� ������//1 ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?��? �?�?O)/OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�?�?�_�_o�_ 3O=oOoaoso�o�o�o �o�o�o�o'9 K]o����_�_ ����+o5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� �������ӟ���	� #�-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ����7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߹��������� �%�/�A�S�e�w�� ������������ +�=�O�a�s������� ���������'9 K]o����� ���#5GY k}�	����� �/1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? ��?�?�?�?/O)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�?�_�_�_ �_O�_!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �_�_����o� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o�������ɟ ۟���#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߝ��߹� ���������%�7�I� [�m��������� �����!�3�E�W�i� {��߇���������� /ASew� ������ +=Oas����� �����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?���?�?�?�?� �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�?�_ �_�_�_�?�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m�_u����_ ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�� ������u������ +�=�O�a�s������� ��ͯ߯���'�9� K�]�w���������ɿ �����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g߁� �ߝ߯���ۿ����	� �-�?�Q�c�u��� �����������)� ;�M�_�y߃������� ������%7I [m����� ��!3EWq� c��������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?i{�?�?�? �?��?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_�? s?}_�_�_�_�?�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qk_u�� ��_�����)� ;�M�_�q��������� ˏݏ���%�7�I� cQ���������ٟ ����!�3�E�W�i� {�������ïկ������/�A�[� �$�ENETMODE� 1p��_�  k�k��f�����j�OAT�CFG q�����Ѵ��C����DATA 1�rw�Ӱ���*	�*��'�9�K�]�"l�dlύ�e��� ����������'ߡ� ��]�o߁ߓߥ߷�1� ��U����#�5�G�Y� ���ߏ��������� ��u��1�C�U�g�y� �����)�������	 -����cu�����j�RPOS/T_LO��t�[�
׶#5Gi�R�ROR_PR� �%w�%L�XTA�BLE  w��ȟ����RSE�V_NUM ��?  ���  ��_AUTO_ENB  ���Xw_NO5! uw����"  *�*x �x �x �x + �+w �/�/�/Q$FLsTR=/O&HIS#�]�J+_ALM �1vw� �[x,e�+�/Q?c?u?��?�?�?�/_"W   w�v!���:j��TCP_VER �!w�!x�?$E{XT� _REQ�&s�H)BCSIZKO�=DSTKhIf%��?BTOL  �]Dz�"�A =D_BWD�0�@�&��A���CDI�A �wķ���]�KST�EP�O�Oj�POP�_DO�Oh�FDR_GRP 1xw��!d 	�?�_��yP�s�Y�Q'��M"���l���T� �����VyS�_�]�TA8���AU��@�d��_�_ okGo2o�Wo}oho�o�o�om?����@p�?��=����n
 L��z$b �`�o���3:�o^I̂hA@`�t@S33�uh}@�q�gx��yPF@ ���|yPG�  @�Fg�fC�8RL���}?��`i��~6��X����875t���5���5`�+��~��� ������� �Zk�� �����FEATU�RE y���@���Hand�lingTool� �]Eng�lish Dictionary��4D St��ar�d��Analo�g I/O>�G�g�le Shift�Z�uto Sof�tware Up�date�mat�ic Backu�p���groun?d Edit ���CameraU�F�Y�CnrRndI�m���ommon� calib U�I��nˑ�Mo�nitor$�tr~�Reliabn���DHCP �[�a�ta Acqui�s3�\�iagno�s��R�v�ispl�ayΑLicen�sZ�`�ocume�nt Viewe�?�^�ual Ch�eck Safe�ty��hanc�ed���s�F�rܐ�xt. D7IO /�fi��@�wend�Err>�QL��\�4�s[�rP��K� �@
�FCTN_ Menu��vZ����TP In��f�acĵ�GigE�־�Đp Mas_k Exc�g=��HT԰Proxy� Sv��igh�-Spe�Ski��� Ť�O�mmun�ic��onsV�u�r����q�V�ײconnect 2���ncrְstruH!��ʴ�eۡ��J���X�KAREL C�md. L�ua����Run-Ti�<�Env�Ȟ�el� +��s��S/W��ƥ���r�Boo�k(System�)
�MACROs�,M�/Offse�u�p�HO���o�u�M�R8�4���Mech/Stop+�t����"p�im�q���x�R�쪐��odo�wit#ch�ӟ�.��4�OptmF��,�f�il䬳�g��p�ulti-T�Γ�PCM fun��¼�o��������Re�gie�rq���ri�ݠF���S�Num� Sel��/�:� Adjua�*�W�q�h�tatu��ߪ��RDM Rob�ot�scove�'���ea��<�Freq Anlyq�'Rem��O�n5���>��ServoO�!�~�SNPX b-�vv�SN԰Cliܡ<?r�Libr&�_��� ��q +oJ�t��ssag��X�@a ����	�@/Iս>�MILIB��?P Firm����P��AccŐ͛T�PTXk��eln���������or�quo�imulah=��|u(�Pa&���ĐX�B�&+�ev�.���ri��T�USB port- �iPf�aݠ&?R EVNT� nexcept�`����%5��VC�rl�c���V���"h�%q�+SR SCN��/SGE�/�%UI~	�Web Pl�� >��A43��ۡ���ZDT Applxj�
�{1EOAT�౔�&0?�7Gri�d�񾡬=�?iR��".5� F���/גR�X-10iA/L��?Alarm C�ause/��ed�(�All Smo�oth5���C�sc�ii+�V�Load�䠌JUpl�@w�t�oS ��rity�AvoidM(�sb7�t�@�ycn�`����_�CS+����. c��XJo ���-T3_H�.RX���U���Xcolla3bo����RA�:�.9D��in���gNRTHI
�On��e Hel����ֿ������1trU�R?OS Eth$��A@������;,�G �B�,|HUpV�%�fW�t ԰�_iRS��ݐ�64MB D�RAM�o�cFROp���L8F FlD������2M �A:�op�m�ԕex@V�
�sh��q��wce�u��p,��|tyn�sA�
��%�r����J��^�.v� P)Q/sbS�`�p��O�N��mai���U���R�q�T�1�^FC+Ԍ%̋F�s9�ˌk̋��Ty-p߽FC%�hױV�:N Sp�ForްK��Ԭ�lu!����cp�OPG j�֡�RJ:�[L`Sup"}�0�֐f��crFP��3lu� ��al�����r��i�
q�4�@а�uest,IMPLE ׀6*�|HZ���c0�BTe�a(�|���$rtu8���V�9HMI�¤���UIFc�pono2D�BC�:�L�y� p���������ʿܿ	�  ��?�6�H�u�l�~� �Ϣϴ��������� ;�2�D�q�h�zߧߞ� ���������
�7�.� @�m�d�v����� �������3�*�<�i� `�r������������� ��/&8e\n �������� +"4aXj�� ������'// 0/]/T/f/�/�/�/�/ �/�/�/�/#??,?Y? P?b?�?�?�?�?�?�? �?�?OO(OUOLO^O �O�O�O�O�O�O�O�O __$_Q_H_Z_�_~_ �_�_�_�_�_�_oo  oMoDoVo�ozo�o�o �o�o�o�o
I @Rv���� �����E�<�N� {�r�������Տ̏ޏ ���A�8�J�w�n� ������џȟڟ��� �=�4�F�s�j�|��� ��ͯį֯����9� 0�B�o�f�x�����ɿ ��ҿ�����5�,�>� k�b�tφϘ��ϼ��� �����1�(�:�g�^� p߂ߔ��߸�������  �-�$�6�c�Z�l�~� ������������)�  �2�_�V�h�z����� ����������%. [Rdv���� ���!*WN `r������ �//&/S/J/\/n/ �/�/�/�/�/�/�/? ?"?O?F?X?j?|?�? �?�?�?�?�?OOO KOBOTOfOxO�O�O�O �O�O�O___G_>_ P_b_t_�_�_�_�_�_ �_oooCo:oLo^o po�o�o�o�o�o�o	  ?6HZl� �������� ;�2�D�V�h������� ˏԏ���
�7�.� @�R�d�������ǟ�� П�����3�*�<�N� `�������ï��̯�� ��/�&�8�J�\��� ��������ȿ����� +�"�4�F�Xυ�|ώ� �ϲ���������'�� 0�B�T߁�xߊ߷߮� ��������#��,�>� P�}�t������� ������(�:�L�y� p��������������� $6Hul~�����  H552�v�21R78{50J614�ATUP'545z'6VCAMwCRIbUIF'�28cNRE5�2VR63SC�HLIC�DO�CV�CSU8�69'02EIOuC�4R69V�ESET?UJ7�UR68MAS�KPRXY{7.OCO#(3?�+ &3j&J6%5u3�H�(LCHR&�OPLG?0�&M�HCRS&S�'MC�S>0.'552MgDSW+7u'OPu'GMPRv&��(0&7PCMzR0q7+ �2� �'51J51��80JPRS"'6�9j&FRDbFR�EQMCN9=3&SNBA��'/SHLBFM1G��82&HTC>T�MIL�TPA��TPTXcFEL�F� �8J�95�TUTv'9�5j&UEV"&UE�CR&UFRbVCuC
XO�&VIPnFwCSC�FCSG���IWEB>HTT>R6��H;�RVCGiWIGQWI�PGS�VRCnFD�Gu'H7�7R66�J5'R�8R5U1
(6�(2�(5VR�J8�86�L=Ih% �84g662wR64NVD"&�R6�'R84�g7�9�(4�S5i'J[76j&D0�gF x�RTSFCR�gC;RXv&CLIZ8I�CMS�Sp>STuYnG6)7CTO>���7�NNj&O�RS�&C &FCBn�FCF�7CH>wFCR"&FCI�VKFC�'J�PO7GBf�M�8OLaxENDvS&LU�&CPR�7ULWS�xC�STx�TE�gS60F�VR�IN�7IH aF�я�����+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi{ ������� /ASew�� �����//+/ =/O/a/s/�/�/�/�/ �/�/�/??'?9?K? ]?o?�?�?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_ �_�_�_�_�_�_	oo -o?oQocouo�o�o�o �o�o�o�o); M_q����� ����%�7�I�[� m��������Ǐُ��  H5�52��21�R�78�50�J6{14�ATUP7��5457�6�VC�AM�CRI��U�IF7�28��NR�E�52v�R63��SCH�LIC�ƚDOCV�CS]U�8697�0F��EIOCǛ4�R{69v�ESETW�vu�J7u�R68��MASK�PRXuY��7�OCO���3W����6�3�J�65�536�H$�L{CHƪOPLGW��0�MHCRǪS���MCSV�0��5=5F�MDSW���;OP��MPR��㐺6�06�PCM��R�0E˓�F���6�51�f�51��0f�PR�S��69�FRDކ�FREQ�MC�N�936�SNByAכ%�SHLB��ME��ּ26�HT=CV�TMIL�6��TPAV�TPTXF��ELړ�6�8%��#��J95��TU�T��95�UEVUECƪUFR���VCCf�O��V�IP��CSC��C�SGƚ$�I�WE�BV�HTTV�R6�՜��S���CG��I�G��IPGS'�RmC��DG��H7�˗R66f�5�u�R���R51f�6�2��5v�#�J׼��6B��LU�5�s�v�4���66F�R64�N�VD��R6��R8�4�79�4��S�5�J76�D0�uFRTS&�C�R�CRX��CL9I&�e�CMSV�s�V�STY��6�C�TOV�#�V�75�NN�ORS����6�wFCBV�FCF�˻CHV�FCR��F[CIF�FC��J#�j�G
M��OL��ENDǪLU��C�PR��Lu�S�C�$�StTE�S6�0�FVRV�IN��IH���m??�? �?�?�?�?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_e_w_�_�_�_�_�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9K]o� �������� #�5�G�Y�k�}����� ��ŏ׏�����1� C�U�g�y��������� ӟ���	��-�?�Q� c�u���������ϯ� ���)�;�M�_�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�e�w������� ������+�=�O�a� s��������������� '9K]o� ������� #5GYk}�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a��s���������͏ߏ��STD�LANG��� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ�ܰ���RBT
�OPTN������'�9� K�]�o�����������DPN	��� )�;�M�_�q������� ��������%7 I[m���� ����!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O �O�O�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o	-?Qcu �������� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ �����/�A�S�e� w���������ѿ��� ��+�=�O�a�sυ� �ϩϻ��������� '�9�K�]�o߁ߓߥ� �����������#�5� G�Y�k�}������ ��������1�C�U� g�y����������������	-?Qc��f�������99��$FEA�T_ADD ?	����  	�#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ���������DEMO y~   � L�B�T߁�xߊ߷߮� ����������G�>� P�}�t������� ������C�:�L�y� p��������������� ?6Hul~ ������ ;2Dqhz�� ���� /
/7/./ @/m/d/v/�/�/�/�/ �/�/�/?3?*?<?i? `?r?�?�?�?�?�?�? �?O/O&O8OeO\OnO �O�O�O�O�O�O�O�O +_"_4_a_X_j_�_�_ �_�_�_�_�_�_'oo 0o]oTofo�o�o�o�o �o�o�o�o#,Y Pb������ ����(�U�L�^� ����������ʏ�� ��$�Q�H�Z���~� ������Ɵ�����  �M�D�V���z����� ��¯ܯ��
��I� @�R��v��������� ؿ����E�<�N� {�rτϱϨϺ����� ���A�8�J�w�n� �߭ߤ߶�������� �=�4�F�s�j�|�� �����������9� 0�B�o�f�x������� ��������5,> kbt����� ��1(:g^ p�������  /-/$/6/c/Z/l/�/ �/�/�/�/�/�/�/)?  ?2?_?V?h?�?�?�? �?�?�?�?�?%OO.O [OROdO�O�O�O�O�O �O�O�O!__*_W_N_ `_�_�_�_�_�_�_�_ �_oo&oSoJo\o�o �o�o�o�o�o�o�o "OFX�|� �������� K�B�T���x������� ۏҏ����G�>� P�}�t�������ןΟ �����C�:�L�y� p�������ӯʯܯ	�  ��?�6�H�u�l�~� ����Ͽƿؿ���� ;�2�D�q�h�zϔϞ� ���������
�7�.� @�m�d�vߐߚ��߾� �������3�*�<�i� `�r���������� ���/�&�8�e�\�n� ���������������� +"4aXj�� ������' 0]Tf���� ����#//,/Y/ P/b/|/�/�/�/�/�/ �/�/??(?U?L?^? x?�?�?�?�?�?�?�? OO$OQOHOZOtO~O �O�O�O�O�O�O__  _M_D_V_p_z_�_�_ �_�_�_�_o
ooIo @oRolovo�o�o�o�o �o�oE<N hr������ ���A�8�J�d�n� ������яȏڏ��� �=�4�F�`�j����� ��͟ğ֟����9� 0�B�\�f�������ɯ ��ү�����5�,�>� X�b�������ſ��ο ����1�(�:�T�^� �ςϔ��ϸ�������  �-�$�6�P�Z߇�~� �߽ߴ���������)�  �2�L�V��z��� ����������%��.� H�R��v��������� ������!*DN {r������ �&@Jwn �������/ /"/</F/s/j/|/�/ �/�/�/�/�/??? 8?B?o?f?x?�?�?�? �?�?�?OOO4O>O kObOtO�O�O�O�O�O��O__0]  'XF_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o�o "4FXj|�� �������0� B�T�f�x��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰπ��������
��.�  /�)�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ���(:L ^p������ � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?V?h?z?�? �?�?�?�?�?�?
OO .O@OROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo\o no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x����� ����ҏ�����,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� ������&�8�J�\� n��������������� ��"4FXj| ������� 0BTfx�� �����//,/ >/P/b/t/�/�/�/�/ �/�/�/??(?:?L? ^?p?�?�?�?�?�?�? �? OO$O6OHOZOlO ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_ �_�_�_�_�_�_
oo .o@oRodovo�o�o�o �o�o�o�o*< N`r����� ����&�8�J�\� n���������ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T�f�x����� ����ү�����,� >�P�b�t��������� ο����(�:�L� ^�pςϔϦϸ����Ϡ�� ��$�4�8� +�N�`�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�o�o �o�o�o&8J \n������ ���"�4�F�X�j� |�������ď֏��� ��0�B�T�f�x��� ������ҟ����� ,�>�P�b�t������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��� �2�D�V�h�z� �ߞ߰���������
� �.�@�R�d�v��� �����������*� <�N�`�r��������� ������&8J \n������ ��"4FXj |������� //0/B/T/f/x/�/ �/�/�/�/�/�/?? ,?>?P?b?t?�?�?�? �?�?�?�?OO(O:O LO^OpO�O�O�O�O�O��O�O __$_6Y�$�FEAT_DEM�OIN  ;T��fP�<PNTINWDEX[[jQ�NP�ILECOMP �z����Q�iRIU�PSET�UP2 {�U��R�  N ��Q�S_AP2BC�K 1|�Y G �)7Xok%�_8o<P�P&oco9U�_ �oo�oBo�o�oxo �o1C�og�o�� ,�P����� ?��L�u����(��� Ϗ^�󏂏�)���M� ܏q������6�˟Z� ؟���%���I�[�� ������D�ٯh��� ���3�¯W��d��� ���@�տ�v�Ϛ� /�A�пe����ϛ�*� ��N���r���ߨ�=� ��a�s�ߗ�&߻��� \��߀��'��K��� o���|��4���X��� ���#���G�Y���}� �����B���f������1�Y�PP�_ }2�P*.VR8���*�������l PC���FR6:�2�V�TzPz��w�]PG���*#.Fo/��	��:,�^/�STM@i/�/ /�-M/�/�H�/?�'?�/8�/g?�GIFq?�?��%�?D?V?�?�JPG�?O�%O�?�?oOF�
JSyO�O��5C��OMO%
Java?Script�O�?�CS�O&_�&_�O �%Cascad�ing Styl�e Sheets�R_��
ARGNA�ME.DT�_��� \�_S_�A�T�_�_}�PDISP*�_���To�_�QLaZo�oCLLB.Z�Iwo2o$ :\�a\��o�i�AColl�abo�o�o
TP�EINS.XML��_:\![o�QC�ustom To�olbarbiPASSWORDQo~��FRS:\��dB`Passwo�rd Config���/��(�e� �������N��r�� ���=�̏a������ &���J���񟀟��� 9�K�ڟo�������4� ɯX��|���#���G� ֯@�}����0�ſ׿ f������1���U�� y��ϯ�>���b��� 	ߘ�-߼�Q�c��χ� ߽߫�L���p��� ��;���_���X��$� ��H�����~����7� I���m���� �2��� V���z���!��E�� i{
�.��d ����S�w p�<�`�/ �+/�O/a/��// �/8/J/�/n/?�/�/ 9?�/]?�/�?�?"?�? F?�?�?|?O�?5O�? �?kO�?�OO�O�OTO �OxO__�OC_�Og_ y__�_,_�_P_b_�_ �_o�_oQo�_uoo �o�o:o�o^o�o�o )�oM�o�o�� 6��l��%�7� �[����� ���D� ُh�z����3�,� i��������ßR���v������$FI�LE_DGBCK� 1|������ <� �)
SUMM?ARY.DG!�͜OMD:U���ِ�Diag Su�mmary����
CONSLOG���n���ٯ���Co�nsole lo�g���	TPACCN�t�%\������TP Acco�untin;����FR6:IPKD?MP.ZIPͿј�
�ϥ���Exc?eption"�ӻ���MEMCHEC�K��������-�M�emory Da�ta����:n =)��RIPE�~ϸ��%ߴ�%�� �Packet L<:���L�$�c���STAT��߭�� %A�St�atus��^�	F�TP����	���/�mment T�BD2�^� >I)�ETHERNE�w�
�d�u�﨡E�thernJ�1�figuraAϩ��?DCSVRF&����7����� ve�rify all�:��� 44��DIFF/��'���;�Q�diff��r�d�>��CHG01�������A����it�2���270���f�x3���I� �p�VT�RNDIAG.LASu&8����O Ope��L� ���nostic��Y��)VDEV�DAT�������Vis�De�vice�+IM�G��,/>/�/:��i$Imagu/+�UP ES/�/�FRS:\?Z=���Updates� ListZ?���� FLEXEVEAN��/�/�?���1 UIF EvM��M���-vZ)�CRSENSPK�/˞�\!O����CR_TAOR_P�EAKbOͩPSRBWLD.CM�O�͜E2�O\?.�PS�_ROBOWEL<S���:GIG��@_��?d_��GigE��(O��N�@�)}UQHADOW__�D_V_�_��Sha�dow Chansge����5dt�R?RCMERR�_�_��_oo��4`CFG� Erroro t�ailo MA��k�CMSGLIBgoNo`o�o|R�e���z0ic�o�a�)�`ZD0_O�osn��ZD�Pad��l �RNOTI��Rd���Notific����,�AG��P�ӟt� ��������Ώ]��� ��(���L�^�폂�� ����G�ܟk� ���� 6�şZ��~������ C�د�y����2�D� ӯh��������¿Q� �u�
�ϫ�@�Ͽd� v�Ϛ�)Ͼ���_��� ��ߧ�%�N���r�� �ߨ�7���[����� &��J�\��߀��� 3����i����"�4� ��X���|������A� ����w���0��= f�����O� s�>�bt �'�K��� /�:/L/�p/��/ �/5/�/Y/�/ ?�/$? �/H?�/U?~??�?1? �?�?g?�?�? O2O�? VO�?zO�OO�O?O�O cO�O
_�O._�OR_d_ �O�__�_�_M_�_q_ oo�_<o�_`o�_mo �o%o�oIo�o�oo �o8J�on�o�� 3�W�{�"�� F��j�|����/�ď�֏e������0��$�FILE_FRS�PRT  ��������?�MDONLY� 1|S�� �
 �)MD:�_VDAEXTP.ZZZ1�⏹�ț�6%NO �Back fil�e ���S�6P �����>��K�t��� ��'���ί]�򯁯� (���L�ۯp������ 5�ʿY�׿ Ϗ�$ϳ� H�Z��~�Ϣϴ�C� ��g���ߝ�2���V� ��cߌ�߰�?����� u�
��.�@���d�������C�VISBC�Kq�[���*.V�D����S�FR:�\��ION\DA�TA\��v�S��Vision VD���Y�k���� y��B�����x��� 1C��g���, �P����? �Pu�(�� ^��/��M/� q/�/>/�/6/�/Z/�/ ?�/%?�/I?[?�/?�?�?2?D?�?9�LU�I_CONFIG7 }S����;� $ �3v�{ S�;OMO_OqO�O�O�I#@|x�?�O�O�O_ _%\�OH_Z_l_~_�_ '_�_�_�_�_�_o�_ 2oDoVohozo�o#o�o �o�o�o�o
�o.@ Rdv���� ����*�<�N�`� r��������̏ޏ�� ���&�8�J�\�n��� �����ȟڟ쟃��� "�4�F�X�j������ ��į֯����0� B�T�f����������� ҿ�{���,�>�P� b����ϘϪϼ����� w���(�:�L�^��� �ߔߦ߸�����s� � �$�6�H���Y�~�� �����]������ � 2�D���h�z������� ��Y�����
.@ ��dv����U ��*<�` r����Q�� //&/8/�\/n/�/ �/�/;/�/�/�/�/? "?�/F?X?j?|?�?�? 7?�?�?�?�?OO�? BOTOfOxO�O�O3O�O �O�O�O__�O>_P_ b_t_�_�_/_�_�_�_ �_oo�_:oLo^opo��o�o$h  x��o�c�$FLUI�_DATA ~�����a�(a�dRESU_LT 3�ep� �T�/�wizard/g�uided/st�eps/Expert�o=Oas���������z��Continu�e with Gpance�:�L� ^�p���������ʏ܏,� � �b-�a�e>�0 �0`���c�a?��ps ���������ҟ��� ��,�>�P��0ow� ��������ѯ���� �+�=�O�a�?�1�C�zU�e�cllbs� ֿ�����0�B�T� f�xϊϜ�[������� ����,�>�P�b�t� �ߘߪ�i�{��ߟ�]�e�rip(pſ-� ?�Q�c�u����� ��������)�;�M� _�q����������������������`��e�#pTimeUS/DST	��� ����!3E~�Enabl(� y��������	//-/?/Q/�b��)�/M_q24 |�/�/??)?;?M? _?q?�?�?Tf�?�? �?OO%O7OIO[OmO O�O�Ob/t/�/�/Z��"qRegion �O5_G_Y_k_}_�_�_�_�_�_�_�America!�#o5o GoYoko}o�o�o�o�o�o�o��Ay�O�O3��O_qEditor�o����������+�=� � T�ouch Pan�el rs (re�commenp�) K�������Ə؏��� � �2�D�|�%���I[qaccesoܟ� ��$�6��H�Z�l�~�����C�onnect t�o Network��֯�����0��B�T�f�x�����x�B�@��}����,!���s Introduct!_4�F�X�j�|� �Ϡϲ��������� �0�B�T�f�xߊߜ�`����������  ɿ��"�i�{�� ������������� /�A� �e�w������� ��������+="�H�3��+� O�����  2DVhz�K�� ����
//./@/ R/d/v/�/�/Yk} �/�??*?<?N?`? r?�?�?�?�?�?�?� �?O&O8OJO\OnO�O �O�O�O�O�O�O�/_ �/1_�/X_j_|_�_�_ �_�_�_�_�_oo0o BoS_foxo�o�o�o�o �o�o�o,>�O _!_�E_���� ���(�:�L�^�p� ����So��ʏ܏� � �$�6�H�Z�l�~��� O��s՟���� � 2�D�V�h�z������� ¯ԯ毥�
��.�@� R�d�v���������п ⿡��ş'�9���`� rτϖϨϺ������� ��&�8���\�n߀� �ߤ߶���������� "�4��=��a��M� ������������0� B�T�f�x���I߮��� ������,>P bt�E��i�� ��(:L^p �������� / /$/6/H/Z/l/~/�/ �/�/�/�/���� /?�V?h?z?�?�?�? �?�?�?�?
OO.O� ROdOvO�O�O�O�O�O �O�O__*_<_�/? ?�_C?�_�_�_�_�_ oo&o8oJo\ono�o ?O�o�o�o�o�o�o "4FXj|�M_ __q_��_���0� B�T�f�x��������� ҏ�o���,�>�P� b�t���������Ο�� ���%��L�^�p� ��������ʯܯ� � �$�6�G�Z�l�~��� ����ƿؿ���� � 2��S��w�9��ϰ� ��������
��.�@� R�d�v߈�G��߾��� ������*�<�N�`� r��Cϥ�g���ύ� ��&�8�J�\�n��� �������������� "4FXj|�� ��������- ��Tfx���� ���//,/��P/ b/t/�/�/�/�/�/�/ �/??(?�1U? ?A�?�?�?�?�? O O$O6OHOZOlO~O=/ �O�O�O�O�O�O_ _ 2_D_V_h_z_9?�?]? �_�_�?�_
oo.o@o Rodovo�o�o�o�o�o �O�o*<N` r������_�_ �_�_#��_J�\�n��� ������ȏڏ���� "��oF�X�j�|����� ��ğ֟�����0� ���u�7������� ү�����,�>�P� b�t�3�������ο� ���(�:�L�^�p� ��A�S�e��ω��� � �$�6�H�Z�l�~ߐ� �ߴ��߅������ � 2�D�V�h�z���� �����������@� R�d�v����������� ����*;�N` r������� &��G	�k-� �������/ "/4/F/X/j/|/;�/ �/�/�/�/�/??0? B?T?f?x?7�?[�? �?�?OO,O>OPO bOtO�O�O�O�O�O�/ �O__(_:_L_^_p_ �_�_�_�_�_�?�_�? o!o�OHoZolo~o�o �o�o�o�o�o�o  �ODVhz��� ����
���_%o �_I�s�5o������Џ ����*�<�N�`� r�1������̟ޟ� ��&�8�J�\�n�-� w�Q���ů������ "�4�F�X�j�|����� ��Ŀ�������0� B�T�f�xϊϜϮ��� ��������ٯ>�P� b�t߆ߘߪ߼����� ����տ:�L�^�p� ����������� � �$������i�+ߐ� ������������  2DVh'��� ����
.@ Rdv5�G�Y��}� ��//*/</N/`/ r/�/�/�/�/y�/�/ ??&?8?J?\?n?�? �?�?�?�?��?�O �4OFOXOjO|O�O�O �O�O�O�O�O__/O B_T_f_x_�_�_�_�_ �_�_�_oo�?;o�? _o!O�o�o�o�o�o�o �o(:L^p /_������ � �$�6�H�Z�l�+o�� Oo��sou����� � 2�D�V�h�z������� ����
��.�@� R�d�v���������}� ߯����ٟ<�N�`� r���������̿޿� ��ӟ8�J�\�nπ� �Ϥ϶���������� ϯ��=�g�)��ߠ� ������������0� B�T�f�%ϊ����� ��������,�>�P� b�!�k�Eߏ���{��� ��(:L^p ����w���  $6HZl~� ��s�������/�� 2/D/V/h/z/�/�/�/ �/�/�/�/
?�.?@? R?d?v?�?�?�?�?�? �?�?OO���]O /�O�O�O�O�O�O�O __&_8_J_\_?�_ �_�_�_�_�_�_�_o "o4oFoXojo)O;OMO �oqO�o�o�o0 BTfx���m_ �����,�>�P� b�t���������{oݏ �o��o(�:�L�^�p� ��������ʟܟ� � �#�6�H�Z�l�~��� ����Ưد����͏ /��S��z������� ¿Կ���
��.�@� R�d�#��ϚϬϾ��� ������*�<�N�`� ���C���g�i����� ��&�8�J�\�n�� ����u�������� "�4�F�X�j�|����� ��q�������	��0 BTfx���� �����,>P bt������ �/����1/[/ �/�/�/�/�/�/�/ ? ?$?6?H?Z?~?�? �?�?�?�?�?�?O O 2ODOVO/_/9/�O�O o/�O�O�O
__._@_ R_d_v_�_�_�_k?�_ �_�_oo*o<oNo`o ro�o�o�ogOyO�O�O �o�O&8J\n� ��������_ "�4�F�X�j�|����� ��ď֏�����o�o �oQ�x��������� ҟ�����,�>�P� �t���������ί� ���(�:�L�^�� /�A���e�ʿܿ� � �$�6�H�Z�l�~ϐ� ��a���������� � 2�D�V�h�zߌߞ߰� o��ߓ��߷��.�@� R�d�v������� ������*�<�N�`� r��������������� ��#��G	�n� ������� "4FX�|�� �����//0/ B/T/u/7�/[]/ �/�/�/??,?>?P? b?t?�?�?�?i�?�? �?OO(O:OLO^OpO �O�O�Oe/�O�/�O�O �?$_6_H_Z_l_~_�_ �_�_�_�_�_�_�? o 2oDoVohozo�o�o�o �o�o�o�o�O_�O% O_v����� ����*�<�N�o r���������̏ޏ�� ��&�8�J�	S- w���cȟڟ���� "�4�F�X�j�|����� _�į֯�����0� B�T�f�x�����[�m� ���󿵟�,�>�P� b�tφϘϪϼ����� �ϱ��(�:�L�^�p� �ߔߦ߸������� � ��ѿ�E��l�~�� ������������ � 2�D��h�z������� ��������
.@ R�#�5�Y�� ��*<N` r��U����� //&/8/J/\/n/�/ �/�/c�/��/�? "?4?F?X?j?|?�?�? �?�?�?�?�??O0O BOTOfOxO�O�O�O�O �O�O�O�/_�/;_�/ b_t_�_�_�_�_�_�_ �_oo(o:oLoOpo �o�o�o�o�o�o�o  $6H_i+_� O_Q����� � 2�D�V�h�z�����]o ԏ���
��.�@� R�d�v�����Y��} ߟ񟵏�*�<�N�`� r���������̯ޯ� ���&�8�J�\�n��� ������ȿڿ쿫��� ϟ�C��j�|ώϠ� ������������0� B��f�xߊߜ߮��� ��������,�>��� G�!�k��Wϼ����� ����(�:�L�^�p� ����S߸�������  $6HZl~� O�a�s�����  2DVhz��� �����
//./@/ R/d/v/�/�/�/�/�/ �/�/���9?�`? r?�?�?�?�?�?�?�? OO&O8O�\OnO�O �O�O�O�O�O�O�O_ "_4_F_??)?�_M? �_�_�_�_�_oo0o BoTofoxo�oIO�o�o �o�o�o,>P bt��W_�{_� �_��(�:�L�^�p� ��������ʏ܏�� �$�6�H�Z�l�~��� ����Ɵ؟꟩�� /��V�h�z������� ¯ԯ���
��.�@� ��d�v���������п �����*�<���]� ���C�EϺ������� ��&�8�J�\�n߀� ��Q������������ "�4�F�X�j�|��M� ��q��������0� B�T�f�x��������� ������,>P bt������ ������7��^p ������� / /$/6/��Z/l/~/�/ �/�/�/�/�/�/? ? 2?�;_?�?K�? �?�?�?�?
OO.O@O ROdOvO�OG/�O�O�O �O�O__*_<_N_`_ r_�_C?U?g?y?�_�? oo&o8oJo\ono�o �o�o�o�o�o�O�o "4FXj|�� �����_�_�_-� �_T�f�x��������� ҏ�����,��oP� b�t���������Ο�� ���(�:���� �A�����ʯܯ� � �$�6�H�Z�l�~�=� ����ƿؿ���� � 2�D�V�h�zό�K��� o��ϓ���
��.�@� R�d�v߈ߚ߬߾��� ������*�<�N�`� r���������� ����#���J�\�n��� �������������� "4��Xj|�� �����0 ��Q�u7�9�� ���//,/>/P/ b/t/�/E�/�/�/�/ �/??(?:?L?^?p? �?A�?e�?�?�/ O O$O6OHOZOlO~O�O �O�O�O�O�/�O_ _ 2_D_V_h_z_�_�_�_ �_�_�?�?�?o+o�? Rodovo�o�o�o�o�o �o�o*�ON` r������� ��&��_/o	oS�}� ?o����ȏڏ���� "�4�F�X�j�|�;�� ��ğ֟�����0� B�T�f�x�7�I�[�m� ϯ������,�>�P� b�t���������ο�� ���(�:�L�^�p� �ϔϦϸ����ϛ��� ��!��H�Z�l�~ߐ� �ߴ���������� � ߿D�V�h�z���� ��������
��.��� ���s�5ߚ������� ����*<N` r1������ &8J\n� ?��c������/ "/4/F/X/j/|/�/�/ �/�/�/��/??0? B?T?f?x?�?�?�?�? �?��?�O�>OPO bOtO�O�O�O�O�O�O �O__(_�/L_^_p_ �_�_�_�_�_�_�_ o o$o�?EoOio+O-o �o�o�o�o�o�o  2DVhz9_�� ����
��.�@� R�d�v�5o��Yo��͏ ����*�<�N�`� r���������̟�� ��&�8�J�\�n��� ������ȯ��я���� ��F�X�j�|����� ��Ŀֿ�����ݟ B�T�f�xϊϜϮ��� ��������ٯ#��� G�q�3��ߪ߼����� ����(�:�L�^�p� /ϔ��������� � �$�6�H�Z�l�+�=� O�a���������  2DVhz��� �����
.@ Rdv����� ������/��</N/`/ r/�/�/�/�/�/�/�/ ??�8?J?\?n?�? �?�?�?�?�?�?�?O "O��/gO)/�O�O �O�O�O�O�O__0_ B_T_f_%?w_�_�_�_ �_�_�_oo,o>oPo boto3O�oWO�o{O�o �o(:L^p ������o� � �$�6�H�Z�l�~��� ����Ə�o珩o��o 2�D�V�h�z������� ԟ���
���@� R�d�v���������Я �����׏9���]� �!�������̿޿� ��&�8�J�\�n�-� �Ϥ϶���������� "�4�F�X�j�)���M� ���߅�������0� B�T�f�x������ �������,�>�P� b�t���������{��� ������:L^p �������  ��6HZl~� ������/�� ��;/e/'�/�/�/ �/�/�/�/
??.?@? R?d?#�?�?�?�?�? �?�?OO*O<ONO`O /1/C/U/�Oy/�O�O __&_8_J_\_n_�_ �_�_�_u?�_�_�_o "o4oFoXojo|o�o�o �o�o�O�O�O	�O0 BTfx���� �����_,�>�P� b�t���������Ώ�� ����o�o�o[� ��������ʟܟ� � �$�6�H�Z��k��� ����Ưد���� � 2�D�V�h�'���K��� o�Կ���
��.�@� R�d�vψϚϬϾ�Ͽ ������*�<�N�`� r߄ߖߨߺ�y��ߝ� ����&�8�J�\�n�� ������������� ��4�F�X�j�|����� ������������- ��Q����� ���,>P b!������� �//(/:/L/^/ /A�/�/y�/�/ ? ?$?6?H?Z?l?~?�? �?�?s�?�?�?O O 2ODOVOhOzO�O�O�O o/�/�/�O_�/._@_ R_d_v_�_�_�_�_�_ �_�_o�?*o<oNo`o ro�o�o�o�o�o�o�o �O_�O/Y_� �������� "�4�F�X�o|����� ��ď֏�����0� B�T�%7I��m ҟ�����,�>�P� b�t�������i�ί� ���(�:�L�^�p� ��������w������� ��$�6�H�Z�l�~ϐ� �ϴ��������ϻ� � 2�D�V�h�zߌߞ߰� ��������
�ɿۿ� O��v������� ������*�<�N�� _��������������� &8J\�} ?�c����� "4FXj|�� �����//0/ B/T/f/x/�/�/�/m �/��/�?,?>?P? b?t?�?�?�?�?�?�? �?O�(O:OLO^OpO �O�O�O�O�O�O�O _ �/!_�/E_?	_~_�_ �_�_�_�_�_�_o o 2oDoVoOzo�o�o�o �o�o�o�o
.@ R_s5_��mo� ����*�<�N�`� r�������gȍޏ�� ��&�8�J�\�n��� ����c��џ��� "�4�F�X�j�|����� ��į֯������0� B�T�f�x��������� ҿ�������ٟ#�M� �tφϘϪϼ����� ����(�:�L��p� �ߔߦ߸������� � �$�6�H���+�=� ��a���������� � 2�D�V�h�z�����]� ��������
.@ Rdv���k�}�������$FMR�2_GRP 1���� ��C4  B�.��	 ��9K^6F@ a@��6G�  �Fg?�fC�8R�y�?�  ��66��X���875�t��5���5�`+�yA�  �/+BH�w-%@'S339%�5[/l-6@6!�/xl/�/ �/�/�/?�/&??J?�5?G?�?k?�?��_�CFG �T�K�?�? OO�9NO� 
F0�FA K@�<RM_C�HKTYP  ���$&� RO=Ma@_MINg@��W���@�R X�SSB�3�� 7�O���C�O�O�5TP_D�EF_OW  ��$WIRCO�Mf@_�$GENOVRD_DO�F���E]TH��D �dbUdKT_ENB�7_ KPRAVC���G�@ �@Y�O�_�?oyo�&oI* �QOU*�NAIRI<�@��oGo��o�o�o��C�p3@��O:��B��+sL�i�O�PSM�T��Y(�@
t��$HOSTC�219��@�5� MC��R{����  27.�00�1�  e �]�o�������K�ď�֏��������	a�nonymous@!�O�a�s����� �4��������D� !�3�E�W�i������� ��ï柀�.���/� A�S���课�П��� �Ŀ����+�r�O� a�sυϗϺ����� ����'�n������� �ϓ�ڿ���������� F�#�5�G�Y�k���� �����������B�T� f�C�z�g��ߋ����� �������	-P� ����u����� �(�:�<)p�M_ q�������� /$ZlI/[/m// �/����//�/D !?3?E?W?/?�?�? �?�?�/�?./OO/O AOSO�/�/�/�/�?�O ?�O�O__+_r?O_ a_s_�_�_�O�?O�_��_oo'o�t�qEN�T 1�hk P�!�_no  �p \o�o�o�o�o�o�o �o�o:_"�F �j�����%� �I��m�0���T�f� Ǐ��돮��ҏ3��� ,�i�X���P���t�՟ ��៼�
�/��S�� w�:���^���������ฯ�ܯ=� �QU�ICC0J�&�!�192.168.O1.10c�X�1��v�8��\�2�ƿؿ�9�!ROUTER:��!��a��?PCJOG��e�_!* ��0��~U�CAMPRT��ƶ�!�����RT�S���x� !S�oftware �Operator? PanelU߇����7kNAME �!Kj!ROBO�����S_CFG �1�Ki ��Auto-s�tarted�DFTP�Oa�O�_ ���O����������E_ �.�@�R�u�c�	��� ��������cN:�L�^� ;r���R���� ����%H� [m���jO|O �O�O4!/hE/W/i/ {/�/T�/�/�/�/�/ /�//?A?S?e?w?�? ����??�?</O +O=OOO?sO�O�O�O �O�?`O�O__'_9_ K_�?�?�?�?�O�_�? �_�_�_o#o�OGoYo ko}o�o�_4o�o�o�o �of_x_�_g�o ��_�����o� �-�?�Q�tu���� ����Ϗ�(:L^ `�2��q��������� ��ݟ���%�H�ʟ [�m�����������  �ί4�!�h�E�W�i� {���T���ÿտ�
� Ϟ�/�A�S�e�w�����_ERR ���ڇϗ�PDUSI�Z  �^6�����>��WRD �?(����  �guest ���+�=�O�a����SCD_GROUoP 3�(� ,��"�IFT��$P�A��OMP��� ��_SH��ED��� $C��COM���TTP_AUT�H 1��� <�!iPenda�nm�x�#�+!K?AREL:*x����KC�������VISION SET��(����?�-�W�R���v������������������G�C�TRL ����a�
��F�FF9E3���FRS:DEFA�ULT�FA�NUC Web ?Server�
t dG����/� �2DV��WR_C�ONFIG �.��������IDL_CPU_kPC� �B����� BH�MIN�����GNR_I�O������ȰHM�I_EDIT =���
 ($/C/ ��2/k/V/�/z/�/�/ �/�/�/?�/1??U? @?y?d?�?�?./�?�? �?�?OO?OQO<OuO `O�O�O�O�O�O�O�O�__;_�NPT_�SIM_DO��*NSTAL_S7CRN� �\UQ�TPMODNTOqL�Wl[�RTYbXp�qV�K�ENB�W��ӭOLNK 1�����o%o7o�Io[omoo�RMAS�TE��Y%OSLAVE �����eRAMCACH�E�o�ROM�O_CcFG�o�S�cUO'���bCMT_OPp�  "��5sYCL�o�u� _ASG 19����
 �o� ������"�4��F�X�j�|����kwrN�UM����
�bI�P�o�gRTRY_�CN@uQ_UP)D��a��� �bp�b��n��M��а�P}T?��k ��._������ɟ۟� �S���)�;�M�_�q�  �������˯ݯ�~� �%�7�I�[�m���� ����ǿٿ�����!� 3�E�W�i�{�
ϟϱ� �������ψϚ�/�A� S�e�w߉�߭߿��� ������+�=�O�a� s���&�������� ����9�K�]�o��� ��"����������� ����GYk}�� 0����� CUgy��,> ���	//-/�Q/ c/u/�/�/�/:/�/�/ �/??)?�/�/_?q? �?�?�?�?H?�?�?O O%O7O�?[OmOO�O �O�ODOVO�O�O_!_ 3_E_�Oi_{_�_�_�_ �_R_�_�_oo/oAo �_�_wo�o�o�o�o�o `o�o+=O�o s�����\n ��'�9�K�]�����������ɏۏi�c�_�MEMBERS �2�:� �  $:� ����v���1���R�CA_ACC 2��� �  [����"�� !G� �� 6�l��5l�l��&[�� ������ � il���a�BUF�001 2�n�=� ��u0u0�  ��u0X��h��u0<0�9 ��u0jh�
ȼu0'�oM����**�U8*�H*�V*�e*�Us*��*��*��*�U�*��*��*��*���������(ꚤ7��J��Yu0�p���gu0�(�L��tu0�ahȽa���ꚤ�������u0�.PF���u�0��u0_p���ݚ��u0	�`kн��0u� �����2� �2�,2�9�4�F2�R�2�`2�l2�x2���2��2�q�4��2���2��F�  F�K�r���i��q����u0�e@���
���u0�8U�ߙ2���8{��I�+���P
� �*K (�:�L�^�p������������ѡ8L�ءc��p��-�G���a�h��@i�(�p 0��p88�J�\��n��Y���t� x������ҙ���x���ҩ�F� 0���¿xe�ع!�S�ߙ3����l�� ����l� �.�2� .�:�.�Z�G�.�R�.� Z�.�b�.�j�.�r�.� ���.��.��.�� .��l��������� ����������ɠ��Ѡ ��٠��s��������� �������	������ ���!���)�l�0��� Bҗ�Jҗ�Rҗ�K�a� ��jҗ�rҗ�q���y� �Ё��Љ���>򙲧� >��������{� ȱ�Ѱ�ٲ����~d�CFG 2�n�� 4l��
l�Jl�<l�47���HIS钜n� ��� 2025�-12-�l� 64������h   7 _p  �xl�y;s�14 �l�z7 ��9 ��ՠ
����� � 3 	 U��� $� =[~�q�q1-3� �  # &f?  ' "����  P
X
`L
�   ��  C} �  8 ��@�	��}! , )�!  89�  �d�q4[}�RM29}	�R/d/v/��/�/�/�/�-) �% 9  -�R  *gl��,B��=/*?<? N?`?r?�?�?�?�?�? ??OO&O8OJO\O nO�O�O�O�?�?�O�O �O_"_4_F_X_j_|_ �O�O�_�_�_�_�_o o0oBoTo�O��[m
7d_o�o�o�o�� _� %g>�� "��"	�b  3"!�b�)"1"9:�a>A*  FI[8 cm8��� ���c��b��b� _+  X�  � UX|c	,: J|"0  Q!_1 
 RNx: 	b(aq`%/7/m�� ������Ǐُ��(5��c12Zt,�� 1� \�_�_I�[�m�� ������ǟٟ럑_4� !�3�E�W�i�{����� ��ï���Я��/� A�S�e�w�����ү� �������+�=�O� a�s�aoN�Ѐo�o
�3��������r:$qpBq� Dq�!Hq.pN�Iq>pJq!f�Npf�Vpf�:�V�� iqn[	
qm!����ߧ ���p�ҽ��p��p?�G�O� 2_�g��'J�Vp.�Z� ��J�\��� �������������*x��6�� �澿п r��������������� K�]�J\n� ������#5 "4FXj|�� ����//0/�B/T/f/x/�/�/��_�I_CFG 2���� H
Cy�cle Time��Busy��Idl�"�mi�n�+1Up|�&�Read�'Dow8?bp� 1�#Count>�	Num �"�����<p>�qaP�ROG�"�������)/sof�tpart/ge�nlink?cu�rrent=me�nupage,1133,�gOO&O�8O<b5leSDT_�ISOLC  ����p�/J23_DSP_EN>��vK0�@INC ���Ms�@A  � ?&p=���<�#�
�A�I:�o&��N_t�O<_�GOB�0C�C"�1�F�VQG_GROUP� 1�vKIr<���Cy�_D_?"x�?�_pQ�_o .o@o�_dovo�o�ow�,_NYG_IN_�AUTO �MPO�SRE^_pVKANJI_MASK v��HqRELMONG ��˔?Uby_o x�����.6r�3%��7�CUd�u�o��DKCL_L�`N�UM(��EYLO�GGING �����Q�E�0LANGU�AGE ���~��DEFA�ULT ����LGf�!��:2�?�M�80VЬU`�'��  � 
��Ua�U`GOUF ;���
��(UT#1:%�� � �-� ?�Q�h�u���������ϟ���Ub(g4�8�i�N_DISP ���O8�_�_��L�OCTOL��UaD�z<�A�A��GBO_OK ���d�1
�
�۠����� �#�5�G�Y�i���3{�W�	��쉞QQJ�¿Կ1��_BU�FF 2�vK 	�U`25
�ڢVB�&�7 Coll�aborativ �=�OΗώϠϲ��� ������'��0�]�T��fߓߊߜ��DCS ��9�B�Ax����Rh�%�-�?�Q���I�O 2��� ���Q���� ����������*�<� N�b�r����������������&:e�E_R_ITMsNd�o ������� #5GYk}����������hS�EV�`�MdTYPsN�c/u/�/
-��aRST5���SC�RN_FL 2�
s��0����/??`1?C?U?g?�/TPK��sOR"��NGNA�M�D��~�N�UPS�_ACR� �4D�IGI�8+)U_�LOAD[PG �%�:%T_NO�VICEt?��MA?XUALRM2��a����E
ZB�1_�P�5�` ��y�Z@CY��˭�O+���ۡ��D|PP 2�˫ �Uf	R/_
_C_ ._g_y_\_�_�_�_�_ �_�_�_oo?oQo4o uo`o�o|o�o�o�o�o �o)M8qT f������� %��I�,�>��j��� ��Ǐُ�����!�� �W�B�{�f������� ՟����ܟ�/��S� >�w���l�����ѯ�� Ư��+��O�a�D����p���RHDBGDEF ��E�ѱO���_LDXDIS�A�0�;c�MEMO�_AP�0E ?�;
 ױ��3� E�W�i�{ύϟϱ�Z@�FRQ_CFG k��G۳A ���@��Ô�<��d%��� ������B��K{��*i�=/k� **:tҔ� g�y�ߔ��߱����� �����J�Es��J d�����,( H���[�����@�'� Q�v�]����������������*NPJI�SC 1��9Z� ������ܿ������	Zl_MST�R �#-,SC/D 1�"͠{ �������� //A/,/e/P/�/t/ �/�/�/�/�/?�/+? ?O?:?L?�?p?�?�? �?�?�?�?O'OOKO 6OoOZO�O~O�O�O�O �O�O_�O5_ _Y_D_ i_�_z_�_�_�_�_�_ �_o
ooUo@oyodo �o�o�o�o�o�o�o�?*cN�M�K���;љ$�MLTARM��u�N��r ���հ��İMETP�U��zr��CN�DSP_ADCO�L%�ٰ0�CMNT6F� 9�FNb�f�>7�FSTLI��x�4 �;ڎ�s�����9�POSCFz��q�PRPMe���STD�1�;; 4�#�
v��q v�����r�������� ̟ޟ ���V�8�J� ��n���¯��������9�SING_CH�K  ��$MODA���t�{�~~2�DEV 	��	MC:f�HS�IZE��zp�2�T�ASK %�%�$1234567�89 ӿ�0�TR�IG 1�; lĵ�2ϻ�!�bϻ�F��YP����H�1��EM_INF 1��N�`)AT&FV0E0g����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ��2��H6�^���R����A�߶�q�������� ��5������ ߏ�B߳�������� ���1�C�*�g��,� ��P�b�t������ R�?���u0�� ������������� M q���Z� ��/�%/��[/  2�/�/h�// �/�/�3?�/W?>?{? �?@/�?d/v/�/�/O �//OAOx?eO?�ODO��O�O�O�O_�NIT�ORÀG ?z� �  	EXESC1~s&R2,X3,XE4,X5,X��.V7,X8,X9~s'R�2�T +R�T7R�TCR�TOR�T [R�TgR�TsR�TR�TT�R�S2�X2�X2�XU2�X2�X2�X2�XU2�X2�X2h3�X�3�X37R2�R_G�RP_SV 1��� (�>�����F���=5�[����濢ca���_�D�B���cION_�DB<��@�zq W �zpzp Y�21uǱ�>w�Zpzpi���@N=po�p�p>{��p5q�r-ud1������8�PG_JOG S�ʏ�{
�2��:�o�=���?����0� B��~\�n������`��H�?��C�@�ŏ�׏���  Nt��qL_NAME �!ĵ8��!�Default �Personal�ity (fro�m FD)=q1�R�MK_ENONL�Y�_�R2�a 1��L�XLy�8�gpl d�� ��şן�����1� C�U�g�y��������� ӯ���	����
�<� N�`�r���������̿޿� :��)� ;�M�_�qσϕϧϹ� ��������%�7�I� [�m�ߑߣߵ����� �����!�3�E�W�i� {������������ ��/�A�S�e�w��� ������������+��<�Sew� ������^��A�a��B�Bw��Pf�� ����/!/3/E/ W/i/{/�/�/�/�� �/�/??/?A?S?e? w?�?�?�?�?�?�?�? �/�/+O=OOOaOsO�O �O�O�O�O�O�O__�'_9_&O�S���x_�]�rdtS���_�] �_�_�W�����S"oe_8oXoa ��qo goyo�o�o�o�o�ouP��p"|����	`@[oUgy8qK�A\�p���s� A �P�y@h�Q�Q��"����Tk\$���  ��P�PE~�xC�  �I� @oa�<o��p�������@ߏ
f�Q*�����0���PCr� �� 3r �.� @D7�  A�?�G�-��?.I�.@I��A����  ;�	�lY�	 �X  ������� �,� � �����uPK��o�����]K���K]�K	�.��w�r_	�<���@
�)�b�x1�����I�Y�����T;fY��{S���3�����I�>J���;Î?�v�>��=@��'���E��Rѯע�Z���wp��u�� �D!�3��7pg�  �  ��9�͏W���	'� �� u�I� ?�  ��u���:�È��È=���ͱ���@���ǰ�3��\�3��E�&���N�pC�  �'Y�&�Z�i�b�@f�i�n�C����I��C����b���r���`����B �p�Ŕq���}ر�.DzƏ<ߛ�`�K�p�ܖ����������А 4�P����.z��d � �Pؠ?��ff�_��	�� 2p>�P���8.f�t�C>L���U���(.��P��������
ĉ���� x��;e�m���KZ;�=g�;�4�<<�0���%�G��3����p?fff?ذ?y&S���@=0e�?��q�+�rN� Z���I���G���7��� (�����!E0i�T����+��F�p���#��D ��w���� ���//=/(/a/ L/�/p/��/�p�6 �/Z#?�/ ?Y?k?}? ��?�?>?�?�?�?�?�?1O�����KD�y^K�CO�OO�O����ذO�O�O�Oai�b��J��}�DD1����.�D��@�AmQa���9N,ȴA;�^�@��T@|j@$�?�V�>��z�ý���=#�
>\)�?��
=�G��-]�{=����,��C+��B�p���P��6���C98R����?N@��(���5-]G�p��Gsb�F�}��G�>.E�V�D�Kn����I�� F�W��E��'E����D��;n����I��`E��G��cE�vmD���-_�oQ_�o �o�o �o$H3 X~i����� ����D�/�h�S� ��w��������я
� ��.��R�=�v�a�s� ����П����ߟ�� (�N�9�r�]������� ��ޯɯۯ���8�#� \�G���k�������ڿ ſ���"��F�1�C� |�gϠϋ��ϯ����������P(�Q34�] �����Q�	�9�<Oߵ53~�mm�ߎaҀ5Q�߫�aғ�����ߵ1�������1��U�C�y�g��%P�P���! �/��'���
���.������4�;�t�_� �������������� :%��/�/d�������� 7%[Imȏ��027�  cB�S@J@�CH#P	zS@�0@ZO/1/C/ U/g/y/�-�#��/`�/�/�/�/�3?�3V�� @�3��0��0�13��5
 ?f?x?�?�?�? �?�?�?�?OO,O>O�PO�Z@1 ���ۯ��c/�$MR_�CABLE 2�~�� ��TT�����ڰO���O�) �@���C_���_O_ u_7_I__�_�_�_�_ �_o�_�_oKoqo3o Eo{o�o�o�o�o�o�o �o�oGm/�K!�"���O�������$�6���*�Y�** �COM �ȖI�����  �"�4�%% 23456�78901���� ���Ï��� � !�� �!
���M�not sen�t b��W���TESTFEC�SALGR  e�g�*!d[�41�
,k�������$pB����������� 9�UD1:\mai�ntenances.xmlğ����C:�DEFA�ULT�,�BGRP� 2�z�  �� O��%  �%�!1st cle�aning of� cont. v��ilationW 56��ڧ�!0�����+B��*������+��"%��m�ech��cal �check1�  �k�0u�|��ԯ����Ϳ߿�@�~��rollerS�e�w�ū��m�ϑ���ϵ�@�Basi�c quarte�rly�*�<�ƪ,�\�)�;�M�_�q�8��MJ��ߓ "8��� ���ߕ �����+�=��C�g����ʦ�߹���������@�Overh�au�ߔ��?� !x� I�P����}� ��������� $n��� ����)l�ASew ������ � +=O�s�� �����/R� 9/�(/��/�/�/�/ �//�/�/N/#?r/G? Y?k?}?�?�/�??? �?8?OO1OCOUO�? yO�?�?�O�?�O�O�O 	__jO?_�O�Ou_�O �_�_�_�_�_0_oT_ f_;o�__oqo�o�o�o �_�oo,oPo%7 I[m�o��o�o ����!�3��W� �������ÏՏ� 6����l����e�w� ��������џ�2�� V�+�=�O�a�s��� ���ͯ����'� 9���]�������⯷� ɿۿ���N�#�r��� YϨ�}Ϗϡϳ���� ��8�J��n�C�U�g� yߋ��ϯ������4� 	��-�?�Q��u��� ���ߞ��������� f�;���������� �������P���t� I[m����� �:!3EW �{��� �� �//lA/��w/ ��/�/�/�/�/X*�"	 X�/?.?@?�)B a/o?m/o%w?�? �?}?�?�?OO�?�? OOaOsO1OCO�O�O�O �O�O__'_�O�O]_ o_�_?_Q_�_�_�_�_ܫ_�\ Џ!?�w  @�! M? HoZolo�&4o�o�o�o�(*�o** F�@ �Q�V�`o '9�o]o�����/^&�o�� ���/�A�S�e�� �#�����я���� �+�q�����7����� ��k�͟ߟ��I�[� ��K�]�o���C������ɯ��o$�!�$�MR_HIST �2��U#�� 
� \7"$ 23456789013�(;���b2�90/�� ��[���./����ǿ ٿF�X�j�!�3ρϲ� ��{��ϟ�����B� ��f�x�/ߜ�S����� ���߭��,���P���t��=��$�SK�CFMAP  .�U&��b
��� ����ONREL  �$#�������EXCFEN�B�
����&�FN�C-��JOGOVLIM�d#�v���WKEY�y���_PAN������WRUNi�y����SFSPDTYPxM����SIGN�>�T1MOTk�����_CE_GRoP 1��U�� +�0�ow�#d� �����&� 6\�7y�m ���/�4/F/-/ j/!/t/�/�/�/{/�/��/�/?�+��QZ_�EDIT
����T�COM_CFG 1���0�}?�?�?� 
^1SI ЄN����?�?���?$O����?XO78�T_ARC_*��X�T_MN_M�ODE
�U:_�SPL{O;�UAP�_CPL�O<�NO�CHECK ?^�� �� _ #_5_G_Y_k_}_�_�_ �_�_�_�_�_oo���NO_WAIT_�L	S7> NTf1�����%��qa_E�RRH2�����@��?o�o�o�o��O�Gj�@O�cӦm|�"��GAA�Y����[��2#��@"� N_l,��<���?���)��n��bPARAM�b�.���tGO�p8
�.�@� = n� ]�o�w�Q������������Ϗ�)��7��[�m� �����OD�RDSP�C8�O�FFSET_CAqRI0�OǖDISԟ�œS_A�@ARK�
T9OPEN_FILE��1T6�0�OPTION_I�O����K�M_PR�G %��%$*؄���'�WO��Ns�ǥ��G ��u����	 ����Ӧ������RG_DS�BL  �����jN���RIENTkTO���C������A ��U�@IM�_DS���r��V~��LCT �{m P2ڢ�3̹��dҩ���_PEX�@���R[AT�G d8��>̐UP װ�:����S�e�Kωϗ���$�r2G�L��XLȚ�l㰂������� '�9�K�]�o߁ߓߥ� �����������#�5�G���2��v������������ e�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?V?�q1�~?�? �?�?�?�?�?�?O Ox2ODO�yA�a�t@n?~M��~O�O�P�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �O�Oo$o6oHoZolo ~o�o�o�o�o�o�o�o  �_oVhz� ������
���.�@�R�d�QOES�Q�����B�d�ӏ �ʏ��������Y�D�}�0��r����� ����ԟڟ���p���h=�M��q�	`���������c�:�o��¯ԯ����A��  �k�C�C��ڰ"ڰ���~O��  ����-���)�C�  �t�k���g����� Կ��ѿ
�5���_:�����OU���6�_�6�H��n�� � ^��\� @D� M p�?�v�\�?:px�:qC4r�p�(�Ͽ  ;�	l��	� �X � ������ ��, � �������Hʪ�����H����Hw�zH����ϝ�8�B���B�  Xѐ�`�o�*�O�3����t�>u����fC{ߍ��:pB\��
�Ѵ9:q�'�K�t�� ������$���*��� �DP�^��b�g�  �  ��h�����)�	'� �� ��I� ?�  ��'֏=�������t�@����!�b��^;"b�t�U�(�N��r�O  '��E�C����t�C�И��ߗ���jA�@�����%�B�� ��,���H:qDz�k�ߏz����������А #4P���:uz:����	f��?��ff'�&8� ]�m�8:p��C>L�����$�(:p�P��	������:�� x�;e��m"�KZ;�=�g;�4�<<a���E/Tv��b�|��?fff?��?&� )�@=0�%?��%_9�� }!��$�x��/v��/f' ��W,??P?;?t?_? �?�?�?�?�?�?O�? (OOLO�/�/�/EO�O AO�O�O�O�O_�O_ H_3_l_W_�_{_�_�_ 1��_A���eO+o�ORo oOo�o�o�oK/�o�o mo�o*'`+�",�zt���CL�xH��}?������
������u����D1�/n�t��p�q��@I��h~,ȴA;�^�@��T@|j@$�?�V�n��z�ý���=#�
>\)�?��
=�G�����{=���,��C+��B�p����6���C98R����?}p��(���5��G�p��Gsb�F�}��G�>.E�V�D�KL�����I�� F�W��E��'E����D��;L�����I��`E��G��cE�vmD���\�՟��ҟ ���/��S�>�w�b� ������ѯ������ �=�(�:�s�^����� ����߿ʿ�� �9� $�]�Hρ�lϥϐϢ� ��������#��G�2� W�}�hߡߌ��߰��� �����
�C�.�g�R� ��v��������	� ��-��Q�<�u�`�r� �������������'M�(�34�]O!���8h<~�%3~�m�����5Q��������!���  `N�r���	eP@"P��Q �_/V/9/$/]/H)����c/j/�/�/ �/�/�/�/�/!??E? 0?i?T?"&�_�_�?�?�8��?�?O�?O BO0OfOTO�OxO�O�OȾO�O2f?_  cB��pyp$QCHR�	z�p@�N_`_r_ �_�_�_�]c�O�_`�_oo+o?�BcV� @d4��QJc�D
 2o�o�o�o�o�o �o%7I[m���oa ������c/�$PAR�AM_MENU �? ��  DE�FPULSE���	WAITTMO{UT�{RCV�� SHELL�_WRK.$CU�R_STYL�p�"�OPT8Q8�P�TBM�G�C�R_DECSN�p��� �����������-� (�:�L�u�p���������qSSREL_IOD  ��̕�USE_PROG %�z%���͓CCR�pޒ��s1��_HOST !F�z!6�s�+�T�=���V�h���˯*�_TIME�rޖF���pGDEBUG�ܐ�{͓GINP_�FLMSK��#�T�R2�#�PGAP� 2��_b�CH1�"��TYPE�|�P ��������0�Y� T�f�xϡϜϮ����� �����1�,�>�P�y� t߆ߘ��߼�����	� ��(�Q�L�^�p���%�WORD ?	��{
 	PR<�p#MAI��q"gSUd���TE���p#��	1���CO�Ln%��!���L�� U!��F�d��TRACECTL� 1� �q� �{ |#�����_�DT �Q� ��z�D� � � K`��c`��_`���� ������1CU gy������ �	-?Qcu �������/p/)/;/M/ � b �@P"M`P" k`P"��h/z/�/�/�/ �/�/�/�/
??.?@? R?T/~?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_�_�_�_��Z5o o*o<oNo`oro�o�o �o�o�o�o�o& 8J\n���� �����"�4�F� X�j�|�������ď֏ �����0�B�T�f� x���������ҟ��� ��,�>�P�b�t��� ������ί���� (�:�L�^�p������� ��ʿܿ� ��$�.� oP�b�tφϘϪϼ� ��������(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
 .@Rdv��� ����*< N`r����� ��//&/8/J/\/ n/Dϒ/�/�/�/�/�/ �/?"?4?F?X?j?|? �?�?�?�?�?�?�?O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZl ~������� � �2�D�V�h�z�����������$PGT�RACELEN � ��  ������Ά_�UP ���e��������΁_CFG ۦ��烸�
����*�:�D�O���O��  �O��DEFSPD ��������΀H_�CONFIG ����� ��j��dĔ�݂ ���ǑP^�a�㑹���΀IN�TRL ���=�8^���P�E��೗����*�ÑO�΀LID����	T�LLB� 1ⳙ 5��BӐB4��O� 䘼����Q� << ��?�������M� 3�U���i���������@ӿ��	�7�T�Ϣ k�b�tϡ�诚���������S�GRP 1�爬���@A!����4I���A� �Cu�C�OCjVF�/��Ȕa�zي�ÑÐ�t��ޯs���#´�ӿߨ�B�����������A�S�?&�B34�_�������j����� �����	�B�-���Q����M�������  Dz����.�����& L7p[��� ����6!Z�h)w
V7.10beta1*��Ɛ@�*�@��) @�+A� Ē?��
?fff>�����B33A�Q�0��B(��A���AK��h�����//'/9/P�p*�W�ӑ�n/�/�%����R�fh����*���P2� LR��/�/�/�/�/H?$�Ĕ�I�u�&: ���?��x?�?A���lP!\3 Bu�B��?��5BH�3[4���o��4��[45��/B\3x3Dx�?YO�?aOkO}O�<<�R@� �O�C�O�O�O�O�DA��X�KNOW_M � Z�%�X�SV 賚ڒ�� �_�_�_?�_�_�_o�����W�M+�鳛� ��	@�3#����_�o�\A���
]bV4�@ u��u��e�o�l,�X�+MR+��JmT3?���W�1C{�OADB�ANFWDL_V�S�T+�1 1����P4C���[�� i/�����?�1� C���g�y�������� ӏ�*�	��`�?�Q��c��w2�|Va�up�#<ʟ���p3��Ɵ؟Ꟃw4��+�=���w5Z�l�~����w6 ����ѯ㯂w7 ��$�6��w8S�e�w���V�wMAmp�������OVLD  ⩻yo߄rPAR?NUM  �{+ø��?υqSCH�� �
��X���{s��UPDX�)ź��Ϧ�_CMP_@`���p�|P'yu�ER_wCHK���yq0bb3��.�RSppN?Q_MOm��_}�~��_RES_G�p쩻
�e�����0� #�T�G�x�k�}��� �����������׳���������:�Y�^� ��Y�y������Ӭ��� ������������ R�6UZ�ӥ�u�<���V 1�Fvp�Va@k�p��T?HR_INRp���(byudMASS6 Z)MNG�MON_QUEUE �uyvup\!U��N�UZ�NW��END��߶�EXE����BE����OPTIO���ۚPROGR�AM %z%��~ϘTASK�_I��.OCFG� �z+�n/� D�ATACc�+�@ �KP@2 �??/?A?S?]51 s?�?�?�? �?�6p1�?�?�?O"O�,F�!INFOCc��-��bdlO~O�O�O �O�O�O�O�O_ _2_ D_V_h_z_�_�_�_�_��_�/A@FD��, �	��!��K_�!�8�)fN!fENB��0m���Pf2YokhG�!2��0k X,	�	d�=��·o�	��e�a$�pd��i�i��g_EDIT ���/%7�����*SYSTEM*�upV9.4010�7 cr7/23/�2021 A���Pw��PRG�ADJ_p  h� $X[�p W$Y�xZ�xW�x�қtZқtSPEE�D_�p�p$NE�XT_CYCLEΝp���q�FGތp ��pAL�GO_V �pNYQ_FREQ�WIN_TYP�q])�SIZ1�O��LAP�r!�[��M�+����qCREATsED�r�IFY�rn@!NAM�p%h��_GJ�STATU|��J�DEBUG�r�MAILTI��ΰ�EVEU��LA�ST�����tELE�M� � $�ENAB�rN�EA�SI򁼁AXIS�p$P߄����~�qROT_RA" ��rMAX ��qEZ��LC�AB
����C D_LVՁ`�B�AS��`�1�{���_�� ��$x���R�M� RB�;�DIS<����X_SPo�΁������t�P� |� 	� 2 m\�AN�� ��;�����Ӓ�� ��0�PAYLOx��3�V�_DOU�q�S���p�tPREF�� ( $GWRID�E
���iR���Y� �p�OTOƀ�q  �p��!�p��k��OXY� � w$L��_POp|�נVa�SRV���)���DIREC�T_1� �2(�3�(�4(�5(�6(�7�(�8� ��F��A��� $VAL|u�GROUP��ݑ��F�� E!��@!�������RAN泲����R��/���TOTA���F��PW�I|=!%�REGEN#� 8�������/���ڶ�nTzЉ���#�_S����8�(�V[�'���4���GRE��w����H��D�����V_H���DAY3�V��S�_Y�Œ;�SUM�MAR��2 �$CONFIG_�SEȃ���ʅ_R�UN�m�C�С�$C�MPR��P�DE�V���_�I�Z�P�*Ӥ���ENHAWNCE�	�
�q��1���INT�B�qM)b�q�2K��n��OVRo�PGu��IX��;���OVC�T�����v�
 4 �����a˟��PS�LG"�� \ ��;��?�1���S8Ɓϕc�U�����Ò�4�U�q]�Tp>� (`�-���rJ<�O� CK�I'L_MJ���VN�+�&�TQn{�N5���MC�ULȀD�V(��C6�P_�຀@�M�W�V1V�V1d�2�s�2d�3s�3d�4s�4d��'�	��������p	�IN	VI#B1qp1� 2!pqT/,3 3,4 4,�p?��;��A����N�������PL��TORr3�	���[�SAV���d�MC_FO�LD 	$S�L�����M,�I��L� �pL�b���KEEP_HNADD	!Ke�UoCCOMc�k0��
�lOP����pl��lREM�k��΢���uU��ekHPW� ;KSBM��Š?COLLAB|�Ӱhn��n�+�IT��O��$NOL�F�CALX� �DON��r���� ,恠FL���$SSYNy,M�C=�����UP_DLYz�qs"DELA� �����Y(�AD���$TABTP_R��# �QSKIP�j% ����OR0� �6�� P_���  �)���p7��%9�� %9A�$:N�$:[�$:h��$:u�$:��$:9�q�{RA�� X������MB�NFL#IC]��0"�U!�o���NO_H� �\��< _SWITCH�k�RA_PARA{MG� ��p��U��WJ��:CӾ��NGRLT� O�O�U�����X�<A��Tc_Ja1F�rAPS��WEIGH]�J43CH�aDOR��aD���OO��)�2�_FJװ���sA�AV��C�H�OB.�.�`�J2��0�q$�EX��T$�'QIT��'Q�pG0'Q-�GADC�m" � ��<��
�R]��
H���RG�EA��4��U�FLaG`g��H��ER�	�SPC6R�rUM�_'P��2TH2N�o��@Q 1 ����0����  D �وIi�W2_P�25cS��|��+�L10_CI�q�pe� �p k����UՖD��zaxT�p�Q(�;a� �c��޲+�i�_h���` P`DESsIGRb$�VL1:i�1Gf�c�g10�_�DS��D�ׁw�POwS11�q l�p`r��x1C/#AT��B��U
WusIND��}�mqCp�mq`B�	�HOME�r 	aBq2GrM_q���� ?t3Gr��� ��$���?t4GrG�Y�k��}�����!�?t5Gr�ď֏������w6GrA�S�e�w������!@s7Gr��П�P����*�8Gr;�@M�_�q�����*�S >�q    �@s�M��P<s�K@��!� T`M��M�IO���m�I��2�OK _�OPy��� »Q*�P�OWE" �7�x EQ 8� � �#s%Ȳ$DSB�o�GNA�b� Cx�P2�BS232S�'$ �iP��xc�gICE<@%�PE`�2� @IT��P�OPyB7 1�FLOWУTRa@2��U$�CqUN��`�AUXT��|2Ѷ�ERFAC3�ڰUU�QRS;CH��% t<�_9�EЎA$FR?EEFROMЦ��A�PX q�UPD�"YbA�PT.�pEE�X0����!�FA8%bҬ��RV�aG� &  C�E�" 1�AL�  ��+�jc'��D�  ?2& �S\PcP?(
  �$7P�%��R�2� ��T�`A9XU���DSP���@@�W���:`$��RNPн%�@����K��_McIR�����MT��AP���P"�qD��QSYz������QP=G7�BRKH����� AXI�   ^��i���1 ����OBSOC���N��DUMMY16�1o$SV�DE���I�FSPD_OV%R79� D���ӓOR��֠N"`��F�_����@OV��SFN�RUN��"F0�̊���UF"@G�TO�d�LCH�"�%REGCOV��9@�@W�`@&�ӂH��:`_0��  @�RTINsVE��8AOFS��9CK�KbFWD���`���1B��TR�a�B �FD� ��14= B1pBL� �6� A1L�V��Kb�����#��@+<�AM�:��0��j��_M`@ ~�@h���T$X`�x ��T$HBK ���F��A�����PPA�
��	�������DVC_DB�3@pA�A"D��X1`�X3`@��S�@�`�0��U���h�CABPP
R�S  #��c�B�@���G�UBCPU�"��S �P�`R��11)A�RŲ�!$HW_�CGpl�11� F&A1�Ԡ@8p�$UNI�Tr�l e ATT�RIr@y"��CYC�5B�CA��FLTR_2_FI�������2bP��CH�K_��SCT��F�_e'F_o,�"�*FqS�Jj"CHA�Q��'91Is�82RSD�����1���_T`g�`� i�EM��NPMf�T&2 8px&2- �6DIAGpE?RAILACNTB�Mw�LO@�Q��7&��PS��� � ���PRBSZ`�`�BC4&�	��FUuN5s��RIN�P`Zaߠ�07Dh�RAH@���`� `C�@�`C��Q�CBLCUR�uH�DA�K�!�H�HD�Ap�aA�H�C�ELD@������C��jA�1��CTIBUu�8p$CE_RIA�QVJ�AF P��>S,�`DUT2�0C��}�;OI0DF_aLC�H���k�LML}F�aHRDYO���RG�@HZ0��ߠ|�@�UMULSE�Pt�'3iB$J���J����FAN_�ALM�dbWRNeHARD��ƽ�	P��k@2aN�r�J�Y_}�AUJ R+4~�TO_SBR���~b�Іje 6?A�cM/PINF��{!�d��A�cREG�NV���ɣZ�D��NF9LW%6r$M�@� ���f� �0 h'uC�M4NF�!�ON 	 e!e#�(b*r3F�3G �	 ���q)5�;$�$Y�r���u�_��p*$ �/�EG@����F�qAR��i���2�3��u�@<�AXE��R�OB��RED��W�R��c�_���SY�`��q� ?�SI�WR1I���vE STհ��(� d���Eg!���t8��^a��B���񐆹9�3� OTO�a����ARY��ǂ�1������FIE����$LINK�QGT5H��T_�������30���XY�Z���!*�OFF������ˀB��,Bl���e���m�FI� ��C@Iû�,B��_J$�F������S`����3-!$ 1�w0���R��C��,�DU���3�P�3TUR`XS.�Ձ�b1XX�� ݗFL�d�`��pL�0���34��^�� 1)�K��	M�5�5%B'��ORQ�6��fC����0B�O;�D�,��p����a�OVE��rM�����s2��s2� �r1���0���0�g /�AN=!�2�DQ�q� ��q�}R�*��6���0�s��V���ER��jA�	�2E��.�C��A���0��XE�2Ӈ�A��AAX��F��A� N!�SŴ1_��Q_Ɇ� ^ʬ�^ʴ�^��0^ʙ�^ʷ�^�1&�^ƒP[� �PkɒP{ɒP�ɒP�� �P�ɒP�ɒP�ɒP������ɪ �R>�DEBU=#$8ADc�2����
�AB�7����9V� <" 
��i �q��-!��%��׆��� ���״����1�י������JT��DR�m�LA�B��ݥ9 FGR�O� ݒ=l� B_ �1�u���}��`����pޥ��qa��AND������qa�  �Eq��1��A@�� ��NT$`��c�VEL �1��m��1u���QP��Fm�NA[w�(�CN1�� ��3줙� ��SERVEc�p+� $@@d@��!���PO
�� _�0T� !��򗱬p�,  $T�RQ�b
(� -�DR2,+"P�0_ . l"@!�&'ERR��"I� q𜍴~TOQ����L��p]�e���0G��%����RE�@ �/ ,��/I -���RA� 2.3 d�& �" 7 0�p$&��2dtPM� �pOC�A�8 1  pC�OUNT���FZ�N_CFG2 4B �f�"T�:#��Ӝ� 
`�s/3 ���M:0�R��qC@��/�:0�FA1P��?V�X������r���� �P�:b
HELpe�4 5��B_wBAS�cRSR�f� @�S�!QY 1T�Y 2|*3|*4|*U5|*6|*7|*8��L!RO�����NL�q �AB���0Z �ACK��INT�_uUS`�Pta9_cPU�>b%ROU��PH@�h9#�u`w�9��TPFWD_KA1R��ar RE���PqP��A]@QUE�i@&��	�f�>`QaI`���9#�j3r��f�SCEME��6��PA�7STY4SO�0�DI'1�`���18�rQ�_TM�cMANR�QXF�END��$KEYSWIT�CHj31:A�4HE�	�BEATM�3PE�pLE��1��H�U~3F�42S?DD_O_HOMBPO:a60EF��PRr��(*�v�uC�@O�Qo ��OV_Mϒ��E�q�OCM���7��� 7&HK�q5 �D��g�Uj�2M��p�4R��FORC.�cWAR����:#�OM�p 6 @��Ԣ�v`U|�P�p1(�V'p�T3�V4�� ���S#O�0L�R7<��hUNLOE0h-dEDVa ���@�d8 <pAQ9�>l1MSUPG�Ua�CALC_PLA5Ncc1��AYS1�1�:b�9 � X`��P �q;a�� ��w��2��j�M$P��`���fyt$��rSC�M�pm�q ���aq���0�tYzZzEU�Q�b�� T!�Hr�p�Pv	NPX_AS�f: 0g ADD|��$SIZ%a�$VA��MU/LTIP�"ns�P�A�Q; � A$T9op�B���rS���j!C~ �vFRIF��2S�0�YT�pN=F[DODBUX�B�0�u&�!���CMtA�������������|Z ��< � �pƛTEg�����$SKGL��T��X�&{𷃥㰀��STMT<e�ЃPSEG�2���BW���SHOW�؅�1BAN�`TP�O���gᣥ�������
V�_G�= ��$PC���O�kFB�QP\�SP�01A&0^�.VDG���>� �cA00�����P���P��P�P���P��5��6��U7��8��9��A�� b`���P��w᧖��!F����h���1��v�Th�י1�1�1��U1�1�1%�12�U1?�1L�1Y�1f�U2��2��2��2ʙU2י2�2�2��U2�2�2%�22�U2?�2L�2Y�2f�U3��3��3��3ʙ3י3�3���Ȫ�3�3%�32�3�߹3L�3Y�3f�4���4��4��4ʙ4�י4�4�4��4��4�4%�42�4�߹4L�4Y�4f�5���5��5��5ʙ5�י5�5�5��5��5�5%�52�5�߹5L�5Y�5f�6���6��6��6ʙ6�י6��6�6��6��6(�6%�62�6�߹6L�6Y�6f�7���7��7��7ʙ7�י7��7�7��7��7(�7%�72�7*߹7L�7Y�7f�OR�V�`_UPD��?s �c 
A�����@ x $gTOR�1T�  �caOP �, ZQ_7�RE^��� J��S�sC�A��_Ux�p�7bYSLOA"A � �u$�v���w�@���@��bVALUv10�6�=F�ID_L[C:�HI5I�R$FI�LE_X3eu4$��C��SAV��B� hM �E_BL�CK�3�ȁ�D_CPU��p��p5�hzmpY��R3R �C � PW���� 	�!LAށ�SR�#.!'$RUN�`G@%$D!'$�@ G%e!$e!'%HR03$�� '$���T2�Pa_LI�RD � � G_O�2>�0P_EDI�Rlp�T2SPD�#E��"i0ȁ�p	���DCS9@G)F� � 
$JPC�71q�� S:C;C�9$MDL7�$5P>9TC�`@7U�F�@?8S� ?8CO�Bu �@��"|�L�G��P;;� 9�:;`�TABU�I_�!L�HGb�% �FB3G$��3A�sR�LLB_AVAI�B�Q�3�!I $� SEL� NẼ�@RG_�D N��Ta?��3SC��PJ �1/AB2�PT�R<D_M]`L��K \M f/QL_���FMj��PGi�Ut9R�6��PS_��P\� �p�EE7B��TBC2�eL ����``�`b$�!F�T�P'T�`TDCg�� BPLp�sNU;WTH��qhTgtW�R�2$�pERV�E.S�T;S�Tw�R_�ACkP MX -$�Q�`.S�T;S��PU@�`IC�`LOMW�GF1�QR2g��`��p�S�ERTIA�d^0iP�PEk�DEUe�LACEMMzCC#c�V�B�rpTf�edg�aTCV8�l�adgTRQ�l�e��j|�Scu��edcu�J7_ 4J!��Se)@qde�Q2�0����1�PRcuPJKlvV�K<�~qcQ~qw�spJ�0��q�sJJ�sJJ�sAAL�s�p�s�pȲv���r5sS�`N1@�l�p�k�`5dXA_́�QCF�BN =`M GROU ���bh�NPC0sD�R�EQUIR�R� E�BU�C�Q�6g0 �2Mz��Pd�QS�GUO�@�)AP�PR0C7@� 
$:� N��CLO� ǉ�S^U܉Se
Q�@A.�"P �$PM]P�`8�`sR�_MGa!��C���+��0�@,�B{RK*�NOLD*�SHORTMO�!Hm�Z��JWA�SP�t p`�sp`�sp`�sp`�s(p`�A��7��8sQ|�RTQ� m���R.Q�cQ�PATH�*� �*��X&����P�NT|@A��"p��� �IN�RU�C4`a��C�`UM��Y
`�)p��>��Q��cP���p��PA�YLOAh�J2LN& R_Am@�L ������+�R_F�2LSHR�T/�L�O���0���>���ACRL0z�p�y�ޤsR9H5b$H+���oFLEX��XPJVR P��_._��_�_����US :�_�Vd`0�G��_`tQd`�_�_lF1G� �ũ�o0oBoTofoxo��E�o�o�o�o�o�o �o ����wz3lt�����3EWF�^zT!��X�'qju�� uu~�W؁���p�u��u�u�u���� 9	��(�T �P5�0G�Y�' AT��l��pEL0�_B��s�J��Sz�JEW�CT�R7B`NA��d�H�AND_VB��(��TUO@`+�`TSW8F�A�V� $$M� �e G�AV�Qs�De�oAA��@�	�$�A5�G�AU�A�d�� 6��G�DU�D�d�PD�G/ -ST�I�5V�5Ng�DY F ��+�x����P&� G�&�A��lw�o�Q�k�P������ʕӕܕ���QJUW 7 �� ��3%遞?!ASYMT���m�T�V�o�A�t�_SH�~������$ ����Ưد�J񬢐��#39"���_VI���`8�q0V_UCNIrS�4��.�Jmu �2��2A��4X��4�6 a�pt�������&E_��������E��CH~( X ̱l���TOc�PPСVsSvD�US�RU�P������z@�D�A}@_�5�U��P�EyAa��RP�ROG_NA��}$�$LAST����CANs�ISz@XYZ_SPu�DW]R@Ͱ,VSV@�E1QsENc��DCUR�H�����HR_T��YtQ9S�d���O�T�&uP?�Z) ��I�!A�D�� �Q���#�S����3��vP [ � ME�O��R#B�!T�PPT0F@1�a��̰� h1a�%iT0� $�DUMMY1��o$PS_��RF���% $lfװFL�A*�YP�bc?$GLB_TI �Up�e`ձ��LIF(!�\����g`OW��P��eVOL#qLb �a_2��[d2[`����b�P�cZ`T�C��$BAUD,v��cST��B�2g`�ARITY0sD_[WAItAIyCJ�2�OU6�ZqyyT�LANS�`�{S�SyZc��BUF_�r��fиx�PyyCHK]_�@CES��� +JO`E�aA�x�bUBYT���� �r�.�.� ��aA���M�������Q] �Xʰ����ST����SBR@M21�_@��T$SV_cER�b����CL�`ʐ�A1�O�BpPGL�h0EW(!^ 4 �$a$Uq$�q$W�9�A��@R��)�ӃUم_� "��D$GI���}$ف �^
Ӄ�(!` L��.��"}$F�"E�6�NEAR��B�$F}��TQL�����J�@R� �a7�$JOI�NTa�)�ԂMS�ET(!b  +�Ec�2�^�ST�Ĕ^�(!_c�  ��U��?���LOCK_�FO@� �PBGLmV��GL'�TE�@sXM���EMP���:�K��b�$U�؂a�2_���q��`<� �q�^��C�E/�?��� $KA�Rb�M�STPDRqA܀����VECX������IUq�av�H=E�TOOL����V��REǠIS3d��6��ACH̐�m b^QONe[d3����IdB�`@$R�AIL_BOXE:a���ROB�@D��?���HOWWA�R0Aa�i`-�ROLMtb��$�*���T��`ܱ���O_FU�!>��HTML58QS��� e�MBՀ�(!d ����@�(!e��������Ĕ}p(!'f t��m�^a��Xt��B�PO��A	IPE�N���O�����q��AORDEaD�m �z�XT`���A)�bPMO�P �g D �`OB�����ǯ�Uc�`���� ��SYS��A�DR��pP`U@^  �h ,"��f$�A��E��E�QP�VWVA�Qi Ǥ �@ق�UPR|�B�$EDI�A�d�VSHWRU��z���IS�Uq�pN�D�P7���G�HEA�D�! @���!i�K�EUqO`CP)P��J�MP��L�U' RA[CE�Tj����IL�S��C��NEx���TICK�!MKQC_��H=Nr�k @���HWC��PHVF��`S�TYeB+�LO�aPg���[�C�l3�
�@��F%$A��D=��S�!$�1�p a�e��q�ePv HVSQU̩�#LO�b_1TE�RC`! S?�m 5���R�m@3����ܡ�O`	c IZ�d�A�eha�qtb�}�hA}pP~r��_D)O�B�X�pSSQ�S'AXI�q��v�bS��U�@TL���RE3Q_ܠ��ET���`��CY%��FY'��A,f\!\d9x�P� E�SR$$nl-�w �����c
�uV
Qh(�AA���dC`�A�@�	�Y��D���p�E"�	CC�C���/�/�/	4NASS}C�` o h��cDSm��Q[`SP�@&�AT� 
R��L��XbADDR�s�$Hp� IF�Ch�_'2CH���pO����- �TUk�Ir p�CUCp#�V��I�Rq�4��T�c��
K�
��V*����Pr \z�D�� ��|,K� P�"CN���*CƮ��!�TX_SCREE��s�Pp@�INA˃<�4��D�a����`t Tᫀ�b����O Y6`���º�U4h�RR��������R1�TC�UE���u �j �qz`S�́��RSML��U`����V�1tPS_���6\��1�9G\���C8��2@4 2��0�Ov�R��&F�AM_TN_FL*�`Q�W� ��PBBL_r/�WB`�Pw ���j�BO ��BLE"�Cg�R"�DRIGH�tRD��!CKG�RB`�ET���G�AWIDTHs���RB�h�a�r<@I��EYհRx d�ʰ����z�`y�BACK��h��>U���PFO��nQWLAB�?(�PyI��$URm��~P��P�PHy1 �y 8 $�PT!_��,"�R�PRUp��s5���TO%!t�z�V�ȇ�pU�@�SR ���LUM�S�� GERVJ�� PP���T{ � " G�E�Rh� �¯�LP$AeE��)^g��lh�lh�ki5ik6ik7ikpP`�Z�x�����$u1��p�Q wzQUSRلO| <z��PU2��a#2�FOO 2�PR�I*m9�[�@pTR�IPK�m�UN[DO��})���0Yp��y����h�����p ~�Rp�qG ��T���-!�rOS2��vR��2�s�CA�����r`�$��h�UIaCA���p�3Ib_�sOFFA�*D@���Ob�r�a��L�t��GU���Ps������+QS�UB`� ��E_�EXE��VeуsW]O� �#��wF��WAl�p΁fP=
 V_DB��$Z!pT�pO�V░̷��3OR/�5�RA�U@6�TK���_<_���� |j ��OWNj�34$S#RC�0`���DA���_MPFI����ESP��T�$0��c���g� n�z�E!�# `%�ۂ34J���7COP��$`��p�_���/�+�6���C�T�Cہ�ہ�� ��DCS��P�4�COMp�@�;��O`�=��b�K�^�/�VT�qU'���Y٤Z���2���@p�w#SB�����2�\0˰_��M8��%!]�DIC#��sAY�3G�PEE�@T�QS�VR1���eQL�� a��P�D  ��f�z��f�> ����6���A�t�b# �~L2SHADOW���#ʱ_UNSCA�d�׳OWD�˰DG�DE#LEGAC�)�q'
�VC\ C>��� v����だm�RF07���7�d`C2`7�DRIVo���ϠC�A]�(��` ���MY_UBY�d?Ĳ��s��1�� $0�����_ఆ����L��BM�A$n�DEY	�EXp@,C�/�MU��X��,���0US����;p_R@"1�0p#�2�G�PACIN*���RG��c�y�:�y��sy�C/�RE�R"!�qq�y�D@� L 
!�G�P�"��0�	R�pD@�&P�Px1Q���	.���RE��SMWq�_Ar�u@+�{�Oq�AA/�3�h�EZ�U���� �y@�HK���P�J��_/�Q0{�EA�N��ۀ2�2�C�MwRCVCA� �:`GORG��Q�dR	��8L�����REFoG�� ���!�+`	�p��������<���q�_ ����r�����`C���p��Q�@D� ��0��!��#q�š�OUx����?� ����2�J@0� 1�*p�������0 UmL�@��CO�0f)��� NT� [��Z�Qf�af% L飏��Q��a��VIAچ� ̈́ÀHD7 6P$�JO�`oB�$�Z_UPo��2Z_LOW��$�QiB<n��1$EP�s��y�� 1!f m�� 1¦4� 5��PA�A �C7ACH&�LO�w@�ВQB���Cn�%I#F^��Tm��N��$HO2�32{��Uÿ2O�@���R`o��=a��ƐVP��<X@A"_SIZ&�K$�Z$�F(�G'���CM]Pk*FAIo�G���AD�)/�MR1E���"P'GP�0����9�ASYNBUFǧRTD�%�$P!��COLE_2D_D4�5W�sw�~�U��QO��%ECCU��VEM��v]2�VIRC�!5�#�2��!_>�*&�pWp��AuG	9R�XYZ@�3�W���8��4+Q2z0T"��IM�16��2P�GRABB��q��;�LERD�C ;�F_D��F�fC50MH�PE�R[����l�JRLAS��@��[_GEb�� �H൑~23�ET@����"���b��I�D��ҙ6m�BG_LEVnQ{�PK|Л6\q���GI�@N\P4� ��P��!g�dr�IS� �NRT��Lʁc�Ų��#a��c"!D�qDE����Xа(�X�� ��2��
d��pzZ���d�c*���D4q���2puT��U&�� $�ITPr9p[Q��Փ�V�VSF$�d� a fp/�f�UR&�kR`MZu�dr���ADJ`C�� Z�DVf� D�XA�L� � 4 PER�IKB$MSG_Q3$Q!o%�p��p'��dr:g�qQ�.��XVR\t��B�p�T_\��R�ZABC"����Sr����
sA�aACTVS�' � � �$|u�0�cCTIV�Q!IOu¥s&D��IT�x�DVϐ�
x�P���!��&�pPS���� �#��p!���q!LSTD��!�  �_ST����wrq�CHx�� L-�@��u��Ɛ*���P GNA�#�C�!q�_FUqN�� �ZIPu�3�HR�$L���}�AZMPCF"���`bƀ�rX�ف��LNK��

Ł�0#�?� $ !��^ބCMCMk�C8��C"����P{q O$J8�2�D6! >�O�H���T���2������M���UX�1݅UXE1Ѡ��1C���Y����������˗7�FT�FG>������Z���� �k�� W�YD'@_ � 8n�R� �Uӱ$HEIGHd�:h?(! 'v���P���� � 1Gd��qp$B% � <E��SHIF��hRVn�F�`�HpC� 3�(�8H`O�ѡ��C��+%D	�"�C�E�pV�1Qp��PH�ERs� � ,�! M�c�u��$P�OWERFL  )�p|����|�p��RG�`  7������AЋ  ��?�p���pdv��NSb ����?� � Bz|� l�  �<@�|�Z�|�%� ��˃����ŵ��� 2ӷ�� 	UH��l&��౿>���A |�ɻt$��*��/�� **:���p��ȥ��͘���������ɘ��|����� 5�������%ߟ�I� [߉�ߑ������� ����w�!�3�a�W�i� ����������O��� �9�/�A���e�w��� ����'���� �=O}s��� ����k'U K]������ C/��-/#/5/�/Y/ k/�/�/�/?�/�/? �/?�?1?C?q?g?y? �?�?�?�?�?�?_O	O�OIO?OQO�� 	 �O�O�O_�E��3_����O`_�O�_�_÷P?REF Ӻ�p��p
��IORI�TY ?p|����p����pSPL`z����W�UT�VqÈ�ODU,~�����_?�OG��Gx��R��,f�HIBqOy�|kTOENT 1��~yP(!AF_t��`�o�g!tc�p�o}!ud��o)~!icmX�0bXY̳�kw �|�)� �����p����u ������N�5� r�Y�������̏�����*/c̳ӹ���xE�W�|�>���F���/��4���|���,�7�A��,  ��P����%�|�'���Z��h�z�茯��|��ENHANCE 	#��7�A9�d����� ' �,f�T
�_�Sz����PORTe��rb�@�U��_CARTREP�P|r|brSKSTAgޛkSLGS�`�k����@Un?othing�� ����Ϳ>�P�b�To���TEMP �?isϨE/�_a_?seibanm_�� i_�����0��T�?� x�cߜ߇ߙ��߽��� ����>�)�N�t�_� ������������ �:�%�^�I���m��� �������� ��$ H3lWi��� ����D/ hS�w���u�>��VERSI�P=g�  dis�able��SA�VE ?j	�2670H705��k/!�m//*�/ 	�(%b�O�+	�/�Se?6?H?Z?l?z:%<�/�?4�*']_j` 1�kX �0ubuE�?OqG�P/URGE��Bp`�ncqWF<@�a�TӒ*f�W�`]Daa�WRU�P_DELAY �z�f�B_HOT %?e'b��O�nER_NORMA�L�HGb�O%_�GSE�MI_*_i_�QQS�KIP�3.��3x ��_��_�_�_�]?e o+goKo]ooo5o�o �o�o�o�o�o�o�o 5GYi�}� ������1�C� U��y�g����������я����-�?�7%��$RACFG ��[ќ�3�]�__PARAM�Q3y��S @И@`\�G�42C۠��2M��CbFB�B]��BTIF���J]�C_VTMOU������]�DCR�3��Y ��UB�h�B�@���4>V�h9w�X;�]�>�>��v��_����;e��m���KZ;�=�g;�4�<<����f@����� �5�G�Y�k�}��������ſ׿���xUR�DIO_TYPE�  �V�5��ED_PROT_a�&g>��4BHbC�EސSǆQ2c� ��B�ꐪϸ� ��ϐ����&�ݹ� W�V_~�o����߱� ��������A�O�m� r���9������� �������=�_�d��� ������������� ��'I�Nm�� �������# EJi+k�� ����//4/F/ /g//�/y/�/�/�/ �/�/	?+/0?O/?c? Q?�?u?�?�?�?�?�?�?;?,O��S�INT� 2�I���l�G;� jO|K��鯤O�f�0 �O�K�? �O�?___N_<_r_ X_�_�_�_�_�_�_�_ �_&ooJo8ono�ofo �o�o�o�o�o�o�o" F4j|b�� �������B��O�EFPOS1 �1"�  xO��o×O����ݏ 鈃���Ϗ0��T�� x����7���ҟm��� �����>�P����7� ������W��{���� �:�կ^�������� ��S�e��� ��$Ͽ� H��l��iϢ�=��� a��υ�� ߻���� h�Sߌ�'߰�K���o� ��
��.���R���v� ��#�5�o������� ���<���9�r���� 1���U����������� 8#\����? ��u��"�F X�?���_ ��/�	/B/�f/ /�/%/�/�/[/m/�/ ?�/,?�/P?�/t?? q?�?E?�?i?�?�?O (O�?�?OpO[O�O/O �OSO�OwO�O_�O6_ �OZ_�O~_�_+_=_w_ �_�_�_�_ o�_Do�_�Aozocf�2 1 r�o.oho�o�o
o .�oR�oO�#� G�k����� N�9�r����1���U� ���������8�ӏ\� ��	��U�����ڟu� ����"����X��|� ���;�į_�q����� �	�B�ݯf����%� ����[���ϣ�,� ǿٿ�%φ�qϪ�E� ��i��ύ���(���L� ��p�ߔ�/�A�Sߍ� ������6���Z��� W��+��O���s��� ������V�A�z�� ��9���]������� ��@��d��#] ���}�*� '`���C� gy��&//J/� n/	/�/-/�/�/c/�/ �/?�/4?�/�/�/-? �?y?�?M?�?q?�?�? �?0O�?TO�?xOO�O<�o�d3 1�oIO [O�O_�O7_=O[_�O __|_�_P_�_t_�_ �_!o�_�_�_o{ofo �o:o�o^o�o�o�o �oA�oe �$6 H�����+�� O��L��� ���D�͏ h�񏌏�����K�6� o�
���.���R���� �����5�ПY���� �R�����ׯr����� ����U��y���� 8���\�n������� ?�ڿc�����"τϽ� X���|�ߠ�)����� ��"߃�nߧ�B���f� �ߊ���%���I���m� ��,�>�P������ ���3���W���T��� (���L���p������� ����S>w�6 �Z����= �a� Z�� �z/�'/�$/]/ ��//�/@/�/�O�D4 1�Ov/�/�/ @?+?d?j/�?#?�?G? �?�?}?O�?*O�?NO �?�?OGO�O�O�OgO �O�O_�O_J_�On_ 	_�_-_�_Q_c_u_�_ o�_4o�_Xo�_|oo yo�oMo�oqo�o�o �o�o�oxc�7 �[����>� �b����!�3�E�� ��ˏ���(�ÏL�� I������A�ʟe�� �������H�3�l�� ��+���O���ꯅ�� ��2�ͯV����O� ����Կo�����Ϸ� �R��v�Ϛ�5Ͼ� Y�k�}Ϸ���<��� `��τ�߁ߺ�U��� y���&�������� ��k��?���c���� ��"���F���j���� )�;�M��������� 0��T��Q�%��I�m��/�$5 1�/���mX ���P�t�/ �3/�W/�{//(/ :/t/�/�/�/�/?�/ A?�/>?w??�?6?�? Z?�?~?�?�?�?=O(O aO�?�O O�ODO�O�O zO_�O'_�OK_�O�O 
_D_�_�_�_d_�_�_ o�_oGo�_koo�o *o�oNo`oro�o�o 1�oU�oyv� J�n����� ��u�`���4���X� �|�ޏ���;�֏_� �����0�B�|�ݟȟ ���%���I��F�� ���>�ǯb�믆��� ���E�0�i����(� ��L���翂�Ϧ�/� ʿS�� ��LϭϘ� ��l��ϐ�ߴ��O� ��s�ߗ�2߻�V�h� zߴ�� �9���]��� ���~��R���v�����#�	6 1 &������������� ��}���<��` ����CUg� �&�J�n	 k�?�c��/ ���	/j/U/�/)/ �/M/�/q/�/?�/0? �/T?�/x??%?7?q? �?�?�?�?O�?>O�? ;OtOO�O3O�OWO�O {O�O�O�O:_%_^_�O �__�_A_�_�_w_ o �_$o�_Ho�_�_oAo �o�o�oao�o�o�o D�oh�'� K]o�
��.�� R��v��s���G�Џ k�􏏏���ŏ׏� r�]���1���U�ޟy� ۟���8�ӟ\����� �-�?�y�گů���� "���F��C�|���� ;�Ŀ_�迃������ B�-�f�ϊ�%Ϯ�I� �����ߣ�,���P�<6�H�7 1S��� �I��߲������� 3���0�i���(�� L���p�����/�� S���w����6����� l�������=���� ��6���V�z � 9�]�� �@Rd��� #/�G/�k//h/�/ </�/`/�/�/?�/�/ �/?g?R?�?&?�?J? �?n?�?	O�?-O�?QO �?uOO"O4OnO�O�O �O�O_�O;_�O8_q_ _�_0_�_T_�_x_�_ �_�_7o"o[o�_oo �o>o�o�oto�o�o! �oE�o�o>�� �^�����A� �e� ���$���H�Z� l�����+�ƏO�� s��p���D�͟h�� �����ԟ�o�Z� ��.���R�ۯv�د� ��5�ЯY���}�c�u�8 1��*�<�v� ��߿��<�׿`��� ]ϖ�1Ϻ�U���y�� �ϯ�����\�G߀�� ��?���c����ߙ�"� ��F���j���)�c� ���������0��� -�f����%���I��� m������,P�� t�3��i� ��:���3 ��S�w /� �6/�Z/�~//�/ =/O/a/�/�/�/ ?�/ D?�/h??e?�?9?�? ]?�?�?
O�?�?�?O dOOO�O#O�OGO�OkO �O_�O*_�ON_�Or_ __1_k_�_�_�_�_ o�_8o�_5ono	o�o -o�oQo�ouo�o�o�o 4X�o|�; ��q����B� ���;�������[� ������>�ُb������!�������MA_SK 1 ��������ΗXNO � ݟ���MOT�E  ���S�_C�FG !Z����N�����PL_RA�NGV�N������O�WER "���Ϡ��SM_DRY�PRG %����%W��եTART� #Ǯ�UME_PRO���q����_EXEC_EN�B  ����GScPDJ�������gTDB����RMп���IA_OPTI�ON������~�NGVERS���`�řI_�AIRPUR�� �R�+���ÛMT_�֐T X���ΐO�BOT_ISOLEC����������/NAME8��H�Ě�OB_CATEG�ϣ,��S�[�.��ORD_NUM �?Ǩ��H705  N��ߨߺ�ΐPC_T�IMEOUT�� �xΐS232s�1�$��� L�TEACH PENDAN��o���)���V�T�M�aintenance ConsN��&�M�"B�P�No Use6�r�8�������̒��N�PO$��Ҏ�"�^��CH_LM�Q�朕	a�,�!U�D1:��.�RՐVgAILw��粥�*�SR  t�� ���5�R_INoTVAL����� ���V_DAT�A_GRP 2'|���� D��P�������	�� ����B0 RTf����� �/�/>/,/b/P/ �/t/�/�/�/�/�/? �/(??L?:?p?^?�? �?�?�?�?�?�?O O "O$O6OlOZO�O~O�O �O�O�O�O_�O2_ _ V_D_z_h_�_�_�_�_ �_�_�_o
o@o.oPo�vodo�o��$SA�F_DO_PUL�SW�[�S���i�SC�AN�������S�Cà(6��7���S�S�
������(q�q�qN� �L ^p���5��`� ��$��+�E�r2M�qqdY��P�`�J�	t/� @��������ʋ|���� r ք��_ @N�T ��'�9��K�X�T D�� X���������ɟ۟� ���#�5�G�Y�k�}��������䅎������Ǧ  "�;�oR� ����p"�
�u���Di���q$q�  � ���uq %�\�������ҿ��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6�H�Z����珈��� ����������g�;� D�V�h�z��������� ������(�Ӣ0�r� i�y���$�7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/?r�+?=? O?a?s?�?�?�?�?�? 8��?OO'O9OKO]O oO�O��$�r�O�O �O�O	__-_?_Q_c_ u_�_�Y�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o�o "4FXj|�c�路g������ �0�B�T�f�x�����@����ҏ�������:�Ҧ��y��3�	�	1234�5678��h!�B!�� \��p0���� Ο�����(�:�@� �c�u���������ϯ ����)�;�M�_� q�����R���ɿۿ� ���#�5�G�Y�k�}� �ϡϳ����ϖ���� �1�C�U�g�yߋߝ� ����������	��-� ��Q�c�u����� ��������)�;�M� _�q���B�������� ��%7I[m �������� !3EWi{� ������// //�S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?D/�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O*����O	_�E�?5_G_�Y_�yCz  A}��z   ��x�2�r }��)�
�W�/  	�*�2�O�_��_ oo"l�#\� �_hozo�o�o�o�o�o �o�o
.@Rd v����Mo�� ��*�<�N�`�r��� ������̏ޏ����&�8�J��X #P$P�Q:�R<u� k��Q?  �������S�P���Q�Qt C �PÙ۟�P(� `,b����]�P�Fl�$SCR_G�RP 1*7+�74� �� �,a ��U	 v��~������d����%���ɯ���h]���P�D1� �D7n��3��Fl�
CRX-10i�A/L 2345_67890�Pd�i r��Pd�L ��,a
1o�������-�[ ¶~�+fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@�R��d�t���H�~�Ă�m��ϴ��� ���ϼ��,a��1�P��U�[�G�imXhuP�,[��뾥B�  BƠߞҷԚ�9A�P��  @1`��暡@����� ?����H����ښ�F?@ F�`A�I� @�m�X��|����� ������������:�0%�7�I�[�B�i��� ��������������- Q<u`��En �ٯ���W�P�"+f@_�5��1`b���x����ͣ�O�,dA����ߒ��Fa�,a ��#!"/4/E-!pZ(f/x/G/ (�P�!(� �/�/�/��/�/?#9b����S7�س�M�ECLVLw  ,a��ݲ��Q@f1L_DE�FAULTn4b1��1`�3HOTSTR�=��2�MIPOWERF�m0pU�5�4WF�DO�6 �5L�E�RVENT 1+�u1u1�3 L!DUM_EIP#?�5H�j!AF_�INE�0SO,d!�FT)O�NIO�O!����O ��O�O!�RPC_MAI�N�O�H��O>_SV�IS_�I�-_�_!OPCUf�_�W�y_�_!TP&�PPU�_<Id�_"o�!
PMON_POROXY#o?Feo�no�R<o8Mf]o�o!�RDM_SRV�o<Ig�o!RȠ�"=Hh�oR!
�PM�o9LiA�!RLSYNC���y8��!R3OS(O��4�6��!
CE�PMTC�OM7�?Fk%���!=	K�CONS��>G�lq�Ώ!K�WA'SRC�o?Fm���;!K�USB�=H�n	�f�!STM�0��;JoU����O֟��c����CICE_�KL ?%K �(%SVCPR#G1��G�1�2G�L�"6�3o�t�6�4����"6�5��į6�6��6�7��6���W�R�	9_�d�3���6� 9���6�a�ܿ6���� 6���,�6�ٯT�6�� |�6�)���6�Q���6� y���^����^�ʿD� ^��l�^�ϔ�^�B� ��^�j���^����^� ��4�^���\�^�
߄� ��2���6��/��� �V��<�'�`�K��� o������������� &J5nY�� ������4 F1jU�y�� ���/�0//T/ ?/x/c/�/�/�/�/�/ �/�/??>?)?P?t?�_?�?
�_DEV �I�MC�:�84���4GRP 2/E�0+��bx 	� W
 ,@�0�?OD!OKODdOvO ]O�O�O�O�O�O�O�O _�O_N_5_r_Y_�_(�_/CE�0�_�_ �_o�_'ooKo]oDo �oho�o�o�o�o�o�o��o�o5Y�_D	�0i@���� ��� �=�$�a�s� Z���~��������؏�lD6OS�D�~�1O������ן
� ������U�<�y� `�������ӯ*��V � �	A�_:�ů^�E��� ��{�����ܿÿտ� ��6��Z�l�Sϐ�� 	A�q����%��Ϲ��� �υ��'߅�v�]ߚ� �߾��߷������*� 5�N��r����� ���������&�8�� \�C���g�y������� ����g�4-j Q�u����� B)fx_ ����)��/ ,//P/7/t/[/m/�/ �/�/�/�/?�/(??�L?^?E?�?�7d ��[~
�6 s��pA;*=�� 6?�=����D�>�����g�:�0��ī���|@�-��@�5_�e�A5�-�=BG+�h�&���6)�AB�m����`x��=�?7O�%TELEOP|8OcN[~y��5��o�ʾTF������������|��ҝ�����E�1��E@�*�A`��~�n�!�ǿ$�A���M��Y<T�������C=�J����Gc��M�cO��IJO/_�[~��6r _�1�<�׻��y�;��	A`����1bP��N	V�A��&@в@���@)E�]��1�����0���� x���Q���U?�Q���O�__ _oDU��NU9��6>����E�bQ��2]�j_ ���rAS�AT��@��@G�$�_ ��ywC� �Pr}��Q�� 2i?�R��_�o�_�_�oDU�K��5��l�������S���`�
�� 3>v��ĚM@�@��V�@�%@���Ŀ�q����]V�N��N�!�C(uµ��� �®�ɒow�o�o�DU��b�5?���T�@O�P��%�*�-���Ƒ�N�PA�����
Q@����q�A�����M�{�B&��br'C9�rt�1��^ѺfK��������pm�5>����@«��͙~��E�A������c�N'pA�(�AC8A�D����A��y�Nd�A���R��ֺ������s��`�_�^��\�n�S�BW��c�v"��?/����H?���4@� �+7�9��$ΏA8�	AAlܾc`�f�@�c+�N�e?6A�z2���LQ� f��t���`�D���2�D�)�DT�m���6M�W�1�������F0��<
u���8��NW`@�^}A1�Nu@X�ƿ�P�A%��N��j!��g(�E��uB��y�!F�`G�/������:�p��6
������\��w�������ku�f@�In_�PI�3�@K�@��"���P�������NuN�A���Q¸!C=�������º�����ٯ�п;�t�2�0�Bq̾���?P�������lG-���~�u�A�R��@&G A�z���:�A�X���NzQBA������V�������uC���׿�����ϒ���6 *����f�?#� ;����>b8�34�=+F':��V�?��r@���/>�@?[����n�MA���q����
]��@���3�xA?8m^�C߂���y�<���5�1*a��:�����2�  ������!�����OLp�A���� ����!�`������V�h�M�Ż���5���]��_?��A������+@��t�M?�<n@���@�o����[��A��
ޭ�@�C���/���=ؕ�{Ӎ� S�(�:��BU�I�IN��<�r�`���������%�'���ho��(L :p^������� ���$H6l ���\���� � //D/�k/�4/ �/�/�/�/�/�/�/? ^/C?�/?v?d?�?�? �?�?�?$?	OO�?�? �?<OrO`O�O�O�O�? �O O�O__$_&_8_ n_\_�_�O�_�O�_�_ �_o�_ o"o4ojo�_ �o�_Zo�o�o�o�o �oro�oi�oB� ������J/� n�b��r������� ����"��F�Џ:�(� ^�L�n���������ߟ ���� �6�$�Z�H� j���ҟ�������د ���2� �V���}��� F�h�B����Կ
��� .�p�Uϔ�ψ�vϘ� �Ϭ������H�-�l� ��`�N߄�rߔߖߨ� �� ��D���8�&�\� J��n�������� �����4�"�X�F�|� �����l���h��� ��0T��{��D ������, nS��t�� ���/F+/j� ^/L/�/p/�/�/�// �/?�/�/�/$?Z?H? ~?l?�?�/�??�?�? �?OO OVODOzO�? �O�?jO�O�O�O�O_ 
__R_�Oy_�OB_�_ �_�_�_�_�_oZ_�_ Qo�_*o�oro�o�o�o �o�o2oVo�oJ�o Z�n���
� .�"��F�4�V�|� j����Ǐ������ ��B�0�R�x����� ޏh�ҟ������� >���e�w�.�P�*��� ί�����X�=�|� �p�^�������ʿ�� �0��T�޿H�6�l� Z�|�~ϐ������,� �� ��D�2�h�V�x� ������ߞ������ 
�@�.�d�ߋ���T� ��P���������<� ~�c���,��������� ������V�;z� n\������ .R�F4jX �|������ �/B/0/f/T/�/� �/�z/�/�/�/�/? >?,?b?�/�?�/R?�? �?�?�?�?�?O:O|? aO�?*O�O�O�O�O�O �O�OBOhO9_xO_l_ Z_�_~_�_�_�__�_ >_�_2o�_BohoVo�o zo�o�_�oo�o
�o .>dR��o� �ox����*�� :�`�����P����� ޏ̏���&�h�M�_� �8��������ڟȟ ��@�%�d��X�F�h� j�|�����֯���<� Ư0��T�B�d�f�x� ���տ������,� �P�>�`϶�ܿ��� ���������(��L� ��s߲�<ߦ�8߶��� �� ���$�f�K��� ~�l���������� >�#�b���V�D�z�h� �����������:��� .R@vd��� ������* N<r���b� ����&//J/� q/�:/�/�/�/�/�/ �/�/"?d/I?�/?|? j?�?�?�?�?�?*?P? !O`?�?TOBOxOfO�O �O�OO�O&O�O_�O *_P_>_t_b_�_�O�_ �O�_�_�_oo&oLo :opo�_�o�_`o�o�o �o�o "H�oo �o8������ �P5�G�� ��h� �������(��L� ֏@�.�P�R�d����� �� ��$�����<� *�L�N�`���؟���� ���ޯ��8�&�H� ��į��ԯn�ȿ��� ڿ���4�v�[Ϛ�$� �� Ϟ��ϲ������ N�3�r���f�Tߊ�x� ���߮���&��J��� >�,�b�P��t��� ����"����:�(� ^�L��������r��� n��� 6$Z�� ���J����� �2tY�"� z�����
/L 1/p�d/R/�/v/�/ �/�//8/	?H/�/<? *?`?N?�?r?�?�/�? ?�?O�?O8O&O\O JO�O�?�O�?pO�O�O �O�O_4_"_X_�O_ �OH_�_�_�_�_�_�_�
o0or_Wo�U�P��$SERV_MA_IL  �U�`���QvdOUTPU}T�h�P}@vdRV 20f;  �` (a\o<�ovdSAVE�l�i�TOP10 21��i d 6� s�P
6r _�P:p�a6 *�a2ohz��� ����
��.�@� R�d�v���������Џ ����*�<�N�`� r���������̟ޟ����&�8�iuYP��cFZN_CF�G 2e��c�T�a�e|�GRP� 23��q ,�B   AƠ�QD�;� BǠ� � B4�SRB{21�fHELL�C4ev�`�o��|/�>�%RSR>� ?�Q���u�����ҿ�� ����,��P�;�t��_Ϙϩ����  �¼����Ϸ͊���P�&�'�)ސW��2�Pd��|g��HK 15�� ,ߡ߫ߥ��� ������@�;�M�_� �������������~�OMM 6���?��FTOV_E�NB�d�au�OW_REG_UI_���bIMIOFWD�L*�7.�ɥ��WAIT\�`ٞ����`r���d��TIM��7����VA�`��>��_UNIT[�*vyLCy�TRY���uv`ME�8@���aw֑d ��9�� �����<��X�Pڠ6p`?�  ��o+=`VL�l�fMON_�ALIAS ?e.��`heGo�� ����/)/;/M/ �q/�/�/�/�/d/�/ �/??%?�/I?[?m? ?�?<?�?�?�?�?�? �?!O3OEOWOO{O�O �O�O�OnO�O�O__ /_�OS_e_w_�_�_F_ �_�_�_�_�_o+o=o Ooaoo�o�o�o�o�o xo�o'9�o] o��>���� ��#�5�G�Y�k�� ������ŏ׏����� �1�C��g�y����� H���ӟ���	���-� ?�Q�c�u� ������� ϯᯌ���)�;�� L�q�������R�˿ݿ ��Ͼ�7�I�[�m� �*ϣϵ������ϖ� �!�3�E���i�{ߍ� �߱�\��������� ��A�S�e�w��4�� ����������+�=� O���s���������f� ����'��K] o��>���� �#5GY}�����l�$S�MON_DEFP�ROG &����� �&*SYSTE�M*���REC�ALL ?}�� ( �}
xy�zrate 11� *.* vir�t:\tmpba�ck\V =>19�2.168.56�.1:16260� |!�/�/�/�,}|K'k-5400 j/�|/??1?�#tp?disc 0�/� ��/�/�?�?�?�%t�pconn 0 �T?f?x?	OO-O�'8�copy frs�:orderfil.datY,S?� ЃO�O�O�-/KBmdb:V/oO� {O__,0_�$3xKD:g!Y/��O� �O�_�_�_� 4KUaS_e_�%�_o#o 5oHOZO�O�O�o�o�o �Oao�O|o1D_ �_�_z_����_S e�_	��-�@oRo�o vo�������o�ok��o ��)�<N�r�� ������]����� %���J�\�� ����� ��ȏc��~��!�3� F�ٟ�|�������ğ U�g�����/�B�T� ݯx��ϛϭ���үm� ����+�>�P��t� �ߗߩ߼�ο_��� �'�:?L?�(���ߌ� ���C��2�/d�v�� �+�>�P���tυ��� ������i���' :�L���p���8 ��[m�#5H� Z����������a ��|//1/D�� z�/�/�/�S/e/� 	??-?@R�v�? �?�?��k?�OO )O</N/�/r/�O�O�O �/�/]O�/�O_%_�O J?\?�? _�_�_�_�?�c_�?~_o!o3oDP��$SNPX_AS�G 2:����Va� � b%�7o~o  �?�GfPARAM� ;Ve`a W�	lkP>TDP�>X�d� ���I`OFT_KB_CFG  CS�\eFcOPIN_S_IM  Vk�b�+=OYsI`RV�NORDY_DO�  �eukrQSTP_DSB~��b�>kSR �<Vi � & ?TELEO�e��{v>TW`I`TOP_?ON_ERRxGb~�PTN Ve�P��D:�RING_PRM'���rVCNT_GP� 2=Ve�ac`x 	���DP��я�����BgVD�RP 1>�i�`�Vq؏ 0�B�T�f�x������� ��ҟ�����,�>� e�b�t���������ί ���+�(�:�L�^� p���������ʿ��  ��$�6�H�Z�l�~� �Ϸϴ����������  �2�D�V�}�zߌߞ� ����������
��C� @�R�d�v����� ����	���*�<�N� `�r������������� ��&8J\n �������� "4[Xj|� ������!// 0/B/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?t?�?�?�?�?�?��?�?O�PRG_�COUNT�f�P�)IENBe�+EM�UC�dbO_UPD �1?�{T  
 ODR�O�O�O�O�O_ _A_<_N_`_�_�_�_ �_�_�_�_�_oo&o 8oao\ono�o�o�o�o �o�o�o�o94F X�|����� ����0�Y�T�f� x������������� �1�,�>�P�y�t��� ������Ο��	��� (�Q�L�^�p������� ���ܯ� �)�$�6� H�q�l�~�������ƿ ؿ���� �I�D�V��"L_INFO 1=@�E�@��	 yϽϨ������>�~?zN�>G�q<����� A�Y����[��2#�@�"�Nl��,�����` ?@ <�@���o� C���B���C�_���0C+�r�|��2��p߂�-@Y?SDEBUG:@�@��o�d�I��SP_�PASS:EB?~��LOG A��]�A  o�i��v�  �Ao�UD1:\��}���_MPC�ݚEk�}A&�� �AK�SAV B��IA����*�i�1�SV�B�TEM_TIM�E 1C���@� 0  �n��i�ԝ�*���MEMBK  �E�A�������7X|�@� Z�i����������h�Y9
�� ��@� `r������0�� �@ Rdv�����
Le�//(/:/L/ ^/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?��SKV�[�EAj��?�?��?���@x]2����?i�  0P o�^
:O.@R�O��O�O}N�� ��OBDp�O_'_89_-L2�Y_�_ �_�_�_�_o�U�_�_ �o'o9oKo]ooo�o �o�o�o�o�o�o�o�#5GYk_?T1�SVGUNSPD��� '����p2�MODE_LIMG D��Ҋt2�p�qE�݉uABU�I_DCS H}5���0�G�0��D���|-�X�>���*���� 
��e��"i���r�i������uEDIT �I��xSCRN �J���rS�G �K�.�(�0߅S�K_OPTIONp��^����_DI��?ENB  /�����BC2_GRP 2L����MPC�ʓ�|BCCeF/�N���� ����`�>�W�B� g���x�����կ���� ����S�>�w�b� ��������Ͽ���� �=�(�a�Lυϗ�Ň �϶�������v��
� /�U�@�yߧ��`�i� ���߰�����
���.� �>�@�R��v��� ��������*��N� <�r�`����������� ����̀4FX ��|j����� ��B0fT vx�����/ �,//</b/P/�/t/ �/�/�/�/�/�/�/(? ?L?d?v?�?�?�? 6?�?�?�?O O6OHO ZO(O~OlO�O�O�O�O �O�O�O __D_2_h_ V_�_z_�_�_�_�_�_ 
o�_.oo>o@oRo�o vo�ob?�o�o�o �o<*Lr`�� ������&�� 6�8�J���n�����ȏ ���ڏ��"��F�4� j�X���|�������� ֟��o$�6�T�f�x� ��������ү����� ��>�,�b�P���t� �������ο��(� �L�:�\ς�pϦϔ� �ϸ������� ��H� 6�l�"��ߖߴ����� V������2� �V�h� z�H���������� ����
�@�.�d�R��� v������������� *N<^`r� ������&8 �\Jl���� ����"//F/4/ V/X/j/�/�/�/�/�/ �/?�/?B?0?f?T? �?x?�?�?�?�?�?O �?,O�DOVOtO�O�O O�O�O�O�O�O_ V�4P�$TBCSG_GRP 2O U��  ��4Q 
 ?�  __q_[_�__�_ �_�_�_�_o%k8R?S�QF\d�H�Ta?4Q	 HA����#e>���>�$a�\#eAT��A WR�o�hdjma��G�?Lfg�bpܚo�n�ffhf�̑ͼb4P|j��o*}@���Rhf�ff>G�33pa#e<qB�o�+=xrRp�qUy�rt~��H�y rIpTv�pBȺt~	xf 	x(�;���f���N��`���ˏڋ����	�V3.00WR	�crxlڃ	�*��3R~t��H�H��� \�.�]�  cC.�����V8QJ2?SRF]��~��CFG T U�PQ SPܚ���r�ܟ1��1�W�e�	Pe���v� ����ӯ������� �Q�<�u�`������� ��Ϳ�޿��;�&� _�Jσ�nπϹϤ��� ����WRq@�0�B� ��u�`߅߫ߖ��ߺ� �����)�;�M��q� \������4Q _�� �O ���J�8�n�\� �������������� ��4"XFhj| ������ .TBxf��nO ����//>/,/ b/P/�/t/�/�/�/�/ �/�/�/?:?(?^?p? �?�?N?�?�?�?�?�? �? O6O$OZOHO~OlO �O�O�O�O�O�O�O _ _D_2_T_V_h_�_�_ �_�_�_�_
o�_o@o �Xojo|o&o�o�o�o �o�o�o*N` r�B����� ��&��6�\�J��� n�����ȏ��؏ڏ� "��F�4�j�X���|� ��ğ���֟���0� �@�B�T���x����� ү䯎o���̯ʯP� >�t�b����������� ���Կ&�L�:�p� ^ϔϦϸ��τ����� � �"�H�6�l�Zߐ� ~ߴߢ���������� 2� �V�D�z�h��� �����������
�,� .�@�v�������\� ������<*` N����x�� �8J\( �������� /4/"/X/F/|/j/�/ �/�/�/�/�/�/?? B?0?f?T?v?�?�?�? �?�?�?OO��2ODO �� O�OtO�O�O�O�O �O_�O(_:_L_
__ �_p_�_�_�_�_�_ o �_$oo4o6oHo~olo �o�o�o�o�o�o�o  D2hV�z� ����
��.�� R�@�b���v���&OXO ֏菒�����N�<� r�`�������̟ޟ� ����$�&�8�n��� ����^�ȯ���گ� �� �"�4�j�X���|� ����ֿĿ����0� �T�B�x�fψϊϜ� ����������>�P� ��h�zߌ�6߼ߪ��� �������:�(�^�p� ���R������� ����  &�*� �*�>�*��$TB�JOP_GRP �2U����  ?���KC*�	V�]�Wd������X  *���� �, � ���*� �@&�?��	 �A������C�  �DD�����>v�>�\? ��a�G�:�o��;ߴAT������A�<��MX�����>��\)?;���8Q�����L��>�0 &�;�iG.��Ap�< � F�A�ff��v��� ):VM�.�� S>�o*�@��R�Cр	��������ff�:�6�/�?�33�B   ��/������>):�S����� �/�/@��H�%&/�/�z�=� <#�
*���v�;/�ڪ!?���4B�3?'? 2	��2?hZ?D?R?�? �?�?F?�?�?�?�?O AOO�?`OzOdOrO�O,�O*�C�*���A��	V3.00{��crxl��*�P��%�%c5Z �F� JZH� F6� F^� F�� F�f� F� G�� G5 G<
� G^] G�� G���G�*��G�S G�;o G��ERDu��\E[� E�� F( F-�� FU` F} � F�N F�� F�� Fͺ� F� F�V� G� Gz� Ga 9ѷI�Q�LHefJ4�o,b*�0c1����OH�ED_TCH� Xd�+X2S�2&�&�d$'X�o��o*�1F�TES�TPARS  ���cV�HRpAB�LE 1Yd� AN`*�����g$j
�g�h�h)�1��g	�h
�h�hHu*�U�h�h�h%v'RDI0n�GY k}��u	�O�#�@-�?�Q�c�u�)rS�l� �z6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z���I� ��m�Fwͩ��ȏڏ 쏘�����x)r~��NUM  ��n���2� �Ep�)r_CFG �Z��I���@V�IMEBF_TTqtD��e޶VER������޳R 1[�8{ 8�o*�d%�Q� ��د  9� K�]�oρϓϥϷ��� �������#�5�G�Y� k�}��ߡ߳������� ����1���E�W�i� {������������ ��/�A�S�e�w��� �������������+=O�_���@���`LIF M\��D`�����DR�(FP
�:!p�!p� d� ��MI_CHAN�� � DBGL�VL��fET�HERAD ?u��0`1�_}��ROUT��!�j!��SNMASKY�j255.%S/�//A/S�`OOLO_FS_DIp��CORQCTRL� ]8{��1o�-T �/�/�/??+?=?O? a?s?�?�?�?�?�?�? �?OL�/6O%OZOc�PE_DETAI�7�*PGL_CONFIG c�������/cel�l/$CID$/grp1^O�O�O�O
__|���G_Y_k_ }_�_�_0_�_�_�_�_ oo�_CoUogoyo�o �o,o>o�o�o�o	 -�oQcu��� :�����)�� �_�q���������׮}N����%�7�I�a�KOq�P��M����� ʟܟ� �G�$�6�H� Z�l�~������Ưد ������2�D�V�h� z������¿Կ��� 
ϙ�.�@�R�d�vψ� ��)Ͼ��������� ��<�N�`�r߄ߖ�%� ����������&�� J�\�n����3��� �������"���F�X��j�|��������@��User Vi�ew �I}}12�34567890 ����+=Ex ,�e����2��B� �����`r��3�Oas����x4>//�'/9/K/]/�~/x5 ��/�/�/�/�/?p/2?x6�/k?}?�?�? �?�?$?�?x7Z?O 1OCOUOgOyO�?�Ox8O�O�O�O	__-_��ON_TR lCamera�� �O�_�_�_�_�_�_˂E�_o)o;n��Uogo`yo�o�o�o�)  mV �	�_�o#5GY  o}���o������F_�mV=� k�}�������ŏl� ���X�1�C�U�g�y� ��2�D��"�ן��� ��1�؏U�g�y�ğ ������ӯ�����D� �k��E�W�i�{����� F�ÿտ�2���/� A�S�e��nUY9���� ��������	߰�-�?� Qߜ�u߇ߙ߽߫��� v�D�If��-�?�Q� c�u�ߙ������ ����)�;���D��I ��������������� )t�M_q���N�`�93�� 0B��Sx� 1�����//
�J	oU0�U/g/y/ �/�/�/V�/�/�/� ?-???Q?c?u?/./ tPv[?�?�?�?OO (O�/LO^OpO�?�O�O �O�O�O�O�?oU�k�O :_L_^_p_�_�_;O�_ �_�_'_ oo$o6oHo Zo_;%N��_�o�o�o �o�o �_$6H�o l~����moe ��]�$�6�H�Z�l� �������؏��� � �2��e&�ɏ~� ������Ɵ؟����  �k�D�V�h�z����� E�e��5����� � 2�D��h�z���ׯ���¿Կ���
ϱ�  ��9�K�]�oρπ�ϥϷ���������   ��5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u����� ����������)�;M_q�  
���(  �-�( 	 ���� ���#35G@}k����
� �Y�
//./�� R/d/v/�/�/�/��� �/�/�/A/?0?B?T? f?x?�/�?�?�??�? �?OO,O>O�?bOtO �O�?�O�O�O�O�O_ KO]O:_L_^_�O�_�_ �_�_�_�_#_ oo$o k_HoZolo~o�o�o�_ �o�o�o1o 2D Vh�o�o���	 ��
��.�@��d� v��������Џ�� �M�*�<�N���r��� ������̟�%��� &�m�J�\�n������� �ȯگ�3��"�4� F�X�j����������� ֿ�����0�w��� f�xϊ�ѿ�������� ���O�,�>�Pߗ�t� �ߘߪ߼������� �]�:�L�^�p����߻@ ������������ ��"�frh:\tpg�l\robots�\crx!�10ia_l.xml�� D�V�h�z�������������������0 BTfx���� �����,>P bt������ ��/(/:/L/^/p/ �/�/�/�/�/�/��/ ?$?6?H?Z?l?~?�? �?�?�?�?�/�?O O 2ODOVOhOzO�O�O�O �O�O�?�O
__._@_ R_d_v_�_�_�_�_�_ �O�_oo*o<oNo`o ro�o�o�o�o�o�n ��6� ���<�< 	� ?� �k!�o;iOq �������� �%�S�9�k���o���裏я����(�$�TPGL_OUT?PUT f����w�� � &�8�J�\�n������� ��ȟڟ����"�4� F�X�j�|�������į��p�ր2345?678901��� ��1�C�K����r� ��������̿d�п� �&�8�J��}T�|� �Ϡϲ���\�n���� �0�B�T���bߊߜ� ������j�����,� >�P����߆���� ����x����(�:�L� ^���l����������� t���$6HZl z������ � 2DVh  �������/ ./@/R/d/v//�/�/��/�/�/�/�/ۂ $$��ί<7*? \?N?�?r?�?�?�?�? �?�?OO4O&OXOJO |OnO�O�O�O�O�O�O _�O0_"_T_}�an_@�_�_�_�_�_�]@��_o	z ( 	 V_Do2ohoVo�o zo�o�o�o�o�o
�o .R@vd�� �������(��*�<�r�`���ܦ� ? <<I_ˏ ݏ�������:�L� ֪��}���)���ş�� �����k��C�ݟ/� y���e���������� ���-�?��c�u�ӯ ]�����W���Ϳ�� )χ���_�q��yϧ� �ϓ�����M��%߿� �[�5�Gߑߣ�߫� ��s����!���E�W� ��?���9������ ���i���A�S���w� ��c�u����/��� ��=)s��� ��U���' 9�!o	[�� ���K�#/5/� Y/k/E/w/�/�/�/ �/�/�/?�/?U?g? �/�?�?7?�?�?�?�?�	OO��)WGL�1.XML�_PM��$TPOFF_L�IM ���P����^FN_SV�f@  �TxJP_MON g��SzD�P�P2ZI�STRTCHK �h��xFk_aBVTCOMPAT�H�Q|FVWVAR �i�M:X�D ��O R_�P�B�bA_DEFPRO�G %�I%?TELEOPi_�O�_DISPLAY�m@�N�RINST_�MSK  �\ ��ZINUSER�_�TLCKl�[QUICKMEN:o��TSCREY`���Rtpsc@�Tat`yixB�`_�i�STZxIRACE_CFG j�I�:T�@	[T
?���hHNL 2k�Z���aA[ gR-? Qcu����z�eITEM 2l{� �%$1234567890 ��  =<
�0�B�J�  !P�X�dP���[S���"�� �X�
�|���W���r� ֏����.��0�B�\� f�����6�\�n�ҟ�� ������>���"� ��.�����ίR���� Ŀֿ:��^�p�9ϔ� Tϸ�xϊ���d� ��H��l��>�Pߴ� \�������v� ����� �h�(�ߞ߰�4�L� �ߦ�����@�R�� v�6���Z�l������ ���*���N��� �� ����������X� ��J
n�� �b����"4 F�/|</N/�Z/ ���//�/0/�/? f/?�/�/e?�/�?�/ �?�?�?,?�?P?b?t? �?�?DOjO|O�?�OO O(O�O�O^O_0_�O <_�O�O�_�O�__�_��_H_�_l_~_Go�dS��bm�oLj�  �rLj �a�o�Y
 �o�o�o�o{j�UD1:\|���^aR_GRP �1n�{� 	 @�PRd{N� r����~��p����q+��O�:�?�  j�|�f����� �����ҏ����>� ,�b�P���t����������	e���\cS�CB 2ohk U�R�d�v��������Я�RlUTOR?IAL phk�o�-�WgV_CONFIG qhm�a�o��o��<�OUTPU�T rhi}�����ܿ� ��$� 6�H�Z�l�~ϐϢϴ� z�ɿ���� ��$�6� H�Z�l�~ߐߢߴ��� ������� �2�D�V� h�z���������� ��
��.�@�R�d�v� �������������� *<N`r�� ������& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/� �/�/??0?B?T?f? x?�?�?�?�?�/�?�? OO,O>OPObOtO�O �O�O�O�?�O�O__ (_:_L_^_p_�_�_�_ �_�_f�x�ǿoo,o >oPoboto�o�o�o�o �o�o�O(:L ^p������ �o ��$�6�H�Z�l� ~�������Ə؏�� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я����*�<� N�`�r���������̿ ޿���&�8�J�\� nπϒϤ϶������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ������������,� >�P�b�t�����������������X���#��N�_r ������� &8J��n�� ������/"/ 4/F/X/i|/�/�/�/ �/�/�/�/??0?B? T?e/x?�?�?�?�?�? �?�?OO,O>OPOa? tO�O�O�O�O�O�O�O __(_:_L_^_oO�_ �_�_�_�_�_�_ oo $o6oHoZok_~o�o�o �o�o�o�o�o 2 DVgoz���� ���
��.�@�R� d�u��������Џ� ���*�<�N�`�q� ��������̟ޟ����&�8�J�\�k��$�TX_SCREE�N 1s%; �}�k��� ��ӯ���	���Z ��I�[�m������� ,�ٿ����!�3Ϫ� W�ο{ύϟϱ����� L���p��/�A�S�e� w��� ߭߿������� �~�+��O�a�s�� ��� ���D����� '�9�K���������� ������R���v�#5�GYk}����$�UALRM_MS�G ?����� �n���	: -^Qc������� /�SEV � �2&�E�CFG u�����  n�@��  Ab!   B�n�
 /u��� �/�/�/�/�/�/??�%?7?I?W7>!GRPw 2vH+ 0n��	 /�?� I_�BBL_NOTE� wH*T���lu���w��T �2DEFPROz� %� (%��Ow�	OBO-BTELEOPGO#O�O�O �O�O�O�O�O_�O&_��?�0FKEYDA�TA 1x���0'p W'n��?�_`�_z_�_�_�Z,(�_�on�(POIN	To>o �_coJo�o�no�o�o dTOUCHU`O�o�o�o 7[mT�x� �����!��E���Z��/frh�/gui/whi�tehome.pngQ�������ŏ׏��h�point z���/�A�S��\� ��������ȟڟi��� �"�4�F�X��|��������į֯e�h�t?ouchup����/�A�S�e��h�arwrg������ÿ տ�n���/�A�S� e����ϛϭϿ����� �τ��+�=�O�a�s� ߗߩ߻������߀� �'�9�K�]�o��� ������������#� 5�G�Y�k�}�T���� ���������1C Ugy���� ��	�?Qc u��(���� //�;/M/_/q/�/ �/�/6/�/�/�/?? %?�/I?[?m??�?�? 2?�?�?�?�?O!O3O �?WOiO{O�O�O�O@O �O�O�O__/_�OS_ e_w_�_�_�_�_N_�_ �_oo+o=o�_aoso��o�o�o�oV��k}�b�����o@}�o8J$v,6� {.������� ��/��S�:�w��� p�����я�ʏ�� +��O�a�H���l��� ����ߟ���'�9� Ho]�o���������ɯ X�����#�5�G�֯ k�}�������ſT�� ����1�C�U��y� �ϝϯ�����b���	� �-�?�Q���u߇ߙ� �߽�����p���)� ;�M�_��߃���� ����l���%�7�I� [�m������������ ��z�!3EWi ��������� П/ASew~ ������/� +/=/O/a/s/�//�/ �/�/�/�/?�/'?9? K?]?o?�?�?"?�?�? �?�?�?O�?5OGOYO kO}O�OO�O�O�O�O �O__�OC_U_g_y_ �_�_,_�_�_�_�_	o o�_?oQocouo�o�o �o:o�o�o�o) �oM_q���6 �����%�7��9�����b�t���^�������,��돞����3� E�,�i�P�������ß ���������A�S� :�w�^�������ѯ�� ��ܯ�+�
O�a�s� �������Ϳ߿�� �'�9�ȿ]�oρϓ� �Ϸ�F��������#� 5���Y�k�}ߏߡ߳� ��T�������1�C� ��g�y������P� ����	��-�?�Q��� u�����������^��� );M��q� �����l %7I[��� ���h�/!/3/ E/W/i/@��/�/�/�/ �/�/�??/?A?S? e?w??�?�?�?�?�? �?�?O+O=OOOaOsO O�O�O�O�O�O�O_ �O'_9_K_]_o_�__ �_�_�_�_�_�_�_#o 5oGoYoko}o�oo�o �o�o�o�o�o1C Ugy���� ��	���?�Q�c� u�����(���Ϗ�� ����;�M�_�q���h����~ ���~ ���ҟ���Ο�*��,�[�� �f�������ٯ���� ���3��W�i�P��� t���ÿ���ο�� /�A�(�e�Lωϛ�z/ ����������(�=� O�a�s߅ߗߩ�8��� ������'��K�]� o����4������� ���#�5���Y�k�}� ������B������� 1��Ugy�� ��P��	- ?�cu���� L��//)/;/M/ �q/�/�/�/�/�/Z/ �/??%?7?I?�/m? ?�?�?�?�?�?���? O!O3OEOWO^?{O�O �O�O�O�O�OvO__ /_A_S_e_�O�_�_�_ �_�_�_r_oo+o=o Ooaosoo�o�o�o�o �o�o�o'9K] o�o������ ��#�5�G�Y�k�}� �����ŏ׏����� �1�C�U�g�y���� ����ӟ���	���-� ?�Q�c�u��������@ϯ�����0����0����B�T�f�>�����t�, ��˿~��ֿ�%�� I�0�m��fϣϊ��� ��������!�3��W� >�{�bߟ߱ߘ��߼� ����?/�A�S�e�w� ����������� ���=�O�a�s����� &����������� 9K]o���4 ����#�G Yk}��0�� ��//1/�U/g/ y/�/�/�/>/�/�/�/ 	??-?�/Q?c?u?�? �?�?�?L?�?�?OO )O;O�?_OqO�O�O�O �OHO�O�O__%_7_ I_ �m__�_�_�_�_ �O�_�_o!o3oEoWo �_{o�o�o�o�o�odo �o/AS�ow ������r� �+�=�O�a������ ����͏ߏn���'� 9�K�]�o��������� ɟ۟�|��#�5�G� Y�k���������ůׯ ������1�C�U�g� y��������ӿ��� ���-�?�Q�c�uχ��^P���^P��������ͮ���
���,��;���_�F� �ߕ�|߹ߠ������� ���7�I�0�m�T�� �����������!� �E�,�i�{�Z_���� ���������/A Sew���� ���+=Oa s������ //�9/K/]/o/�/ �/"/�/�/�/�/�/? �/5?G?Y?k?}?�?�? 0?�?�?�?�?OO�? COUOgOyO�O�O,O�O �O�O�O	__-_�OQ_ c_u_�_�_�_:_�_�_ �_oo)o�_Mo_oqo �o�o�o�o���o�o %7>o[m� ���V���!� 3�E��i�{������� ÏR������/�A� S��w���������џ `�����+�=�O�ޟ s���������ͯ߯n� ��'�9�K�]�쯁� ������ɿۿj���� #�5�G�Y�k����ϡ� ��������x���1� C�U�g��ϋߝ߯�����������`���>�`���"�4� F��h�z�T�,f��� ^���������)�� M�_�F���j������� ������7[ B�x���� �o!3EWix� �������� ///A/S/e/w//�/ �/�/�/�/�/�/?+? =?O?a?s?�??�?�? �?�?�?O�?'O9OKO ]OoO�OO�O�O�O�O �O�O_�O5_G_Y_k_ }_�__�_�_�_�_�_ o�_1oCoUogoyo�o �o,o�o�o�o�o	 �o?Qcu��( ������)�  M�_�q��������ˏ ݏ���%�7�Ə[� m��������D�ٟ� ���!�3�W�i�{� ������ïR����� �/�A�Яe�w����� ����N������+� =�O�޿sυϗϩϻ� ��\�����'�9�K� ��o߁ߓߥ߷����� j����#�5�G�Y��� }��������f�����1�C�U�g�>��i��>������������������,��?&cu \������� )M4q�j �����/�%/ /I/[/:�/�/�/�/ �/�/���/?!?3?E? W?i?�/�?�?�?�?�? �?v?OO/OAOSOeO �?�O�O�O�O�O�O�O �O_+_=_O_a_s__ �_�_�_�_�_�_�_o 'o9oKo]ooo�oo�o �o�o�o�o�o�o#5 GYk}��� �����1�C�U� g�y��������ӏ� ��	���-�?�Q�c�u� ����p/��ϟ��� ��;�M�_�q����� ��6�˯ݯ���%� ��I�[�m������2� ǿٿ����!�3�¿ W�i�{ύϟϱ�@��� ������/߾�S�e� w߉ߛ߭߿�N����� ��+�=���a�s�� ����J������� '�9�K���o������� ����X�����#5 G��k}���������������&�HZ4,F/�>/� ����	/�-/?/ &/c/J/�/�/�/�/�/ �/�/�/?�/;?"?_? q?X?�?|?�?�?���? OO%O7OIOXmOO �O�O�O�O�OhO�O_ !_3_E_W_�O{_�_�_ �_�_�_d_�_oo/o AoSoeo�_�o�o�o�o �o�oro+=O a�o������ ���'�9�K�]�o� �������ɏۏ�|� �#�5�G�Y�k�}�� ����şן������ 1�C�U�g�y������ ��ӯ���	��?-�?� Q�c�u���������Ͽ ���Ϧ�;�M�_� qσϕ�$Ϲ������� �ߢ�7�I�[�m�� �ߣ�2���������� !��E�W�i�{��� .�����������/� ��S�e�w�������<� ������+��O as����J� �'9�]o ����F����/#/5/G/�$UI�_INUSER � ���h!��  �H/L/_MENHI�ST 1yh%�  ( �u ��+/SO�FTPART/G�ENLINK?c�urrent=e�ditpage,�TELEOP,1 �/�/?!?�)�/�%�menu�"113�3�/}?�?�?�? �'E?W>71l?�?O�#O5O�(�?W?54 �?�O�O�O�OIO[OmB k?__+_=_�?�O�!2�O�_�_�_�_�Oa_c348,2�_o$o6oHo��Iono�o�o�o�o�o��\a�!\o �o/ASVow �����`�� �+�=�O������� ����͏ߏn���'� 9�K�]�쏁������� ɟ۟j�|��#�5�G� Y�k���������ůׯ ��o�o�1�C�U�g� y�|�������ӿ��� ���-�?�Q�c�uχ� ϫϽ�������ߔ� )�;�M�_�q߃�ߧ� �����������7� I�[�m��� ���� ����������E�W� i�{������������� ����ASew ���<��� +�Oas�� �8���//'/ 9/�]/o/�/�/�/�/ F/�/�/�/?#?5? � 2�k?}?�?�?�?�?�/ �?�?OO1OCO�?�? yO�O�O�O�O�ObO�O 	__-_?_Q_�Ou_�_ �_�_�_�_^_p_oo )o;oMo_o�_�o�o�o �o�o�olo%7�I[F?��$UI�_PANEDAT�A 1{�����q  	��}  frh�/cgtp/fl�exdev.st�m?_width�=0&_heig�ht=10�p�pi�ce=TP&_l�ines=15&�_columns�=4�pfont=�24&_page?=whole�pm~I6)  rim�9�  �pP�b�t��� ���������Ǐ�� (�:�!�^�E�����{������ܟ�՟�I6� �  [0 �J�O�a� s���������ͯ@�� ��'�9�K���o��� h�����ɿۿ¿��� #�5��Y�@�}Ϗ�v���&��Ɠs���� �)�;�Mߠ�q�䯕� �߹�������V��%� �I�0�m��f��� ���������!��E� W����ύ��������� ��:�~�/ASe w������  =$asZ �~����d�v� '/9/K/]/o/�/��/ �/*�/�/�/?#?5? �/Y?@?}?�?v?�?�? �?�?�?O�?1OCO*O gONO�O�/�/�O�O �O	__-_�OQ_�/u_ �_�_�_�_�_6_�_o �_)ooMo_oFo�ojo �o�o�o�o�o�o% 7�O�Om��� ��^_�!�3�E� W�i�{������Ï�� �������A�S�:� w�^�������џDV ��+�=�O�a����� ��
���ͯ߯��� |�9� �]�o�V���z� ��ɿ���Կ�#�
�`G�.�k�ޟ�}�|�@�����������)�� 4ߧ�#�`�r߄ߖߨ� ��!����������8� �\�C���y������������������$UI_POST�YPE  ���� 	 ��s�B�QUICK�MEN  Q��`�v�D�RESTO�RE 1|���  �������������m ASew�,� �����+= Oan��� ��//�9/K/]/ o/�/�/6/�/�/�/�/ �/�??0?�/k?}? �?�?�?V?�?�?�?O O�?COUOgOyO�O6? @O�O�O.O�O	__-_ ?_Q_�Ou_�_�_�_�_ `_�_�_oo)o�O6o HoZo�_�o�o�o�o�o �o%7I[�o�������SC�RE��?���u1sc��uU2�3�4�5��6�7�8��sT;ATM�� ����:�USER�p��r�T�p�ks���4���5��6��7��8���B�NDO_CFG }Q�����B��PDE����None��v�_INFO 2~��5)���0%�D� ��2�s�V�������͟ ߟ��'�9��]��o�R���z��OFF?SET �Q�-���hs��p���� �G�>�P�}�t���Я ��׿ο����C� :�L�^Ϩ����͘����
����av��WO_RK �!������.�@ߢ�u�UFR?AME  ����RTOL_AB�RT�����ENB��ߣ�GRP 1������Cz  A������*�<�@N�`�r��֐�U������MSK  h�)���N��%!���%z����_EV�N�����+�ׂ3݄«
 h��UEV��!td�:\event_�user\�u�C�7z���jpF��n�S�Ps�x�spot�weld��!CA6��������!� ��G|'��5kY �����>� ��1�Ug� ��/��	/^/M/ �/-/?/�/c/�/�/�/��/$?�/H?�/:J�Wf�3�����8C?�?�? �?�?�?�?O +OOOOaO<O�O�OrO �O�O�O�O_�O'_9_�_]_o_J_�_�_�_��$VALD_CP�C 2�« q�_�_� w� �qd�R�*o_oqo��hsNbd�j�`��i�d a{�oav�_�ooo3 BoWi{�o�o�o�o ��o�PA�0� e�w������� ���(�=�L�a�s� 
�������ʏ���� �$�ޟH�:�o����� ����ڟ؟����� � 2�G�V�k�}������� ¯ԯ�����.�� R�S�yϋϚ������ ����	��*�<�Q�`� u߇ߖϨϺ������� ��&�8�M�\�q�� ��߶���n������ "�4�F�[�j������ �����������!0� B�Wf�{������ �����,>t eT������ �/+/:La/p �/�/./�����/ /'?6/H/?l/^?�? �?�/�/�/�/�/?#O �?D?V?kOz?�O�O�? �?�?�?�?_O1_@O RO9_vOw_�_�_�O�O �O_�__-o<_N_`_ uo�_�o�o�_�_�_�_ o&o;Jo\oq�o ����o�o�o� � "7�FXj���� �������!�0� E�T�f�{�������ß ҏ����
�,�A�P� b�����x�����Ο�� ���(�*�O�^�p� ��������R�ܯ� � �Ϳ6�K�Z�l�&ϐ� �Ϸ���ؿ���"� � 2�G���h�zϏߞϳ� ��������
��1�@� U�d�v�]�ߛ����� �����,��<�Q�`� r������������ ��&�;J�_n��� ���������� �$F[j|�� �����0 E/Ti/x��/��/ �/�/�//,/.?P/ e?t/�/�/�?�?�?�? �/??(?:?L?NOsO �?�?�O�?�O�OvO O O$O6O�OZOo_~O�O J_�O�_�_�_�O_ _�F_D_V[�$VAR�S_CONFIG� ��Pxa  FP]S��\lCMR_G�RP 2�xk� ha	`�`  �%1: SC130EF2 *�o$�`]T�VU�P�h`�5_Pa?� W A@%pp*`�Vn' No9xCVX�dv��a��<uSA�%p�q�_R���_R B���#�_Q'��H��l� ;���{�����؏ÏՏ �e��D�/�A�z�-������ddIA_WO_RK �xeܐy�Pf,		�Q�xe���G�P ����YǑRTSYNCSET  xi��xa-�WINUR�L ?=�`� ����������ȯگ�SIONTMOUt9�]Sd� ���_CFG �S�۳�S۵P��` FR:\~��\DATA\�� �� MC�3�LOG@�   oUD13�EXd��_Q' B@ ����x�e_ſx��ɿ�VW � �n6  ����VV��l�q  =���?�]T<�y�}Y�TRAIN��l�N� 
gp?ňCȞ��TK���b�xk (g�����_� ��������U�C�y� g߁ߋߝ߯�������_GE��xk�`_P�
�P�Rꋰ�RE��xe*�`hL�EX�xl`1-�e�VMPHASOE  xec��ecRTD_FIL�TER 2�xk �u�0���� 0�B�T�f�x�����VW �������� $6�HZl_iSHIF�TMENU 1�^xk
 <�\%��������� �=&sJ\� ������'/��	LIVE/S�NA�c%vsf�liv��9/���� 7�U�`\"menur/w//�/�/��d���]��MO�e�y��5`h`ZD4ɘV�_Q<��0��$�WAITDINE�ND��a2p6OK�  �i�<���?Sܺ?�9TIM�����<Gw?M�?*K�?�
J�?
J�?�8RELE��:G6p3���r1_ACTO 9Hܑ�8�_<� �ԙ�%��/:_af�BRDIS��`�N�$XVR���y��$ZA�BC�b1�S; ),��j�I�2B_Zm�I1�@VSPT q�y��eG�
�*��/o�*!o7o�WD�CSCHG �pԛ(��P\g@�P[IPL2�S?i���o�o�o�ZMPCF�_G 1��ii�0@'¯S;Ms�S��i��p'��g��e2���  ?5����3|Y=�y��2�/�6��B��65=����6
*�~��`C��B��_�C�_�I�1�q�>�����F��=5�[����濢c����������Z�~���Ï�>���0C+�r�|�G2��ڏ�ӈ��� ��*�@�N�x��$�6�H�0N�`��Tp����o�_CYLI�ND�� { ���� ,(  * =�N�G�:�w�^����� ��ѯ���7�� ��<�#�5�r������� ����޿y�_����8�@ύ�nπ�㜻ã wQ �5�����S �����(�ٻ�X���r�A��SPH�ERE 2��� ҿ��"ϧ������P� c�>�P�̿t���ߪ� �����'���]�o� L���p�W�i�������������PZZ�F � 6