��   v��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@���&�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	>4SUSRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  wXKaIRTs1�	o`'2 L1���L2�R�	 %,��?���b1`��c�c~a����?�  �o��
 ��a�o�o1CU �oz� ����c�
�� .�@�R��v������� ��Џ�q���*�<� N�`��������̟ ޟm���&�8�J�\� n���������ȯگ� {��"�4�F�X�j��� ������Ŀֿ���`TPTX���ʊ�)�� s ��Ƅ�$/so�ftpart/g�enlink?h�elp=/md/�tpmenu.d�g���ϨϺ��υ�&a�s�pwd���+� =�O߄�s߅ߗߩ߻� ��\�����'�9�K� ���߁��������V���a�f�oC ($p�-����T�?�x���a�a��oŪ����l��c�gH���a�ah���a�h��h�	f���%�������`����`  ���f eOp��h#h��F�bc Xc�B 1�)hR \��`_�� ;REG VED]����wholem�od.htm�	s�ingl	do�ub tri�p8browsQ�����u ���//@/��|�dev.s�l�/3� 1�,	t �/_�/;/i/??/?��/S?e?w?�?�?�?� ��?�?OO%O�7OIO[OmOO�E @ �?�O�O�O�O�O_�F �	�?�?;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omooM'�o �o�o�o�o�o+ =Oas���� �����?>�P�b� t���������Ώ���O �����L�^�_'_ �������ş���� �6�1�C�U�~�y��� ��Ư��ӯ�o��� -�?�Q�c�u������� ��Ͽ����)�;� M�_�-��ϬϾ����� ����*�<�7�`�r� A�Sߨߺ�q���i�� ���!�J�E�W�i�� ������������"� �/���O�I�w����� ����������+ =Oas���� ���,>Pb t���߼��� //�����^/Y/k/ }/�/�/�/�/�/�/�/ ?6?1?C?U?~?y?�? Y��?�?�?�?�?	OO -O?OQOcOuO�O�O�O �O�O�O�O__�R_ d_v_�_�_�_�_�_�_ �_�o*o�_o`oro��j�$UI_TO�PMENU 1�K`�aR� 
d�a*Q)�*default�5_]*lev�el0 * [	 #�o�0�o�'rtpio[23�]�8tpst[1[x)w9�o	�=�h58E01_�l.png��6menu5�y�p�C13�z��z	�4���q��]������� ��̏ޏ)Rr���+��=�O�a���pri�m=�page,?1422,1h��� ��şן����1��C�U�g���|�class,5p������ɯۯ�����13���*�<�N�`�r���|�53������ҿ�����|�8��1�C� U�g�y����ϯ���������"Y�`�a�o/߀�m!ηq�Y�w�avt�yl}Tfqmf[0�nl�	��c[164[w��59[x�qG���/��29��o�%� 1���{��m��!��� ��0�B���f�x��� ������O�����,>����2P�� ���\��' 9K������������1��/$/�6/H/Z/��|�ainedi'ߑ/�/�/��/�/��conf�ig=singl�e&|�wintp ���/$?6?H?Z?	��8�??ٷ�gl[�<��?�߲08��
A���?,OH2��DO�?cO��O�z �� �4s�x�O�O�$��Ol� E_W_i_{_�_�_���_ �_�_�_oo/o�_So@eowo�o�o�o�$;�$�doub5o��1}3��&dual�i38��,4�o&�o9�o�n�o�a8� ��Ao����&� 8��\�n��������� m�����
��.�@� K�d�v���������Z{?�;�M�sc�_;���s��X�}���e�u��0����O_� �J�p�^�6e�u7 �����ｿϿ��� P�)�;�M�_�qσ�� �Ϲ����������"�1�M�_�q߃� �ߠϹ��������� ��7�I�[�m���� ����������!�����6(�]�o��������$��74�������)�C�ߟT�	TPTX[20�=Aw24#GJ���Bw1H������8 �"H���A#��[��tv`�R��@24�K0�11����5S:�$treev'iew3�f3��o}?381,26M/ _/q/0�/�/�/�/�/ �/~/?%?7?I?[?m?�o/܈5�o5%���? �?�?
?#O5OGOYOkO�}O�?�? "2�?8"2@K��O�O_�O��1�?��E�f_x_�_ �6<_ڀedit�a>_ P_�_�_oˉ/���_ �Cooo�o�oB�o�o ��oA�o�+ =Oas��o�� �����(�9��� Q�x���������ҏO ����,�>�P�ߏt� ��������Ο]���� �(�:�L�^�ퟂ��� ����ʯܯk� ��$� 6�H�Z��l������� ƿؿ�y�� �2�D� V�h����Ϟϰ����� �ϕo�o��o@ߧE� c�u߇ߙ߽߬����� O����)�<�M�_�q� ���W��������� &�8���\�n������� ��E�������"4 ��Xj|���� S��0B� fx����O� �//,/>/P/�t/ �/�/�/�/�/]/�/? ?(?:?L?��߂?1� �?���?�?�?�?O $O5OGO�?SO}O�O�O �O�O�O�O�O��2_D_ V_h_z_�_�_�/�_�_ �_�_
oo�_@oRodo vo�o�o)o�o�o�o�o *�oN`r� ��7����� &��J�\�n������� ��E�ڏ����"�4� ÏX�j�|�������a? s?蟗?�sO_/�A� S�e�w���������� �����,�=�O�a� #_������ο��=� �(�:�L�^�pς�� �ϸ������� ߏ�$� 6�H�Z�l�~�ߐߴ� ����������2�D� V�h�z�������� ����
����@�R�d� v�����)����������ƚԔ*de�fault%��*level8��ٯw���? tpst[1]�	��y�tpioG[23���u����J\men�u7_l.png�_|13��5Ж{�y4�u6 ���//'/9/K/]/ ���/�/�/�/�/�/j/ �/?#?5?G?Y?k?�"�prim=|p�age,74,1�p?�?�?�?�?�?�"��6class,13�?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_f_x_{?�218�?�_�_ �_�_�__B6o9o�Ko]ooo�o`�$U�I_USERVI�EW 1֑֑�R 
����o��o�o[m �o'9K] � ����l��� #�5��oB�T�f���� ��ŏ׏鏌���1� C�U�g�
��������� ӟ~�����v�?�Q� c�u���*�����ϯ� 󯖯�)�;�M�_�
� �~������ݿ�� �%�ȿI�[�m�ϑ� 4ϵ��������Ϩ�
� �.ߠ�i�{ߍߟ߱� T���������/��� S�e�w���Fߨ�� ��>���+�=�O��� s���������^����� '����FX�� |������ #5GY�}�� ��p���h1/ C/U/g/y//�/�/�/ �/�/�/�/?-???Q? c?/p?�?�??�?�? �?OO�?;OMO_OqO �O&O�O�O�O�O�O�? �O_ _�OD_m__�_ �_�_X_�_�_�_o!o �_EoWoio{o�o0h