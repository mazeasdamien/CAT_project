��   ?Q�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����MN_MCR�_TABLE �  � $MA�CRO_NAME� %$PRO�G@EPT_IN�DEX  $OPEN_IDa�ASSIGN_T�YPD  qk$MON_NO}�PREV_SUB�y a $USER�_WORK���_�L� MS�*RT�N  �&S�OP_T  �� $�EMG�O��RESE�T�MOT|�H�OLl�� 2��STAR PD�I8G9GAGBzGC�TPDS��REL�&U�s �� �EST�x��SFSP�C���C�C�NB��S)*$8�*$3%)4%)5%)6�%)7%)S�PNS�TRz�"D�  ��$$CLr   O����!������ VERSIO�N�(  �XK�!IRTU�AL�/�!;LDU�IMT  ���� ���4MAX�DRI� ��5
�4.1 �%� � d%
�Vacuum O�ff����i0ACU?UM_OFF?��K���1���0%	k5n�?�9	�5� �O�7ջ6�0�4
�����1 ��Ι�O�8 GOmO ��"�33�13A2 �׸oONO�OrO�5��F2B2 ļ���O�O(_�O�4 �K 9O_�_�_�H�F�_ �_�_�_�[�3�5�_7o �_[o
oo�o@o�odo vo�o�o�o!�o�oW g�<N�r� �����S��� ��8���\�n������� �ȏڏO���s�"�4� n���j�ߟ�����ğ 9����4���0���T� f�ۯ������үG� ��k��,���P���׿ ����ϼ�1���?� y�dϝ�L�^��ς��� �ϸ���?���c��$� ��H߽�l�~߸��� )�����_��o��D� V���z�����%��� "�[�
����@���d� v�������!����W {*<v�r� ���A�< �8�\n��� /��O/�s/"/4/ �/X/�/�/�/�/?�/ 9?�/�/G?�?l?�?T? f?�?�?�?�?�?�?GO �?kOO,O�OPO�OtO �O�O_�O1_�O�Og_ _w_�_L_^_�_�_�_ �_�_-o�_*ocoo$o �oHo�olo~o�o�o )�o�o_�2D ~�z���%�� I��
�D���@���d� v�돚���!�Џ�W� �{�*�<���`���� �����̟A���O� ��t���\�n�㯒�� ��ȯ�O���s�"�4� ��X�Ϳ|���ȿ�Ŀ 9����o��ϥ�T� f��ϊ��Ϯ���5��� 2�k��,ߡ�P���t� �������1�����g� ��:�L������� ���-���Q� ��L� ��H���l�~����� )����_�2D �h����%� I�
W�|�d v��/��
/W/ /{/*/</�/`/�/�/ �/�/?�/A?�/?w? &?�?�?\?n?�?�?O �?�?=O�?:OsO"O4O �OXO�O|O�O�O_ _ 9_�O�Oo__�_B_T_ �_�_�_�_�_�_5o�_ YoooTo�oPo�oto �o�o�o1�o�og �:L�p�� ��-��Q� ��_� ������l�~�󏢏� Ə؏�_����2�D� ��h�ݟ����؟%�ԟ I���
��.�����d� v�믚����ЯE��� B�{�*�<���`�տ�� �����A���w� &ϛ�J�\ϖ��ϒ�߀����=���a��"� �%
Send E�vents�S�SENDEVNT���Q�.�� %	���Data�߶�D�ATA���(��%���SysVar<;��SYSVw���}0O�%Get�x�GET+��1���%Request Menu����REQMENU?���2�]ߞ�Y��� }�+�����.�� d�7I�m� ���*�N� ����i{�� /��/\/G/�/// A/�/e/�/�/�/�/"? �/F?�/?|?+?�?�? a?�?�?�?O�?�?BO �??OxO'O9O�O]O�O �O�O___>_�O�O t_#_�_G_Y_�_�_�_ o�_�_:o�_^ooo Yo�oUo�oyo�o �o $6�ol�? Q�u����2� �V��������� q��������ˏݏ� d�O���7�I���m�� ����ݟ*�ٟN���� ��3�����i���𯟯 �ïկJ���G���/� A���e�ڿ�����"� �F����|�+Ϡ�O� aϛ�����߻���B� ��f��'�a߮�]�����ߓ��$MACR_O_MAXX��Կ���Ж��SOPENBL ���2��ݐѐ�_���"�P�DIMSK�2��<�w�SU���T�PDSBEX  )K��U)�2��� ���-�