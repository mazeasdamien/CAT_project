��   g�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����BIN_CF�G_TX 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG���DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST��NSS�* 8�D�FACE_NUM? �$DBG_LE�VEL�OM_N�AM� !� FTޒ @� LOsG_8	,CMO>�$DNLD_F�ILTER�SUBDIRCAPCp��8 . 4� �H{ADDRT�YP�H NGT1H����z +�LSq D $ROBOTIG ��PEER�� MwASK�MRU~;OMGDEV���PINFO. �  $$$�TI ��R�CM+T �A$( /�QSI�Z�!S� TAT�US_%$MAI�LSERV $�PLAN� <$�LIN<$CLyU��<$TO�oP$CC�&FR�&�YJEC|!Z%E�NB � ALA5R:!B�TP,�#�,V8 S��$VkAR�)M�ON�&����&APPL�&P�A� �%��'POR��Y#_�!�"ALE�RT�&i2URL �}Z3ATTA�C��0ERR_T7HROU3US�9H!��8� CH- c%�4M�AX?WS_|1;��1MOD��1AI�  �1o (�1�PWD  � LAط�0�ND�1TR=YFDELA-C�0<G'AERSI��1vQ'ROBICLK_HqM 0Q'� XML+ �3SGFRMU3T̑ !OUU3 G_�-COP1�F33�A�Q'C[2�%�B_AU��� 9 R�!UP=Db&PCOU{!�C�FO 3 
�$V*W�@c%AC�C_HYQSNA�U�MMY1oW2"$D�M*  $gDIS��SM	 l5�o!�"!%Q7�IZP�%� ��VR�0�UP� _D;LVSPAR��QYN,
3 �_��R!_WI�CTZ�_INDE�3^`O�FF� ~URmiD��  (d�  � t Z!`M�ON��cD��bHOUU#E%A�f�a�f<�a�fLOCA� #�$NS0H_HE����@I�/ ; d8`ARPH&�o_IPF�W_* dO�F``QFAsD890�VHO_� 5R�42PSWq?�TEL� P����90WORAXQE� LV�[R2�ICE��p��$cs  �S���q��
��
�p��PS�A�w�# XK	�Iz0AL`��' �
����F����!�p�i���$� 2Q� �P��������� Q�b��!�q����$� _FLTR  ��\� �����B�����$Q�2���7rSH`D 1�Q� P㏙�f� ��ş��韬��П1� ��=��f���N���r� ӯ�������ޯ�Q� �u�8���\������� 󿶿�ڿ;���_�"� XϕτϹ�|��Ϡ�� �����6�[���B� ��f��ߊ��߮���!� ��E��i�,��P�b� ���������/��� (�e�T���L�����z �_LUA1�x!1.��0��p����1��p�255.�0��r��n���2 ����d %7I[3e��� ����[4���T'9[5U���{���[6���D ��//)/s��Qȁ�MA��MA��P������ Q� ��u.< �/?&?�/J?\?n?A?�?�?m�P�?�?�?�? �?O.O@OROOvO�O�Ou.kOl�q��O�L�
ZDT StatusZO�O5_G_�Y_n�}iRCo�nnect: i�rc{T//alert^�_�_�_�_mW #_oo,o>oPobot�e^�P~2g���go �o�o�o�o�o�o	�-?Qcul�$$�c962b37a�-1ac0-eb�2a-f1c7-�8c6eb56401a8  (�_��_���"�p�1!W��(��"S��J�E�� X��C� ��,$ ���W���ˏ��� ֏��%��I�0�m�� f�����ǟ�������h!��u�R����n� DM_�!�����SMTP_CT�RL 	����%����DF���ۯt�@ʯ��'��Lz�N��� 
j��y�q�>u����Ԙ��#�L�USTOM �j������  |���$TCPIPd��j��H�%�"�E�L�����!���H�!T�b<�n�rj3_tpd7�� ��i�!KC�LG�L�i���5�!CRT�ϔ����"u�!CONS���M�[�ib_smon����