��   #��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	��/GR�P: $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2(��� RING��<�$]_d�REL�3� 1  	�P CLo: �� �AX{  �$PS_�TI����TIME ��J� _CMD,��"FB�VS �&�CL_OV�� F�RMZ�$DED�X�$NA� %��CURL�W����TCK5�wFMSV�M_LIF	��`;8G:w$�A9_0M:_��=�93x6W� |�"�PCCOM���FB� M�0�M7AL_�ECIr�PL!�"DTYk�R_�"�5L#�1EN�DD��o1� �5M�P PL|� W �  $�STAL#TRQ_�M��0KN}FSD� �HY�J� |GI�JeI�JI�E#3AnC�uB�A���$�A{SS> ���	Q������@VER�SI� W�  XKQIR�TUAL_QS �1'X }��� 	 �� �_w_�_�_�_�_�_�_ �_.on2PQbYocQ�ro`o  ������%VZo o�o�f�k�o�o)&8�kkqrZ������d���<���=L��%�L�3?�M���@�m��� ����ȏڏ����"�04�F�X�� EU��p��{���T  2� �����*�<�N�`�r���Nbџ����ү �����,�>�P�b� t���������ο�� ��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z��������<������� �2� D�V�h�z���������FP��(������ ,P;M�q�������(��$&4 1b\��Q��&O����M�yOD��F@ Of��.>G�@��Sn@�\�<���:zV<�$A���) ��	/���\n���/l/�/�/�/�/��R�t.[}~q��/	?z� ��! �/9?�/]?H?�?�?u��%ΐ345678901�?�4�-�1�� �?��O
O@OROǕ�0 rO�O�$ZE�?�O2O�O �O�O_dO5_G_�O�O z_h_�_�_�_�_*_�_ N_`_�_�_.odoRo�o �_�_�oo&o�oro (N�ou��o< ������j;� ����n�����ȏ �0��T�f�4���X� F�h���䏵�ǟ�|� �����B�T���{� Ο��Z�,����ү� ^�p�A�����t�򯘿 ����ο$����Z��� :�(�^�Lςϔ�꿻� � Ϛ�l���$��H� �ϰρ����ϴ�2��� �����d�5�G���� z�h�������*��� N�`����.�d�R��� �������&���r� (N��u���< ����j; ���n������0/T|2&�(/. �8�$PL�CL_GRP 1��� {px5?�  r/ �+|?�/x?�/�/�/�/ ?�/?I?4?m?X?�? x?�/�?