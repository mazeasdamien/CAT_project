��   ��A��*SYST�EM*��V9.4�0107 7/�23/2021 A 
  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41p� d =R��&�J_  4 �$(F3IDX���_ICIfM_IX_BG-y�
_NAMc M3ODc_USd��IFY_TI� ��MKR-  $LINc �  "_SIZc  �� �. �h $USE_FLC 3!�8:&iF*SIMA7#�QC#QBn'SCAmN�AX�+IN�*}I��_COUNr�RO( ��!_TM�R_VA�g#h>�ia �'` �����1�+WA-R�$�H�!�#�N3CH�PEX�$O�!PR�'Io�q7iOqfOoA�TH- P ?$ENABL+��0BT���$�$CLASS  ����A��5z��5�0VERS��G  {XKAIRTU� �O@'/ @E+5�������-@B{FA@A�E��%A �O���O�O����QEI2\K!+_=_ O_a_s_�_�_�_�_�_ �_�_oo'o9oKo�O�+ W?"Hg@ ���j@�o�o�i��� � 2\I  4%Xo��}A�A�o;_q@P������@�A ����8��)�n� M�A@�c$"+ �k�K-@���ń�AЄX }A@A-@�N��
��.� @�R�d�v��������� П���F�A偍A�� (�:�L�^�p����������ʯܯ�DxL��W� 2�l �O�a�s��������� Ϳ߿���'��A� Z�l�~ϐϢϴ����� ����� �2�=�V�h� zߌߞ߰��������� 
��.�@�K�d�v�� ������������ *�<�G�Y�r������� ��������&8 JU�n����� ���"4FX c|������ �//0/B/T/_q �/�/�/�/�/�/�/? ?,?>?P?b?ah�4�0 ���?�p