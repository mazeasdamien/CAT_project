��  
��A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1�TU4QQ  �AR�x1R� � /$TIT91� �� � �Td�T0�ThP�TU5�V6�V7�V8�V9�W0�W�WOQ�U�W�gQ�U�W1�W1�W1��W1�W2�R�SBoN_CF�!@$<!J� ; ;2�1�_CMNT�$�FLAGS]�C�HEK"$�b_O�PTJB � ELL�SETUP � `@HO8@9 P�R�1%�c#�aREPR�hu0D+�@���b{uHM9 MN�B;16 UTOB�J U�0 }49DEVIC�STI/@�� �@b3�4pB�d�"VAL��#ISP_UNI�tp_DOcv7�yFR_F�@|%u13���A0s�C_WAx�t,q�zOFF_T@]N�DEL�Lw0pdq�1�Vr?^q��#S?�o`Q"U��t#*�QTB��bMyO� �E � �[M�����RE�V�BIL���!X�I� v�R  �!D�`��$NOc`M�|����ɂ/#ǆ� �ԅ��ނ�@Ded �p E RD_E���h�$FSSB�6�`KBD_SEV�uAG� G�2Q"!_��2b�� V!�k5�p`(��C�00q_ED|� � � t2d�$!S�p-D%$� ��#�B�ʀ_�OK1��0] P_C�� ʑ0t��U �`LACI�!�a�Y�� ��qCOMM� # $D
� ��@���J_�\R BIGALL;OW� (Ku2:-B�@VAR���!�AB mPBL�@� �� ,K�q���`S�p�@M_O]˥���CCFS_U	T��0 "�A�Cp'���+pXG��b�0 =4� IMCM ��#�S�p�9���i �_D�"t�b��M�1� h$�IMPEE_F�s��s��0� t����D_���J��D��F��%�q_����0 T@L��L�DI�s@G�^� �P��$I�'�����CFed X@G�RU@��Mb�NF�LI�\Ì@UIR�E�i42� SWIYTn$`0_N�`S 2�CF�0M� 	�#u�D��!��v`(����`J�tV��[ �E��.p�`�ʗELBOF� �շ �p`0���3����� F�2T��A`�rq1�J1��z _To!@��p��g���G�� �r0WARNM�p#tC�v`�ç` �� COR-UrF�LTR��TRAT�9 T%p� $AC�CVq��� ��r$�ORI�_&�RT���S<���HG�0I����TW��A�I�'�T��1D���� �202�a1��HSDR�2��2�2J; �S���3��4��5���6��7��8��9�KD׀
 �2 @.� TRQ�$vf��4'�1�<�_U<�G�z�Oec  <� �P�b�t�53>B_�LL�EC��!~�MULTI�4�"u�Q;2�CHILD��;1���@T� "'�S�TY92	r��=��)�2�������ec# |r056$J ђ�a�`���uTO��:�E^	EXTt��p��2��22"y����$`@D	�`&��p������(p�" ��`%�ak�����s�����&'�E�Au��qMw�9 �% ���TR�� ' L@@U#9 ���At�$JOB����P��v}IG��( dp� �����^'#j��~�L�pOR�)� t$�FL�
RN9G%Q@�TBAΰ � v&r�*`1t(��0 �x!�0�+P�p�%���*��͐U��q�!4�;2J�_R��>�EC<J�8&<J D`5CF9���x"�@�?���P_p�7p+ \@RO"pF�0��IT�s�0NOM���>Ҹ4s�2�� @UR<PPgў�P8,|Pn��0�P�9�͗ RA���l�?C�� ��
$TͰtMD3�0T��pU�`�΀e+AHlr>�T1�JE�1\�J���PQ��\Q8��hQCYNT�P���PDBGD̰�0-���PU6$$Po��|�u�AX����T;AI�sBUF,�l��B�1. ����F�`[PI|�-@PvWEMuXM�Y�@�VFvWSIMQSTO�q�$KEE�SPA ��  ?B�B>C�B�A���/�`��MARG8�u2�FACq�>�SLEW*1!0�����
�zs�CW$0'���pJB�Ї�qDECj�eL�s��V%1 Ħ�CH�NR�MPs�$G�_@�gD�_�@s��1g_FP�5�@TC�f FӓC�Й���qC��+�aVK�*��"*�JRx���SEGFR$`I�Oh!�0STN�LIN>�csPVZ�z���@�D2����r 2���hr�r��1��3` +^?���եq�` ��q|`�����t��|aSIZ#�!� ��T�_@%�I��qRS �*s��2y{�Ip{��pTpLF�@�`��C3RC����CCTѲ��Ipڈ�a���b��MI�N��a1순���D
<iC �C/���!uc�0OP4�n j�EVj���UF��_!uF��N�����|a��=h?KNL�A�C2�AVSC	A�@A��r�@�e4�  cSF�$�;�Ir �3�a��
�05��	D-Oo%g ��,,m����ޟ��   �ǀD�6� n���sυ�Uz��R�0HANC���$LG��ɑDQ$ft�NDɖ��AR۰�N��aqg��ѫ�X�M�E��^�Y�[PS�RAg�X�AZ�П���rEOB�FCT��A��`��2t!Sh`0ADI��O��y�s"y�n!�� �����~#C�G3t!N��BMPmt@�Y�3�afAES$������W_;�BAS#X�YZWPR��*�tm!��	VQR_L
 .� 7 ���C�/�Y(zJ�LB�$��3����5�FOR�C��_AV;�M�OM*�)�SԫBP��H�1�HB�ɀE�F|���PYLOAD&$ER��t&3�2��Xrp�!J"zR_F}D�� 8 T`�I�Y3��E�&��Clt��MS�PU
a$(kpD��7��rb�9�B�	EVIѣ
�!e�X�$I��B@X��X<&v�SY5� / �R_HOPe�: >�pALARML�2W̭r#�R_�0; !hb P�q�`M\qJ@O$PL`A��M����0�E��	���V�T�0�]�U�PM3�uU��<�TITu��
%�![q�BZ�_;��3= �B �pQk��6NO_HEADE^az��}ѯ� �`􂳃���dF�ق�t�pn��>�Ю@��uCIRTR�`��ڈ�L��D�CB@4�RJƱ�u�[Q�н�?��2>���OR�r��OxK��T`UN_OO�Ҁ$����T��Њ��I�VaCnp�D�BPXWOY���@�$SKADR�wDBT�TRL��Az�րfpbDs���&6�DJj4 _�DQ�5�APL�qFwbWA��^WcD�A�k�A=�2CUMgMY9��10�&��DB����B�[Q;PR�� 
� ������C �Y1M$�a$8�b`L��D���7����0E�����PC�1F�/�� �PENEJA@Tf�G=/�����RECOR"H�H @��C$L�#D$�PR���+0jp��nq�_D$�qPROSS�
���
��r� -�$TRIG<� �&PAUS�#lt�ETURN�"�M�R��U� Ł� E�W����SIGNA9LA�QR$LA�0O5��1E$PD�F$Pİ�AGc0�A�1C~4�3��DO��D��"�!&GO_A7WAY�"MOZq��Z�u CSG�CS;CBg�I Իa#��<�ERIL0Nn�T�`$������3�2L\�@	BGAG~@R�P����44BD�/ACD�O�F�qF� YF'C�CM�A� X'C�$FRCINI_�5#Ӑ@���$NE�@�F��4L��� J� ���<����R/���}P\ OVR10����$Ҡ�$ESC�_�`uDSBIO�X��(Te���VIB�� `szLZ��LV���pSSW������V	L�:�Lk�ZX����`��QP���USC�PⓂA���A��MP1��U�C�P��Rt`�S5QeU����Sg�Cg �Sd���dcC��g<.���AUTO$�a҃oac�SB����T����C/B��2�f_$VOLT�g��A� ���1D����a���@��ORQ�Ҁr�$DH_THE� PRp� <)t&wALPH&t��o�Jw�  p���.�R��{s�5c`r��A���ED�S\ F�!M��q�sV�r�v�ûvL��R�tk����BTHR����T`�����zVɖ���Q�D)E7 ��1K�2P�C� X�C�f�F��#�g�� QT,0Т�p���f�d@����g����N~��s2>�Y0INHB��ILT� ɡ�T?� �3��/�఩3�P)Q0QАT)PeŖ0Y�AF5�OM�r�o��z��� o�)Pڳ|���o�P��͘o�PL?�x��o�TMOUXc|��o� � w�+��1�H���A��g�Io�����DqI~���'�STI������O��� Hҽ�ANǥ�Q�S8��b͑�h$kЪ���/�1_Ig�yPRAOP�P�.C��kӦMCN�Qe�E�L�VER�Se��bP'PI/�F�{������G�DEN��G����o�F�2H��ӷo�MԺ�F��_ԴM�D��䧭�@ed��3�ea���DO� ���U��2�j�ʹDI ��e�۴��번�������/�F0�����O�N���ȅQI�VAL�ȤCR�_SIZpJ���A&�REQ�R����2���D�CH )���ʹ��z�D��ō��&�S_�>X��/W�FLG����/U$CV�iM�@VQ��FLX��"�B��-�L����ALJP�C��� �bT^�W^� gR�xc� cQ�NDMS��m�K�C{P_M�  �STW.�������h�AL�PY�YQk�����V��e�IAG@�'�d7���T�	A�P� R��A^�� ]� `]�	`]�6[�q_D��g��c����YP�����r�"8Tc� ?�����1��T��ۡ���LH�?`��! �0��LDĀp��U0JFRI�0 �P��I\15�j�IV1U�s1IU�P�PZ�Q��C�L!W���
�PL�C��S��CWC�	/��  �IZ!Fů�T�Q�g!��?���g��p~�
�P�5RSMI�PT��0  b *�lsd2AWda_T
p�5��0NS_PE�A��;����ܢSAV�����7%I��CAR؀�P�!<$f�E"CR�����T[#qEl@I�\"STD;��[!F�`'�x'QOF07�k%B�"RCO҇&RC��v(���1�R�'�=�G%��WMA�Q_naI��AQ���a$2F�%-4I:�*7I>R99�/Q97��k8M�H!C:�`Rp  tp�2F��SDNX�Va���  �G2�AK P $M!��s�S�1 7��3nc%j9f��4[��RA�D�0CY_ �L L!IG1@0'1BV�1@�07H2��NOà���CDE�VIP M�0�$�RBT�FSP0c3�C-T�DBY4�A��G3�3HNDGD��1N H�0GRP�HE�!XL<Uj�S�DF02��4L�` aO�Bp��U�FBQ\�FEN�@�uSV���3 �1P d�@DyO���PMCS���?P��?PuRN�HOT�SW24�DpELE�1�U�:�3�P�RQ T�@I�[r@  fl�o`OL�GHA8F#��c:����3�A�0�R � $MD�Lb 2Q��E Xȃqn6�q� �i�c�e
�cJ]�	�e���#�nX�d�g]PTOa�� xtb1U�4SLAV�� S  n�INAP���F��By�1_��wENU�1T $
��PC_eq�2 �RL�vw��^tSH=O�� U ��A�a�q�2rr�v�u�v�]sCF\ V�` ,�xr�O�G�W�p�%�q �Ype�rI��!�MAX�,�q0 AY�vWA (�gNTV���rVE�0.�uSKIg�T�`$�}�2S���JsX!���C��s��f��_SyV��`XCLUL�: �p�ONLB�߃�Y�T��OT�UHI�_V�!��APPL�Y��HI�P�v�_�ML�� $VGRFY�����M3�IOC_�Z� 1���l���O�@�LS�/"@$DUMMCY4x𛐒�_C L_TPJ�T�#Cc�1CNF�Օ_E���j@�1���D#Q_0������PCPB��� R S��k���kdo�>�� W ��� �RT_�@`[uN;OC�R X;r���TEL������zDG���x`Y D��P_;BA`#c���!�ȥ_ЀҬH�У6Tb�E�� Z�np�R�SARGI��!$���`Yn�S;GN�1[ ��`��IGNQ�G�J�����VJ�d�[�ANNUN��ޕ��_Ex�'wATCH�������Ķd�r�1\� <�0�@����S	$ah���������ַ1EF I�� �] @�0F��IT>�	$TOT! �C������-�M�@N�Iva^,B��r��A�q��DAY�3LOAD�D�&�~�� �EF��+XI@R_\��I��O���a��ADJS_R_!x``���� 2�"�����ŉ`�_��PI�cѝD��AG����1a 0@��\�=� \������U! ���CTR�LN p b;�T�RA��#IDLE_PW��G�XԮQ���V�GV_WЉ`a ��'��Ax`c�� 1$k��P�STAC�#M��Q����R2 A�e����SW��A����dՉ``f�OH�(�OPP��#IRO�� �"BRK�Ө#AB��o�㾢��   ��F�Չ`b����"@�RQDW��M�S��6X�'2�I�FECALƳ� 10tND��M���B�0�� ���CP¢��N� Y���FLA�#��OV Y�HE|O��"SUPPOd���gL�p��Q��"�Xт��Y��Z��W������P����BтX�Zbq�$Y2@CO@P�S��2
報�b D!���"�RI�0�s�d `�@CACH�5�VcS��+0�LA SUFFI���p7�Yq���r��6'�7QMSW��e 8vKEYI�MAG�TM@S���&�""@rQ�RO�CVIEN�6�f ^aBGL[�F���?� 	aR��gڶ��PST��! �b����������^�EMAI�`N��:E���FAU� 7��h^�Yq�Z�U�3|�q 5�i<' $#�USWи�;ITߓBUF����DN��H�SUB-$�DC���"��p"SAVx%:"#�_q��X��'󀤶P$�UORDO�P_- ^%=�.�(OTT��_�P�ӆ�0LM$��$g��'AX�3.�U�X- ���#�_GD�
�0YN_���7�j�D�E���M����T��F�Q�a��DIBEKDT�0Ch�6�k;r�GN!�&E�$`����QvP��FP 7l (�pSV� �T�ć�[�ka�1��m� <�n���#7C_RYIKQ�#B\� D3pRE��1'DSP6BP�`hIIMx#]C�A��1A��U:G��8!CM�I�P\�C��~ \DTH�^ oSPB��T\�]CH9S�3?CBSCi�m ���V�dVP�#T_�D*cCONVˁG *cT^ ZF- FD�A�ad?C�0"1R�SC�ҜDeCMER�T�1F�BCMP�S�0ETn�S nFU��DU! ���6ђ�CDSI�@� ���O����o�G�QR�Q�U=�MS��Z-�D�P�Tz�Q[�A�1p� "��Q�4$ZO�0+�q�$��U��ޔ�ePM��eC�N�$��l�l�iGR#OU�W����S� �MN�ku�eu�ep
||�i�cH�p!�ez��0CYC��shw��c��:�zDE�_D���RO�aP��qf��gv3�O���vO� �w�tU��B�u��8L�p�ALA �1q�� 1z�Г0�PB�����H0ER�T7��Rr ,�0>��%>�G1MLR1qG0�0Rw�Ց�1s�����Ų���)Pv���C����U��A��2��0V`tH *��L��� 	��V°��12�b�2� ��2���2���2��2�7/�8/�9/�D�1��;�1H�1U�1b�1�o�1|�1��1��1J��2��2;�H�2U�U2b�2o�2|�2��U2��2��3��3;��3H�U�3b�3o�3�|�3��3��3��4L���2XT�ѡ1u� �\0xf\0�Ug0}�@eme�FDR��ovT VE��`�!G�RG�RE��9FG�SOVM6CᵽA�TROV�D�T� 
�MX�INp깅�	���IND(�B*�
Tȑ0E0Z0G-1 ����PM�3�D���RIV�Pq�SGE[AR6AIO*�KڲQN�0��1�(��P�0|�aSZ_MCM8 nG��F��UR�R�w���P!? ̄�]p?&�C�?&�E
�.��:!�PR��x�0��Pq���RI� @:#ETUP2_ y b�F9#TD�@
�7%T�`�>є׎�l�:"BAC�Q2z T�:"�4)��:%�PBW�(�I+FIf�W M�����PTP� �L{UI�{ иqd UR��!��Bp�1P0 �sEMP�p�C2$b�S�?x�n�J��� �#VRT|^��0x$SHOc�9L)��ASSP�!8s��@��BG_;���H���U���b���o�F�ORC���Qd-|�FU�1�2��2�1�� �^ (�} �|d�NAV_a��b����ְS�q��$VISI��ۂSC4SELЮ�� �r5V�pOg�$b�ְ,�b�$r�I���@�FMR2��~ ���P{r ���0����������ƨ���ڲ_ɡ��L�IMIT_���TC�_LMƤ϶�DGgCLF_Å�DY�LD>т�5��yϋ�Rp�M���Sj�-	? T�FS� �T�� Pl�	�3E0�$EX_	 	1P!0YPba	3B5Bs�G'Q��� �d�6�RSWa%ONZPÏEBUG��ߵGiR�`g@U{SBK�a�O1� C�P�O ���P��M�t�Ot`SMu�E��"8�:�F�y`_?E � �0i�^;�TERM%�%No�ORI�1 �&�H0SMpOs� ��&�S`Z(�%��U�P�p �� -E�yb�b�)#� �x�G�*� ELTaO7�p�0BPFI*c��1Ѝa�@$�$�$wUFR��$��0�!0�UH OT7BPqT�a��#3NST�p�PAT�q74PTHJ�a�PE�P�3ap�!ARTi �%� i �12�"REL{:�1S�HFT�B�!?1m8_���R�P�SX& c $r'�0�h����]s\1R�0I�0eU�R �p�PAYLO�@nqDYN_#�O��R?14�Ʌ�@ERV:�
AX� �8^�7�p{2ס�eE���RCN�ɅAS?YMFLTRɅ�!#WJ�'^�Z�E^�i1�IX��QU�D�pAm5� YF�5PFP$CFQ�6kOR�pM��i!�����>0� �EaCH�Hs��T�� �%2���POC��!���$OaP���rc��ֱ,��jbRE�PR�#\1X��q?3eH�R=5��U�X�1��e$PWaR���u�=@R_�S0b4d�t�#UD^��WQ�" ���$�H��!L`ADDR
xfH!GA2eaZaSar�R��� Hl�SSC�ף�e壒eU��eb�SE���;��HSCD��� )$N�zP_�p_��2��bPE�D�o�HT�TP_��H�� (��OBJ�pSb��[$^fLE03s>t� � n�Q�Jp�_U�T�arSKP̘�2�KR�gHIT����zP��Par��`^��P�PSS�����JQUERY_�FLA�!_qB_W�EBSOC���HQW���!���`�@�INCPUVd�O  �vq:�7��d8��d8��b��IHMI_{ED] T �7R�H��?$d�FAV�@ �}��IOL]N�ґ 8l�R����0$SL!R$�INPUT_���$�P��P�� SLAz �������|C��|Bx�����`F_AS����$L��5w���1��b�!;ࢃ���@HY|�l�E�SQ� �UOP�� ` 1���^f8�\�8�c����PP�3�P��Αc�ے|Ė8aIP_ME��nm�� X1�IPZ`<V�_NETV�p�d�R|�+���WD�SP��p���BG�V}`g�MgAm�� �l(�3TA"B<pA�TIԕ�E�� ����0PS��BU ID�r����P���a�d���10��v��������N	� 
���IRCA̰!� ט �Sy�CY�`EAT�K�}�P�8��3h�]�RY0�A���A�DAY_w���NTVA7�Ԡ��܂]5��ά�SCA@��CL@��w�,�Ţz�m����^2�'�N_�PC �)�Ţ��n���� C�\�0rw����`��� 2�n!d����m���ғ�0r��LA�B11�� ��UNIr
���C ITY��He�^e��R�����Ҿ?�R_URLF��7$AL��EN�`��e�t �sTh�T_U>]�ABKY_2�2GDIS����#SJ�m���$`ҙE�"�R����O A��2��Jh��FL+]�������Ѭ
�UJ]R��� �SpF3��7��'��Q���J7z��O�B$J8�!7`��
��7����y83� �APHI� �Q�P�DJ7�J8�2i�L_KE~��  �KZ��LM� � <��XR$�-�C�WA?TCH_VA��'@<��,vFIEL�Pc1y}`���� D '11V0@@���CT����%�� LG ���� $=�LG_SIZ[t�2�� 1�,(�1�FD<�I0�G� �>�/� I�;�.�S 7��� ��(���^��� ���A�� _CAM32

F�A�..��T(-��29�S� S(�S^�_IRi�S �k].�RS��N0 } MZIPDU~���aLN��r��� �p2�O���c�rKPL�DAU!�EA�`Z�nT7-GqHoR��4�BOO�a?�� CK���IT�sk^`G�REk��SCR; �sL��DIF�S� �`RGI"$D�̆?��TH��t4�SAs3�W��4�?�JGM'MgNCH�s4�FN{�b&K?'-�=)UFK(��0K(FWDK(HL.�)STPK*VK(��XK(rK(RS�)HPg+<�CT�#�B?��`�9U�a_$�� %���T�R"G/)�0PO V7�*��#5$W�M)�EX;�TUI=%I ��B�G���Ar�3#�3�; ��$Sű�	�ᰟ�0�NO�6AcNA4�{Q²AI4�8Zt�EDCS���c�QC�cQBOWHOcGS�=ӁBnHSzH�IGNG�ŰY�<!�k�ZD�DEV�'LLu���Y�eФ���TU$=���(�A���*�#Al�����P���3��sPOS1IU2�IU3IQ��2R@eЦ# �S{FP,D��� �����a�uq0��V+ST��R8Y$��0~�P �$E�VC�[ep�`�VfL�kS �eЧ L
�Z��� o�0��SxpO��t�`id�����_ � �t�� p޳��c ��MC�� ��SpCLDP��s�TRQLI��u��i�d�FL\��b���c�D���g�LD�e�d�e�ORG{��! r��RESERV;�LtG��LtR��d��� �� 	�e�%�d�e��PIT�`��	0q�t�vRCLMC�tL^�y]��q��MI�#�������$DEBUGMAS]�������%U�T7@��E���MFRQ���� � "�H_RS_RU�aa�^�Al�#5FREQ�8 t$�00�OV�ER��Y�&��V��PnT!EFI̠%Fa�_��٢X�yt� \8
Ќ��$U�P\�g?�pűPSHP
��	��C@�s���r�sU�$�?(���MISC�ծ Yd��QRQ��	I�3TB�̠ ���1���AXsҀ�����E�XCES"���b�Mj�����t�s����c�SC�P � 	HY���_��~���������MK Ա����%�B_�F�LICAdB�QU�IRE�#MOs�O����`�Lc`M�Ų �`z���a��r�`�ND������Q�#���DO�I�NAUT�O�RSM����@N�r��3x塨a�PSTL�w� 4�LOC�V�RI���UEX��A�NG-B-��aODA\��p����Ю�MF�e����Ybb�0ple�� #�SUPhev	�FX��IGG~ � ��pbc�� E�bc	6bd��݂�R4� �PD��PS�4�s3/�Wf�TI��<pEX��vPIN�� t��+MD��IA)��W@����q��H�����D#IA8��Ñ�W��Ĩ/Q�1��D?)`�O��Ӧ��� �C�UG�VОp-�ՑOr�_�=ѹ ��`0�S�����i�{ءP{�� ���Pz�KqE2��H-$B: n֤�ND2�r�����2_TXkdXTR1AWC���r�MԀ4q�`�P.�}X���P��d�SB)`�USW�CS;�Tf���V�PgULS����NS���n�
u�JOIN@�� u�6`"��r=b@��cb���P�r��0��cb��o�TA8�{����� �Er�S�C����J��
�R�P�L	� ���L�O9>л�m��	�l���Bҍ�����RR2g�� �1}�A�q d%$G�I���GEA��y2���p EP�RINE��<$R���SW0�t�sA;BCŸD_J��z�\-���_J3D
>G1SP���-�P>Be3dG�8`-���J�s�mr�qO�AI<��M�CSKP�j�H3�3��J@L�Q������_AZ�r�6EL�A��qOCMP��M����cRTD�a�1����m��P1���0�Z��SMG� ���tJ�G�`SCLɐ��S'PH_�@L���z-���RTER �����A_D@�!�ڰA�@�SL�$DI�L�23U�DF�_�5!LW;(VE�L�aINwb�0^ _BLW@-�f$��qV$�k'�'|%�s� ECyHR�tTSA_�_����E5`���@B��%�B���!5`_S� ��%�"%��$b��9,&V�DHɐt��=��8P$V�����1$�����6��$�A���g���H �$BE�L.�m��_ACC�El!�7�q�0IR�C_ ��?pNT<��S$PSɐ�bL_���5�c���63�F@�6�ѩ9G�3G3�2S�̑_FQs2P@VA���7��1_MG|�D1DsA"��FW�`Q�`�3�E�3�2�HDE�K�PPABN�7�SPEEfBJQ�O�`��JQ���1�!$US�E_G��PP#�CTERTY�@�0�q �YNf�A=V� ��B=QM9�M�o�m@OX AjTINC'Ԓ��B��D���W��ENC�F��-��1�2���0INPO	�I�2�U����NTV#}%NT2c3_9"��cLOJ ��`��Iנ�!f? @�#��g`�U"�C� �VMOSIxA;�Z��VA��L�PERCH#  >c��� �g�� �ck�$b�tk�\T'UH-@U@�A�2�eLT �6���U�$jv:fgTRK�сAY�� �c�Oq�2^uSs��g8��R�MOM)ҍ���MP���C��0jsACR��DU��KB�S_BCKLSH_C�2�u9�_f��ES�,� ��R
�TQ�CLALM�Tl�p%0<��CHK� ����GLRTYo����T���8Q��Td_UM����C���A����@LMTa _Lq0O����ˇEō�؋Ā�5ᅀ�8v �qYQ�`'��hP	C�a�hH���wE���CMC�Ձ@�GCN�_��N�ӆ��SF�1�iV'R���W�[���bʕ_�CAT��SH���D�V��q�V`~�KA~����PA��&�R_P��ys_� ��Vv���fsx�i�JG�ŰT�v��y�z�TORQUPgRcoy�@OUW�jb{�@ݢ_W�uOt�t1��e3���k3��I�I�Ik3F��P��}@�VC�00
Q�tp�1�w�u@��v䀳JRK�w�����pDB�Mls�pMC? DLe1�bGRV���e3��k3ܱH_��ڳ"@)��COS6�i6�LN ��Y�z�`�e0[ɮ[� -��ʅ�K�׵ZT�jfܱMYb���B���J˾��THET0*eN�K23k3 �_3c�C�B%�CB_3C��AS{ I�-�X�e3X�%��SBe3v�0�GTS��ACzR��A��<�ڔ�$DUf�w�����m%��|%Q�a_ ;��Q��0�3�Kv�s(R��A�A�J�(�3�3�LPH6���U�Sz���Œ��⠣Ƽ����R�Vc�V�X�U0{�V��V��V���V��V��V��V��Hc�|��z��������H��H��H��H���H��OT�Oc�OT	y�O��O��O��UO��O��O��O�ƁF�Eѡ	�ŦV�S�PBALANCE�_���LE��H_�SP�!v�����>��PFULC�$�$���*1�uU�TO_a�i�T1T2e�22NH��2�P ���q&��2�3�q�TpO. �1�IN�SEG�2CaREV8�C`�QDIF9u9�1��,"1�,pO!B�,�öw2Ǡ�P�S��LCHWARL�B�2ABH��u�#�C`��\Q�%��X\qP�
�{&:�F2Z� 
p|"ڡ�1�UROB���CR�b�%p�)  ��C�1_d�T �� x $WEgIGHYP�P$T�d�#{�IYQ`IFQN�@LAGJR)�SJR��JRBIL05OD��pF`2ST�02P�,�0 �0��!� ��� 
�P�2KQ�1 � 2�Qd6DEB�U3L@_2��M'MY9�5�N2��4λP$DA�a$��0v�� 	��DO_�0A�!� <� y6o%�KQ7�IBI2A0N�SH_(`�KPf2O9� �/� %��T�P�Q⭁T��4�0TICYK 34 T1�0%qC��pz@N��TC��R��pKQD"�ED"�E�0P�ROMPYSE6� $IR��IQo�8�B�`RMAIᰄQ4[R�E_*0�C�teq]PR�COD~3sFUQP6ID_��.U��B� G_SU;FF-� $3@Q�A�BDO�G��EC0�FGR*3D"lT�C xTD"�UD"�U��lT�4�0�� H _FIv}19�SORDI13 � �236��R|IQ�0$ZDT5U� �f1�5�4{ *�L_NA%A�z@<b�EDEF_I Lh<b�FXd�EP2�FZ4`�F�c�E�e�FIS�@��Ap�D�c�CVdDё�44��!�Z2DX(�rt~3D��O� BLOCKE2�fS�O`�O�G�alRfPUMkU <blT�clT�elT�bxR nswUgcxT�dxRX6�v �a�SO e��U<b�U�c �S�w�hX?@P �dO@�a��0WMxL�Cs���TE7���4�( $1LOOMB_f���02wVIS��ITY2�Av�OJ3A_FR1IU�� SI�a��B	Rw@҇�@҇3�3
2W��W��찰���9_��QEAS3�R@�����p�Bӆ4Љ�5Љ63ORMU�LA_I2�E�T�HR2��G,g��� Ч<8�5COEFF_O^A�Ԕ^A���G
�3S0�2C�A&�?�3$H�3��)bGR� � � $Cp�BXN@TM6wN�CudBXKsh�CER�T,t�+d�0�  NLLt�TpS6�_SVt����p��0������0�� @�SETU�cMEA�@KPi�0�f1�R� � �  ��  �0��'�$�'�q2�Abz@q7q	t����Rb��A�p�apn��� NPREC�Q,�d1�SK_� 4�� �P�!1_USER��"��3 �����VELe���3 �ܵD!�I`��MT?AC�FG���  �|@�Oj"NORE�� $@'��SI�!��w6M"UX�P��A�DE�� $�KEY_�3��$JOGu��SV�����Ñ!Y�5�SW�j"�aaӍ�T4�G�IY:�4 �� �4  �e'2k!X�YZ�S���3k ����_ERR��� � ��=AP�Є1|��{�$BUFf�qXX�� �MOR4�7� H� CU�$A�k!j��Aa����Q'$� ��aW��$P���G6�� � $SI���Y�İVOY���O�BJEZ�ADJyU�2\�ELAY`�4�%��D
�OU�P�Ÿj�JQ�R=i�T�9��8��2DIR�=�E����� DY�N��"��TY�"R�O@I0�"�OPWwORK���,�0�SYSBU1�Y�SCOP��?Җ���U��b�PCp���PAð�,���f"Y�OP�PU�!��!M�$�IMAG/�� 1�Z23IMz�M�IN��~J�RGOVRDv���İ'�P)�I� ��P�s��k"LApB�|��'�PMC_E`?ѭ1N1 M��1�211�2�v�SL���� � $OV�SL��c��a�`c�2j"��_v�#�Pw��#�P-B=�2bC�� >`��q?w�_Z�ER7���Z�$Gd� 3������G� @����%O6PRI\�� 
�P�	�����PL��� � $FREE��E������Lʶ��e�Tg ^0AT�US��TRC_Ta�N�MBR�W@+���c�1,`��� D�1%�fÌ�L���"��0�QJ ����XEQ3������� � PcUPa��`�aPX�@�w"�43�����PG�ڻ�$S�UB?�%�q?�J?MPWAIT�2�W%LO��FeA�R�CVF�A}@R"Z!R�V�R"ACCt R���pB�'IGNR_{PL�DBTB^0P�aS!BWP�$/��U1@�%IG�@I���TNLN�&�"RȖ�<r�N�@��PE�ED�HADO!W^0��/���EK4�")!W`SPD0!� L<A2�X`k0��y3UNI*�{w0�R�|LY`� I}S�PH_PK�����RETRIE��3�)���0�@FI���� ��P�0�4 �2��DBGL�V�#LOGSIZ,]��aKTw!U��0D�D�#� _T���MB��C��R�V@?MRPC|5���CHECK� NX�	�P�0!�#���9a�L#Y�NPEA*pT�2���@�P1 � h $AR#B!R��S�a���O�P��ATT ���"��#FV@2��aSƝ3UX��B�PL9I�"0!� $���OITCHR"�W���AS�-�QSLL�B0!�� $�BA��DsY�BA�M� f�Y��PJ�5u�	��R6�VzQ_�KNOW�C�Rv�UFd�AD�X�v0Dð~iPAYLOA,���p#c_O�,g��,gZb)cL�q��L_�� !�eb�Q��Trd���fF�iC��P`j+�cd��I`hR��H`g;�|dB>���JQ¦�a_Jja۱��AND:�|�tjb~a���*�PL� AL_ �^Pv0���Q���Ce�D(cEd��J�3p1v� T�@P�DCK��>����_�ALPHAs�sBE0��z�AS|���!>�� � ��"oWD_1)j2SdD�AR���u� ���TIA4/�5/�6e�MOM|�;�[�H�h[�U��Bn AD;�p�H��U�PUB��R`���H���U�S��1p��1 �ف2a�� �BRQ���?� e$PI��1��s̱.g$�kHi$�I
0�I>�IL��}�!}�!��}rr�b��/3HIGmS/3o% h4Ɩh4o%� V�Ɩ���՘�!䙥!o%SAMP�o�8�Ɨ9�o%�Ps ��h���  ��w� ��h0�p�� �������8���-pU�H 0��INǬ-p�Ψ �Ťo"Ъ���0�/GAMM��SS�F� ET��K���D�tv��
$4pIBR��2I�$HI��_�f�O�����E�в�A��ϰ��LW���伀Ϲ����r��0jqC��%CHK���  v~I_����� ,r�x,q��z�s����|y�1s �$cx� 1��I� R�CH_D�!� R1N3��#��LEUࡒ����x���0MS�WFL�$ہSCR�(100;�,@v�3 7B[֝��`;���o�h0�~�PI3A�ME�THOB���%��AX �X20��2�ERI��8�3d�R$�0�e	��pFU�9��}�⌣�&�L8��9�;�OOP}���8Qጡ��APP�3�F��@U�v�a岣R	T��0�Oph0.ŧ�0��턱 1�#�터k ��L���RA�@M�G$�VSV��;P�CURA���GRO50��S_SaA�Q��3��NO�pC���t3����4o FoR�����x��R���� �DOg1A��bAw� qڪ����Aϗ�A��1�-��ic'QPM��o � �YL"��a����S�b4�7B�I���a�Ï�a�_��CѣM_W�b��A���=�M@� ��`�0q|$JԐR1I�"�PM$���C �A{ ��WC�$��L1QVaC �tA�tA�tAUt� �ͰN�P��dS��-pX�0O�s,qZ��Py ��� ���M�� x�u���������2�������5L�q_XR� |tq�3�[��&H��& U�3�4��'�&N�sQ}�PKQ��q"
��KPW`�q$P�A�PMON�_QU=� � =8�@QCOU���@7QTH]�HO|807HYSPES�R80�UE#0)�b OVT�  �0P!��T�R_UN_TO�OP9O���� P`�5�C�|A�INDE>��ROGRA� HP�� 2A�NE_NO��4�5IT��0e0IwNFO�1� `Qh�:�1��l!OI�2�� (��SLEQ��� A�� @�6d1S_�EDIT�1� ��P�Kށ����E澰NUpGjHAUT<O�mECOPYށ��(�L��[�M��N�@�K^K�PRUT� �B�NF�0UlR$G��2�D=RGADJn�1� htpX_� AI���#V�#VW!X�P!X�#VϓP��N^p_CYCoS7NS_h3�q 	��LGOXã�NYQ__FREQÂW֠�:ƴQSIZB��L�^`r�P!QV�֠��CcRE����Y�IF>���3NAA�%�T_}G��STATUt <��w7MAIL?��qx=a�34LAST=a��q�TELEM�Q�; �qNABot�EASI|a1l��  X�kb��<�f�ҳ���I�0�īR��;1� �&�bABS1SpE�0Ӑ9V_a�fBAS]r�eď�āU񐳐H�Y$qwRM�R�c ����:s�𐠲Xatg L�T��| �	�b 2�  ���䤏v(r�w]r ����(r�w� �DO�U�3��p��$$C�X`S0�� ��5�c�c� �pY�sSI9����XK�IRTU�����A� _WR�K 2 @�� 0  G�5�w���t�.�� ��	ɀ��ݏc�A��ˏ�����,�8�ȁ>�s���̍�Q�BSSA� 1�"�� <a�ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ���߰������ߝ�CC��@XLMT0������  d��IN�����P�`EXE�'�S�6�^0-r ���@�Q�DV��Svp�@�S�%sel�ect_macr�o�߫���IOgCNV�c	� ��P��Up(㲗��0�V 1^�P $�N���H�B�E�A�?���k h�z������� ��������
.@ Rdv����� ��*<N` r������� //&/8/J/\/n/�/ �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�? �?�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� � 2�D�V�h�z������� ԏ���
��.�@� R�d�v���������П �����*�<�N����LARMRECOV ���6�!�LMDG 1��<�����_IF� 1��d  �YST-040 �Operatio�n mode A�UTO S��ed� P) d ou�t ��for BWD��7�?��S�e��w�������, 
� ��ҿM�>IP�L_FANUC_�SMPLG>  LINE 0 ���ABORTED���JOINT 100 %׿:�!��$�RP_CL�O�@��k�E�S�BN-060 I�nvalid a�ttribute� syntax data����������NGTOL  �j� 	 A �  1�C���PPI�NFO ��� ��v߈ߚ߬��  �����ߕ���� ��)��%�_�I��m����O�������� 	��-�?�Q�c�u����������PPLI�CATION ?}������LR Ha�ndlingTo�ol� 
V9.40P/17B�>��
883�� 
F0F3170�2 
'7D�F5 ���Non}e��FRA��� 6c��_A�CTIVi�]�  ���*�  ��M�ODi���(��CHGAPONL{ +OUPL��;1	ة� hl�~��CUREQw 1
ث  T���	���� $�����//'/�9/�/]/��Κ� �$H��k�*HTTHSKY�/���$\~/ �/>??r/,?J?P?b? t?�?�?�?�?�?�?:O OO(OFOLO^OpO�O �O�O�O�O�O6_ __ $_B_H_Z_l_~_�_�_ �_�_�_2o�_o o>o DoVohozo�o�o�o�o �o.�o
:@R dv�����*� ���6�<�N�`�r� ��������̏&���� �2�8�J�\�n����� ����ȟ"�����.� 4�F�X�j�|������� į�����*�0�B� T�f�x����������L俬TO����DO_CLEAN�8�o�NM   � ����������ߠDSPDR3YRv��HI��@��q߃ߕߧ߹��� ������%�7�I��MAX��V���G�g�XV�fcf�PLUGGVW�cWPRC(�B����`�R���O��1�C�/SEGF/K�� *�ϩ�q�����������$�LAPN�a��# 1CUgy�������*TO�TAL���KUSWENUN�[ <��@鲬RGDIS�PMMC-�!1CL5�y�@@C�[OL��n�9�W_STR�ING 1'
_�M S�
�
�_ITEM1�  n��� //*/</N/`/r/�/ �/�/�/�/�/�/??�&?8?I/O �SIGNAL��
�ײ����������޼��ƭ�خ���ޮ����5���9��������� = 10�0������������۸���� ��1�2�t3�5�3ʰ���ް� t�M?H �װ��A����??=??OQO cOuO�O�O�O�O�O�R��R���O,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^opo�OWOR-���a _�o�o�o�o* <N`r����������&�P	O�e	L��k5�o� ��������ɏۏ��� �#�5�G�Y�k�}���p����şG�DEVO� �c�ݟ�)�;�M�_� q���������˯ݯ﯀��%�7�I�[�m�PALT]���on� ��ο����(�:� L�^�pςϔϦϸ���p���� ߂�GRIl� �8Ѭ��`�r߄ߖ� �ߺ���������&� 8�J�\�n����&�R]��P߶��� (�:�L�^�p������� �������� $6<H��PREG���  ��Z����� &8J\n��������N=�$�ARG_�`D ?�	���/!��  	�$N6	[C(]�C'�N7d)" SBN_CONFIG�0�/+�1�2�!|!C�II_SAVE � N4�!�#" TC�ELLSETUP� /*%  O�ME_ION=N<%?MOV_H� �/�?REP��M?*U�TOBACK� �/)�!FRwA:\n X?,n� '`�0n�8�� �;�  �20/07/�31 12:49:12ne(nO0 OMODO�<��mO�O@�O�O�O�O�On��O _._@_R_d_v__�_ �_�_�_�_�_o�_*o <oNo`oro�oo�o�o��o�o�o��� � �1_p3_\AT�BCKCTL.TM;�Sew��b;INI���5�&j3?MESSAG� �q�!7 �#�!�qODE�_D� �&�%�xOx��j3PAUS`�� !�/+ , 	�e /%d�r�,		\������� ������ڏ��� �J��4�n�X�z���7�A�TSK  G��?��m0UPDT�p�wd���XWZD_�ENB�t�*�ST�A�u/!�!!XIS>� UNT 2ǖ�!�� � 	 ���l�J�7C� ��� ]�� �n
�|������!"��
����,��Я�|��G�P �b �u�+ %M> ?A8R ��N'ȯ�)��M�+^�METV��2j��� P{��B95@�-�A�B4@���A/�yB"�v�7�>�8=�&��=�Q�<�I_=?�*��7_��SCRDCFG �1/%�1 	��%�"E��+�=� O�a�sϚ?n
Q�)� ���������߄�A� ��e�w߉ߛ߭߿�&�`�'p1GRc��%����6pNA0.+	�p4��_ED�p1��� 
 �%{-<pEDT-�߰*:|����Y�#���f�q2o�n
e"�cO6h������2 �);��l�*��q1:�@�������"�
�3�� M�*q���q����`��
�4��= ���=��,�
�5u��	���	/ Pb��
�6A/� �/���j/�//./�/R/
�7?}/Z?�/���6?�?�/�/�??
�8�?��&O��]��OmO �?�?\O�?
�9�OO�O9O`���O9_�O�O(_�O
�CR�H?�_ �_~=�_oJ_\_�_�_���K�NO_DEL�
��GE_UNU�SE��IGAL�LOW 1.��   (*S�YSTEM*4��	$SERV_GqRE{�`A�REG�e�$�c4��`NUMx�js�mPMUi`>4�LAYu�4��PMPAL|�p?uCYC10Jn�]~GpK~�sULS�U=�m_rA��cL���tBOXORI��eCUR_�p�m�PMCNV9v�p10s~%�T4D�LI%���i	*P�ROGRA�dPG_MIK~u����ALU���~���B����n$FLUI_RESUcw��o��!�MR�n�`l o,�e�w��������� џ�����+�=�O� a�s���������ͯ߯ ���'�9�K�]�o����\bLAL_OU�T �k���W?D_ABORdp�n����ITR_RT/N  T��i�?NONSTOB��� ��CCFS_UTIL .����CC_AUXA�XIS 3N� h���Ϧϸ������CE_RIA_IL�`�Кa@�FCFG N��Y�M�
�_LIMv�b2U� �P7� 	��B\��T�P
���Y�Z�U�Y����� �Թ��Yq��Q��$��v�X
_��"��9�PÀGP 1r�#��k�}﨏��`�C�`C�@CU7��J��]��p��}����� C���U���������U������������U���������;���pCk������������������������������� D� DK��K�K�K� ��V?�3�HE8`O�NFI-��m�G_�P�1r�  Uerŷ����������#5m�KPAUSf�q1r�� sr 7}r�k���� ��9Io�U����?�A�ii�4�M�NFO� 1H�$�� �]�9/T^��h�>F�d9��]�/�A/�� D&�t����D�)�´ ²?E�³��z/�'@�O� �*ز!�LLECT_�!0H���3��$ENU�Ÿ�b�Ҳ!NDE�#�#H�Y�12�34567890�I7R�a$�G?Y6��H��S)�?�?�\�?�? �?�[�?�?BOOO1O �OUOgOyO�O�O�O�O _�O�O	_b_-_?_Q_ �_u_�_�_�_�_�_�_�:oo#6B�$�+ ��-'2IO &29��k#Ƽo�o�ol�o�gTR?�2'nm�(�؈2o ~x�(�m*z-��&_MORS�3)r͌a��u]� �y�������rT:�q*r�,}�?f�f�f���Kp���4�%P,2,�/.�e／ Ώ�������8u�k)@o,�k#� � ja�(P�DB.0.ʼ)dc?pmidbg]���L��ʓ:�n��p��|��Ȗ  �n��A��X�!��l����f�mgz�ӯ�� �f¯�� �>-`ud1:@�i��+ꂑDEF -���c)T�cy�b?uf.txtt��u���=�/nm��>�����a�MC&�r20��|cdC�$��s212ͤ!�q�k&�CzkЎ1^�A���hAӡ�A��߈B5O����C�4 y�H+C3/��C%;]C���D}�C����D�F-Ev��@F?�UE�f�E�v�E�/F��n�?���l�<�23nlD�)�h1��!��2�ӧ�5���
&pxc��}���  D4q���λG��  E%�q�F�� E��p͟�F-F�P �E��fF3�H ��GMx����_�>�33���i�G�nc�G�@�#5����G�Ai�k$=L��<#�{u��`V��c:��R�SMOFST �+����P_T1:�4nmA g���MODE 5��Ʊ`��3q�w!;��-�O�I�?����<�MܾTES�T��2����R�"60�/y�uƦ� Al�k(��� b���C6�0B���CE���s���:d�{s +���*!�����^�T_��PRO/G %G�%ӿL|[��`NUSER��`KEY_TBL�  G�!$"�	�
�� !�"#$%&'()�*+,-./R7:�;<=>?@AB�C��GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������&���͓���������������������������������耇���������������������  LCKjp�aj OSTAT�\�X1�_AL-�p1}_AUTO_DO6�o�#FDR 3]8��2hk)U;`/r/�/�$O/�/H� -�k��/5����)�/�/ �/<?>O?5�\�J�N/ �?�?�?�/�?!Oe�T� ��8ObOh3fOPO�O�O nO�O�O�O
]�?/_A_ S_�?d_�_4O�_�_�O �_�_�_�_�_o(o^o po_�o�o�of_�o�o �_*o,Xf <z����o�� #��o4�Y�z�t�� ������Ώ�����.� @��g�y���6����� l��ܟ�����(�6� �J�`�����V�ϯ� 󯞟�)�ԟJ�D�b� d�V�����t���ȿ�� Ͼ�7�I�[��lϑ� <��Ϭ�ʿ�Ͼ���� ���0�f�x�&ϟ߱� ��n����ߤ���2� 4�&�`�n�D����� �����+���<�a� ��|���������� ���� 6H��o� �>���t��� �0>Rh� �^����/1/ �R/L/jl/^/�/�/ |/�/�/??�??Q? c?/t?�?D/�?�?�/ �?�? OO�?"O8OnO �O.?�O�O�Ov?�O_ �?"__:O<_._h_v_ L_�_�_�_�_�Oo!o 3o�ODoio_�o�o�_ �o�o�o�o�o�o> P�_w��Fo�� |o��
��8�F� �Z�p�����fߏ� ���9��Z�T�r� t�f�������؟�  �ΏG�Y�k��|��� L�¯��ڟܯί�� �*�@�v���6����� ӿ~��	ϴ�*�$�B� D�6�p�~�TϒϨ��� �Ϟ��)�;��L�q� ϒߌߪϬߞ����� �����F�X���� ��Nߴ��������� ��@�N�$�b�x��� ��n�������A ��b\z�|n�� ���(��Oa s��T��� ��//�2/H/~/ �/>�/�/�/��/? �2?,?J/L?>?x?�? \?�?�?�?�?�/O1O CO�/TOyO$?�O�O�? �O�O�O�O�O__N_ `_O�_�_�_VO�_�_ �Oo�__ooHoVo ,ojo�o�o�ov_�o �_$I�_jd�o �v������ 0��oW�i�{�&���� \ҏ̏��ޏ�&� ��:�P�����F���џ 㟎����ď:�4�R� T�F�����d������  ���'�9�K���\��� ,�������������� ̿
� �V�h���ϡ� ��^����ϔ�
��"� $��P�^�4�r߈߾� ��~���	����,�Q� ��r�l�ߌ�~���� ������&�8���_�q� ��.����d������� ���� .BX� �N�������! ��B<Z\N�� l���/�//A/ S/�d/�/4�/�/� �/�/�/�/�/?(?^? p?/�?�?�?f/�?�? �/OO*?,OOXOfO <OzO�O�O�O�?�O_ #_�?4_Y_Oz_t_�O �_�_�_�_�_�_�_.o @o�Ogoyo�o6_�o�o l_�o�o�_�o�o(6 J`��Vo�� ��o�)��oJ�D�b d�V�����t���ȏ�� ��7�I�[��l��� <�����ʏ̟����� ܟ�0�f�x�&����� ïn�ԯ������2� 4�&�`�n�D�����ο ࿎���+�֯<�a� ���|Ϛ��ώ����� ���� �6�H���o߁� ��>Ϥ���t������ ���0�>��R�h�� ��^���������1� ��R�L�j�l�^����� |�������?Q c�t�D����� �� �"8n �.���v�/ �"//:</./h/v/ L/�/�/�/�/�?!? 3?�D?i?/�?�?�/ �?�?�?�?�?�?O>O PO�/wO�O�OF?�O�O |?�O�O
O_�O8_F_ _Z_p_�_�_fO�_�_ o�Oo9o�OZoTor_ tofo�o�o�o�o�o  �_GYko|� Lo���o������*�@�v�\��$C�R_FDR_CF�G 9Z���q
UD1�:�w�tJƄ  �Ҁ�|��HIST �3:Z�  �� � ?�rU@�A�B�C�pU�D�E�I�Ug�p�o�w��h���INDT_E�N��t������T1_D�O  �u��z�T�2����VAR 2m;���� h'� A&����&�r��'L�'�L΍C��rZ��ST�OP����TRL_�DELET6�Ɣ �n�_SCREE�N Z����kcscy�U_�MMENU 1<���  <�|% ����tۯ�:��s� =�v�M�_�������� ��˿�*���`�7� Iϖ�m�ϥ��ϵ��� �����J�!�3�Yߒ� i�{��ߟ߱������� �F��/�|�S�e�� �����������0�� �f�=�O�u������� ��������)b 9K�o���� ���L#5� Yk���� /�y~��_MANUA3��e���ZCD��=x㙵�/%  "��r�Ԇ
*n'
*?|�(��pd<'GRP� 2>��B1� h ���"h ��$DBCO��R�IG�����"G_E�RRLOG ?�ʫ�q�/1?C?U? ��!NUMLIM�ē�!��
�!PXWORK 1@ʫ ?�?�?�?�?�?m��DBTB_y� !A=���!;Bl ���DB_AWAYz�#�qGCP ���=�ׇ2UB_AL(s0..�"_�"Yb���p����S@ 0 1B�+ , 
�?�O
$�O_H_M���_L�@�%UONTIM6������GV�I�
}P�GMOTN�EN.�.&}[REC�ORD 2Hʫ� �_�sG�O� �Q�_
+`B	oo-o?o �XGono�_�oo�o�o �oqo�oo4�oX j|�)�!�E ���0��T��x� �������ҏA���e� ���>�P�b�t�㏘� ���+�������� :���3�͟�������� '�ܯǯկ����� J�\�˯��k�y���%� 7����m�"�ϣ�X� ǿٿ�Ϡ�7ϯ���E� ��i�{�0�B�����x� �Ϝ��������ߑ��QBTOLEREN�C^DBȧBl@L���� CSS_CC�SCB 2I�,DP
$�O
.c��� ��?�������(�:� L��p���
+�`��� ��������!3E Wi{����� ��/ASe w������� //+/=/O/a/s/�/��/ ���/�/����+:�LLE�JI��UQ4<C:A C��C�{0.0�ޮF? A�+�p+��C�P�q1�- 	 gA�k0�0B���9?�  �6��?�?�(DP��qP��B���HC[�3OEOWO��{O�(kO�O[O��OO��K��L��d������?8;V��'�[�O���OH_(#21��@��7_�_�_�_��vPA.��_c8.�A �_o�WqQm1�1m1!m�QB�QBoLb�)e�Yo�o�o�oQZPz��`�`0�D20�Ca� @��
��!X�&R[�� 5_��>7�����Yk }�"w�a$1W2�!�"{$5�ךO��O���8�J�\���MaCH�+�>1�?3B�Dz��D~���%O��ď�Hݏ��K	���2%����"CR�A�P�W1_�/�t��=R� t�r�R���ʟ����Пޟ�9��#�q`H��� ������a����*3Ʃ ������!��E�W� 6�{�Z�l���ÿ�o�b��"��q2��Az&�4���B7YB#��@�m@$?Y*���ʿB�T�f�x����"H�� �������ϑȴ�!�� E�W�i��0ߝߐ��� ��r��߮��-�?�Q� ��u������߆� �����)�;���_�>��P���t��s����x� h���0'9 f]o����� ���,��OY �}������ �(//1/K/U/�/���/�/  z/���/ �/??5?(?Y?L?^? �?�?�?�?�?�?�?�?  O1O8UOt/^O�O�O �O�O�O�O�O�O__ $_Q_H_Z_�_FO�_�_ �_�_�_�_oo o2o Doqohozo�o�o�o�o�Է	  �a���`�����pZ�`�/- R=pva�C� �<�q
S�����h�:�2���#��K�x����i�A   ��<��m�@�  Տ�t͂С���Ѡ�=�賖 ��Ͽx�+Ă�C�  M��3�t��Ӄ>��{�����S��@a@�������B�S��>����C�������͂��<�o?��PH�)S�B�����������B!ܿ�ͅ1�+��9��� m�b�i�20K���5�!��@��	�@$X�Ƕ�9��q��]A���
y�@q._^B]��т��¡`  ?��ͥͿ<�u�{?���e�ܱ��Ծ�$DCSS�_CLLB2 2=K����p��~'�NSTCY �2L���  h�믊��� ����ҿ�����,� B�P�b�tϊϘϪϼ���Ϸs)�DEVIC/E 2Mm���(��>�P�}�t߆� �ߪ߼��������� C�:�g�y��������)�HNDGD 3Nm�pCz�k)�_LS 2Om�G� 9�K�]�o������������PARAM �P8����H��RB�T 2Rm� K8�p<	����Ⱥ�Q�T������Rh��1�@� ��CW  �B\@`6�B	�� �����@R���H�b��������.���	>,�Y�kJk����c ��; M�T����0/�//f/�A�S�=D �C��ׂ!т�1@#��@�I&�@R�\@g�;?��j���B�&fB�D�CC3$�C2�oC3Ф����A����B8�yB�BA����.��mB����C�RC3��C4
C3���a�(�35P<8�@ "E/W/�??/m??�? �?�?O�?�?8OO!O 3OEOWOiO�O�O�O�O �O�O�O�O__j_A_ S_�_�_l��_�_�_�_ o	oBoTo?oxo�[? �_�_q_�o�o�o�o�o 4/ASe� �������� �f�=�O���s����� �_o��,��)�b� M���q����o��ŏ� ��۟�:��#�p�G� Y���}������ůׯ $����Z�1�C�U��� y���ؿ����� ϛ� D�/�h�Sό�wω��� ��������.��� )�;�M�_߬߃ߕ��� ����������`�7� I��m������� �����J�\��π�k� ��������������" ��+�=�jAS�w ������ T+=Oas�� ��/��//'/ 9/�/�/�/�/�/�/ ?�/(??L?^?9g/ y/�?}?�?�?�?�?O �?�?OZO1OCO�OgO yO�O�O�O�O_�O�O D__-_z_Q_c_u_�_ =?�_�_
ooo@o+o doOo�oc?u?�_�o�_ �o�o�oN%7 I[m���� ����!�3���W� i�����������yo"� �F�1�j�|�g������ğ�h�$DCSS�_SLAVE �S������ښ_4D � ��AR_M�ENU T�  ��R�d�v��������b�A�֯�֞'�SH�OW 2U� � ��Ձ/�9�@� ^�p�����������ܿ� � (�"�L�I�[� m�ϑϣ�ʿ������ ��6�3�E�W�i�{� �ߴϱ��������� � �/�A�S�e�w�ߛ� �������
���+� =�O�a���������� ������'9K r�[�������� ��#5\�k }������� //1/XU/g/�� �w/�/�/�/�/	?? B/??Q?x/�/�/2?�? �?�?�?�?O,?)O;O MOt?nO�?�O�O�O�O �O�OO_%_7_^OX_ �O_�_�_�_�_�_ _ �_o!oH_Bol_io{o �o�o�o�o�_�o�o 2o,VoSew�� ��o����@ =�O�a�s�������� ͏ߏ� �*�'�9�K� ]�o�����"���ɟ���CFG V������_FRA:\	�L��%04d.CSVj�	��}֟ ���[A O�CHW�z���g�񏋯����u������į֯�u����JP�����������RC_O�UT W�����+�۟_C_F�SI ?Q� �u����� ��޿ٿ���&�!�3� E�n�i�{ύ϶ϱ��� ��������F�A�S� eߎ߉ߛ߭������� ����+�=�f�a�s� ������������ �>�9�K�]������� ����������# 5^Yk}��� ����61C U~y����� �/	//-/V/Q/c/ u/�/�/�/�/�/�/�/ ?.?)?;?M?v?q?�? �?�?�?�?�?OOO %ONOIO[OmO�O�O�O �O�O�O�O�O&_!_3_ E_n_i_{_�_�_�_�_ �_�_�_ooFoAoSo eo�o�o�o�o�o�o�o �o+=fas �������� �>�9�K�]������� ��Ώɏۏ���#� 5�^�Y�k�}������� ş�����6�1�C� U�~�y�����Ư��ӯ ��	��-�V�Q�c� u������������ �.�)�;�M�v�qσ� �ϾϹ�������� %�N�I�[�mߖߑߣ� ����������&�!�3� E�n�i�{������ ��������F�A�S� e��������������� ��+=fas ������� >9K]��� �����//#/ 5/^/Y/k/}/�/�/�/ �/�/�/�/?6?1?C? U?~?y?�?�?�?�?�? �?O	OO-OVOQOcO uO�O�O�O�O�O�O�C��$DCS_C_�FSO ?����Q P �O�O<_e_ `_r_�_�_�_�_�_�_ �_oo=o8oJo\o�o �o�o�o�o�o�o�o "4]Xj|� �������5� 0�B�T�}�x�����ŏ ��ҏ����,�U� P�b�t���������� ����-�(�:�L�u� p���������ʯܯ�  ��$�M�H�Z�l��� ������ݿؿ���%π �2�D�m�h�z�_C/_RPI^._�� ����Ϩ�_���W�X��{�^SL��@L� ���� �����H�C� U�g��������� ���� ��-�?�h�c� u��������������� @;M_�� ������ %7`[m�� �����/8/3/ E/W/�/{/�/�/�/�/ �/�/???/?X?S? e?w?�?�?��9��߬? �?OO+O=OfOaOsO �O�O�O�O�O�O�O_ _>_9_K_]_�_�_�_ �_�_�_�_�_oo#o 5o^oYoko}o�o�o�o �o�o�o�o61C U~y����� ��	��-�V�Q�c� u������������ �.�)�;�M�v�q���𕟾���&�NOCO�DE X=���'�PRE_?CHK Z=�А�A А�< �Ր=�E�W�=� 	 <9������3 y�ïկ�������� A�S�-�w���c����� ��������+�=�� a�s�i�[ϩϻ�U��� ������'���]�o� Iߓߥ�߱��ߵ��� �#���G�Y�3�e�� �ϗ�����q������ ��C�U�/�y���e��� ��������	��-? KuOa��� �����);_ qK������ �/%/�I/[/5/G/ �/�/}/�/�/�/�/? �/E?W?�/{?�?g? �?�?�?�?�?O�?/O AOOMOwOQOcO�O�O �O�O�O�O_+_!?3? a_s___�_�_�_�_ �_�_o'oo3o]o7o Io�o�oo�o�o�o�o �o�oGY3}� I_w������ 1�C��/�y���e��� �������я�-�?� �c�u�O�������� �󟍟�)��5�_� 9�K�������˯ݯ�� �����I�[�5�� ��k���ǿ��ϟ��� ���E��1�{ύ�g� ���ϝ���������/� A��e�w�Q߃߭߇� ���������+��� a�s�M�������� �����'��K�]�7� ����m���������� ��5G=�/}� )������� 1CgyS�� �����/-// 9/c/Yk�/�/E/�/ �/�/�/?)??M?_? 9?k?�?o?�?�?�?�? OO�?OIO#O5OO �OkO�O�O�/�O�O_ �O3_E__i_{_U_g_ �_�_�_�_�_�_o/o 	ooeowoQo�o�o�o �o�o�O�o+�oO a;m�q��� ����!�K�%�7� ����m���ɏ��Տ�� �o5�G��S�}�W� i���ş�����՟� 1���g�y�S����� ����寿�ѯ�-�� Q�c��K�������Ͽ Ώ�����M�_� 9σϕ�oϹ��ϥϷ� ����7�I�#�m�� u�gߵ���a������� 	�3���i�{�U�� �����������/� 	�S�e�?�q����ߣ� ����}�����O a;��q��� ��9K%W �[m����� ���5/G/!/k/}/W/ �/�/�/�/�/�/�/? 1??U?g?A?S?�?�? �?�?�?�?	OO/O QOcO�?�O�OsO�O�O �O�O__�O;_M_'_ Y_�_]_o_�_�_�_�_ o�_o7o-O?Omoo o�o�o�o�o�o�o�o !3?iCU� �������� 	�S�e�?�����Uo�� я㏽����=�O� )�;�����q���͟�� ��ݟ�9�K�%�o� ��[������������ ��#�5��A�k�E�W� ������׿�ÿ��� ���U�g�Aϋϝ�w� ����ɯۯ	�ߵ�'� Q�+�=߇ߙ�s߽��� ���������;�M�'� q��]������������$DCS_SGN [���-��^�>	�29-NOV-�25 10:31� ��6�0- 7-�E�  12:49� `�`� [�}S�n�P�f4�n�j�`��k�2�ե��U�Þ�;"�0>~�  �HO�W \��� `��VE�RSION �%�V4.5.�2��EFLOGI�C 1]���  	������+	���:PROG_E_NB  ��"�c�[ULSE  �@s_AC�CLIM���ud�WRSTgJNT�-���EMOdb�w� INIT ^
����OPT_S�L ?	���
 	R575��VE74J6K7K50o1o +	�|(TO  4���V� DEX҆d-�`�#PA�TH A%�A�\�S/e/��HCP�_CLNTID y?��" ,����/��IAG_G�RP 2c������b�	 �@�  �"ff�?aG��%��� BG�  ?��1� 0�C?1>@c��j2!��7@�z�@^��@
�!���mp2m15 �89012345�67�0���� � ?��?��=q?��
?���R?�Q�?ѯ�?ʼ0��0�?(�?�z���0�`�@�  AG�A�p�0�10A� 0� 0G�B4�� ��4`�
�1@����@��\@~��R@xQ�@q���@j�H@c��
@\��@U�@Mp����?�?�D��#@��7IH���@C\@>L@9���@4x0/\)@)��@#\@{@�jO|O�O�O�O8G�?���?��0��� G@?}p�?u?n{?[@;?\�0Q��O_�_,_>_PX�
=?���0�tP_U� 0z��H?p�0h��?^�R�_�_�_�_��_PX�5�\P�� �� 0� `�0?�tP� � #`o o2oDoVo8G ����oAS�o' q�y��[m� �+�	�O�a��m��ÀqbRB�@jRcQ�`
=?��ʆ�\Pׄ
=�5!��4V����
=�b��a&���U?� @C��``3�=q�=b���=�E1>�J��>�n�>��H�
=<�o ~��s������ �`�C޷`<(�Ub� �4�"��@ß���A@`�?5������ 8�J��Ȼ�V������ද��گ쯖�>J����bN�
=�'�G�6���@{`^��pP��0k�@f�fZ>!T@��33�푒�(��
=C��� ��I�CH��)C.dB؃�
= B׿ݱɼ' �  �
��a'�B3Ğ�,��N�B��`�X���wωϰ���3~���l�_?�(�k�R������!�`�~�lD&t�����D/�`�>�s���o�ߢ˻6�<҂������ ²X����AD
� ��߯ߚ��߾��������n��*Iҥ	��W��!CT_CON�FIG d�'|�d�egA��!STBF_TTS�
s	�����e�:���MAU� h~��MSW_CFv��e�+  @��OCoVIEW��f	�1���/[�m���� ������I����� &8��\n��� �E���"4 F�j|���� S��//0/B/� f/x/�/�/�/�/�/a/ �/??,?>?P?�/t?��?�?�?�?�?^�RC�gΥ��!j?NO ;O*O_ONO�OrO�O���SBL_FAUL�T h�:��AG�PMSK���Gj�TDIAG iz��������UD1: 67890123451R��%Q��EPD�m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�oLV�!V�i�
\_�od�TORECP
_Z
*T CW5{[_Xj|� �������� 0�B�T�f�x��o�o�o����UMP_OP�TIO%��NځT�R���I��PM�E���Y_TEM�P  È�3�B+�O��*�9�U�NI���O���YN_BRK j4�~�EDITOR����(���_�`ENT� 1k�9  �,&IP�ANU�C_SMPLGRP_CLOSEȏ�&FS_MOV_5DEG �'OPE%��������EAS_W�RK2FpG��A�NIMA�_DR�Oq�W��30�K��� �-BCKE�DT- _PIC�ɯ��HOME ��*�&PROG_1 �������|J��MAIN q�>��&DE�C����GETDATA4˿ݿ��1 ���&&�1 �B���AAA �R���&�y϶��TE�� 4?���@�1 ����&�O4�1䜐MGDI_STAb�>�O����NC_INFO� 1l	�������@����ߢ�n�V�1m	� �~�����
�
�d��=�O�a� s����������� ��'�9�K�]�o��� ������������� 	*�8J\n� ������� "4FXj|�� 
�����/!+/ =/O/a/s/�/�/�/�/ �/�/�/??'?9?K? ]?o?�?�?�?��?�? �?�?/#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_ �_�?�_�_�_�_Oo -o?oQocouo�o�o�o �o�o�o�o); M_q���_�_� ���o%�7�I�[� m��������Ǐُ� ���!�3�E�W�i�{� ����ß՟���� �/�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���'�9�K� ]�oρϓϥϷ����� �����#�5�G�Y�k� }ߏߩ���������� ���1�C�U�g�y�� �����������	�� -�?�Q�c�u����ߓ� ���������); M_q����� ��%7I[ m�������� /!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�� �?�?�?�?�OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�?�_�_�_�_ �?�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy�_ �����_�	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q�������˟ �����%�7�I�[� m��������ǯٯ� ���!�3�E�W�i��� ������ÿտ���� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a�sߍ��ߩ߻� �������'�9�K� ]�o��������� �����#�5�G�Y�k� �ߏ������������� 1CUgy� ������	 -?Qc}�o�� ������//)/;/ M/_/q/�/�/�/�/�/ �/�/??%?7?I?[? u��?�?�?�?��? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_�??�_�_ �_�_�?�_�_oo+o =oOoaoso�o�o�o�o �o�o�o'9K ]w_�����_� ���#�5�G�Y�k� }�������ŏ׏��� ��1�C�U�o]��� ����������	�� -�?�Q�c�u������� ��ϯ����)�;� M�g�y�������]�ӟ ݿ���%�7�I�[� m�ϑϣϵ������� ���!�3�E�_�q�{� �ߟ߱�˿������� �/�A�S�e�w��� �����������+� =�O�i�s��������� ������'9K ]o������ ��#5Ga�k }�������� //1/C/U/g/y/�/ �/�/�/�/�/�/	?? -???YK?u?�?�?� ��?�?�?OO)O;O MO_OqO�O�O�O�O�O �O�O__%_7_Q?c? m__�_�_�?�_�_�_ �_o!o3oEoWoio{o �o�o�o�o�o�o�o /�_[_ew�� �_������+� =�O�a�s��������� ͏ߏ���'�9�S ]�o��������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��1�K�9�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�C�� �$ENETM�ODE 1n����  
S�S�N�p߂�R��OATCFG �o�������C���DAT�A 1p_��М.��*��*���!�3�E�T�dT�u몱M�y��������� ������E�W�i�{� �������=����� /A����w�� ����]o+ =Oas��� ���//��K/�]/o/�/�/�/�-R�RPOST_LO��	r��C%
���/??�/?Q�RROR_P-R� %_�%4/q?�@8TABLE  _����?�?�?�+�RSEV_NUM� n�  ��i�@�!_AUT�O_ENB  ���g�@4_NOA �s_ہ�B W *�`@�`@�`@	�`@@+_@yO�O�O�9DFLTR%O7FH�ISCE!g�2K_A�LM 1t_� e�C$`LM�+�O�9_K_]_o_�_�_�O_\�2?@  _�^A����ZR�TCP_V_ER !_�!`?ޣ_$EXT� _R�EQ�F�0I*cSsIZ3o%dSTKPi�NE�'bTOL�  E!Dz�B��A %d_BWD��P�`�F�a�ҢcDI�a u���'��E!�kSTEP�o�oR�>�`OP_DOroP��FDR_GRP s1v_��Ad 	�_xp��aps�Y�q�'�M"����l��T� ����vas��}��tA
�A�I�ZA$@�����{��{/��?��e�P���t����}?���W@/Ơ@�9�?��ܷ�
? F@ �qԁE!@	���R��`��B�-�f�Q�A@�p���@S33��P�@ ����O�؟�ap� ��ŜapG�  (�Fg�fC�8R4��ȝ?�΀Q�Ǟ6��X�x��875t���5���5`�+�ȟH ������%V��ArEATURE �w���`���LR Hand�lingTool� �E"Eng�lish Dictionary���Multi La�nguage (�CHIN)�&�K�ANA/�4D S�t�ard���A�nalog I/�O^�g�gle S�hiftz�uto� Softwar�e Update���matic B�ackup�ͱg�round Ed�it���Came�rau�Fy�Com�mon caliOb UI��n���Monitor�(�tr�Reli�ab����DHCP���Data A�cquis7�`�iagnosɱr�z˿isplay�L�icens^�d�o�cument V�ieweC�b�ua�l Check ?Safety#���?hanced#�����s��Fr����xt. DIO 3�sfi��D�end�ErrB�L��`�8�%s_�rp�O� �`��FCTN Men�u�v^ò�TP ;In��fac�����GigE�����p� Mask Ex�c�'���HT��Proxy Sv���#�igh-Spe�Skiҳ#��SпmmunicȰonsZ�ur�С�u��v���connecwt 2��ncr�Џstru	����e�����J��0�KAREL Cmd. �~��Run-Ti@��Env���el u+̰sʰS/W���������v�Book�(System)��MACROs,~Q�/Offse���0�HSв�s�5�MR�<�8®�M����R�l���MechStoEp/�t����0�iq҄�� x�r�ʰ��o}d��witch.���.��TOpt1mf��0�fi����g��0�-T���PCM fun��:�	a��tiz���o��Regii�r,u��ri��F�4�s�Num Sel���O>� Adju�e�Jw���tat�u0�����RDM� Robot�s�cove��ea��@�Freq Awnlyu�Rem���S�nU���Ser�voS�A ��SNPgX b1�SN���Cli��_.��Li#br�/� � �K&oN�t��ssag�0��P ����a���P/I���%MIL�IB?�"P Fi�rm���.P��Acyc��TPTXo��$eln��?�!���-orqu��i�mulaA���6uH Pa*��.�\�b�&/�ev.�%��r�i��t?USR �EVNTO-@ne�xcept� n���(E9�{�VC�rp�g���V���B<?�E4�+�KSr SCn5�OgSGE�O�EUIa�?Web Pl�^�=!��ET7������ZDT Appln�<�QEOAT�!Ѵ���iPj�ax)�_ Grid����]�_iR�B.U�f����O��RX-10i�A�_m�ll Sm�oothU���c�s�cii/�vLoa9d��tjUpl�`���toS��0rityAvoidM,��sW�t�0g`	�yc����;@�c�CS�/�. c�� xJo=tL�r x��u��� xc��abo���RL�0>�2Y��or��O�0�S�gFit��{tl��nt���wHMI 7Dev�� (S!m� d��in�#?�
�ߞ�sswo\���ROS Eth(��a�!��$�[L%�g 0�b�L%dhUpvE!��%[�t �НiR�s��{�64MB �DRAM��FR�O#����l<f Fl�H����6m �aZ�o�pq���e``v��sh����Ɨc�Õ��Yp�6؜ty��sa�)�r'��j"~ 1.z�pq/sJs�`d� �vx��� 2�ap�pornv���<"V�q�T1*�F1C/��E�Fs=���Hel�U!��Ty-p��FCE h��v�R@St�{����lu�A $ꃨPG j����Rj��No �m �c߷ dOL�;�Sup���0OOPC-UJk"�T�`��5��j��cr.p�lu� �����quir��� Om���%�T0.
���est~L%IMPLE ���VJ'S;�eq�te!x��dhz�I(p��[B�?CPP���E����bTeaH �9���Drtu���v�Y����4���UIFg�p�onsRfstdp�nKe SWIM�EST f� F01ᚥ� bC�:�L�y� p���������	�  ��?�6�H�u�l�~� ������������ ;2Dqhz�� ����
7. @mdv���� ���/3/*/</i/ `/r/�/�/�/�/�/�/ �/?/?&?8?e?\?n? �?�?�?�?�?�?�?�? +O"O4OaOXOjO�O�O �O�O�O�O�O�O'__ 0_]_T_f_�_�_�_�_ �_�_�_�_#oo,oYo Pobo�o�o�o�o�o�o �o�o(UL^ �������� ��$�Q�H�Z���~� �������؏���  �M�D�V���z����� ��ݟԟ��
��I� @�R��v�������ٯ Я����E�<�N� {�r�������տ̿޿ ���A�8�J�w�n� �ϒϤ���������� �=�4�F�s�j�|ߎ� ������������9� 0�B�o�f�x����� ���������5�,�>� k�b�t����������� ����1(:g^ p�������  -$6cZl~ �������)/  /2/_/V/h/z/�/�/ �/�/�/�/�/%??.? [?R?d?v?�?�?�?�? �?�?�?!OO*OWONO `OrO�O�O�O�O�O�O �O__&_S_J_\_n_ �_�_�_�_�_�_�_o o"oOoFoXojo|o�o �o�o�o�o�o KBTfx��� ������G�>� P�b�t�������׏Ώ �����C�:�L�^� p�������ӟʟܟ	�  ��?�6�H�Z�l��� ����ϯƯد���� ;�2�D�V�h������� ˿¿Կ���
�7�.� @�R�dϑψϚ��Ͼ� �������3�*�<�N� `ߍ߄ߖ��ߺ����� ���/�&�8�J�\�� ������������� +�"�4�F�X���|��� ������������' 0BT�x��� ����#,> P}t����� ��//(/:/L/y/�p/�/�/�/�*  H551�#Z�!2�(39�(0�%�R782�'56J�614�%ATUP�'6545'86�%V�CAM�%CUIFv'728c6NRE6�52V6R63�&RwSCH�%LIC�6�DOCV�6CSUv6866J6026�EIOC�746R{69V6ESET?7vU7J7U7R68�&�MASK�%PRXuYo87�&OCOH�3?86@&83^FJq6%8 :�GLCHFF�OPLG?70vFM�HCRGFS�GMA]T�6MCS>80"G{5526MDSW+WviGOPiGMPRjFt�0�H06PCMn7�5qW@26�@�G51�J751�X0J6PR�SG69^FFRD�b6FREQ6MC�N�&97SNBA��7�GSHLBfM�1g�0X26HTC�>6TMIL86T{PA�6TPTXcf#ELf�@�7870��&J95z6TUT�jFUEVFUEC�FFUFRb6VCC��hO�FVIPnfC;SC�fCSG�6�0�I�%WEB>6HTT>6R6�8�h;0Fv�CG]wIGEwIP�GS�vRCnfDG�iGH7�X6�'R7�	GR�XR51�86JvH2vH5V6�0JXʮX6z7L=i�'J8m7"G87�G83J6�R55vF@26R6�4�g5��R6�GR[84��79�H4z6�S5]GJ76^FD�0626F �RTS�fCRDFCRX�jFCLIZXI7CMqS�6S�>6STYng6)WCTO>6�0�7q7�7�0z6ORS�F�7@6FCB�6FC�F�WCH>6FCRnFFCI�vFC�G�J�pOWG*�M�XNOM�6OLWKP�6{OP��SENDGF�LU�FCPR�WL�	wS��C�8ETS�^�T��0zgCP�6T�E%�S60�&FVmR�6IN�WIHag�IPNnfGene �$�(1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�q߃ߕߧ߹��� ������%�7�I�[� m����������� ���!�3�E�W�i�{� �������������� /ASew�� �����+ =Oas���� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ m������ ��!�3�E�W�i�{� ������ÏՏ���� �/�A�S�e�w����� ����џ�����+� =�O�a�s����������ͩ  H�551ϧ�2�3�9��0�R782z�5�J614��ATUP?�545z?�6�VCAM�oCUIF?�28���NRE�52~�R{63�RSCH��LIC��DOCVn��CSU�86��J60N�EIOC���4.�R69~�EgSET_�}�J7}��R68�MASK^�PRXY��7�OCO�3_�.���>�3��J6=����LCH��OPLGz_�0��MHCR���S}�MAT��MC�S^�0��55N�MgDSW����OP��GMPR��۰.�0�PCM��5M��N�l��.�51n�51���0n�PRS~�69���FRD��FRE]Q�MCN�9��SNBAϻ�SH�LB�MM�۰��2��HTC^�TMI�L��TPAN�T7PTX��EL����.�8-�+��J95TUT��UEV�~�UEC��UFR���VCC^O��V�IP��CSC��C�SG���I�WE�B^�HTT^�R6�ͼ��[��
CG�I�G�IPGSRmC��DG��H7m�6�R7m�R��R�51^�6��2��5�~��J�ܞ�6��L�]��J87��87v.�83n�R55��\k�N�R645�+�R6��R84n+7�9�4��S5��J�76��D06N�F�<RTS.�CRD�~�CRX��CLI.�m�CMSN�{0^��STY��6��CTO^��N�7-�˰���ORS�ګ��FC�BN�FCF��CH�^�FCR~�FCI�>FC��J�G��M��NOMN�O�L����OP]KS�END��LU~�C�PR��LmS�<C�ETS�K|<;����CP��TE=;S6�0�FVRN�INv��IH��IPN��Gene�Ψ�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o���� �����#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W� i�{ߍߟ߱������� ����/�A�S�e�w� ������������ �+�=�O�a�s����� ����������' 9K]o���� ����#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G��Y�k�}�������ů � נSTD~ҤLANG� ���0�B�T�f�x� ��������ҿ���� �,�>�P�b�tφϘ� �ϼ���������(� :�L�^�p߂ߔߦ߸� ������ ��$�6�H� Z�l�~�������� ����� �2�D�V�h��z�������RBT�OPTN������ 	-?Qcu��������DPN�);M_ q������� //%/7/I/[/m// �/�/�/�/�/�/�/??ted �ʨ 9?K?]?o?�?�?�?�? �?�?�?�?O#O5OGO YOkO}O�O�O�O�O�O �O�O__1_C_U_g_ y_�_�_�_�_�_�_�_ 	oo-o?oQocouo�o �o�o�o�o�o�o );M_q��� ������%�7� I�[�m��������Ǐ ُ����!�3�E�W� i�{�������ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳����� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q��� ����%7 I[m��������/!/3/E/  �N/l/~/�/�/�/��-99�%�$F�EAT_ADD �?	����!~0  	�( ??/?A?S?e?w?�? �?�?�?�?�?�?OO +O=OOOaOsO�O�O�O �O�O�O�O__'_9_ K_]_o_�_�_�_�_�_ �_�_�_o#o5oGoYo ko}o�o�o�o�o�o�o �o1CUgy �������	� �-�?�Q�c�u����� ����Ϗ����)� ;�M�_�q��������� ˟ݟ���%�7�I� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o�������������$DEMO �w�)   �(4�*�<�i�`�r� �������������� /&8e\n�� ������+" 4aXj���� ����'//0/]/ T/f/�/�/�/�/�/�/ �/�/#??,?Y?P?b? �?�?�?�?�?�?�?�? OO(OUOLO^O�O�O �O�O�O�O�O�O__ $_Q_H_Z_�_~_�_�_ �_�_�_�_oo oMo DoVo�ozo�o�o�o�o �o�o
I@R v������ ���E�<�N�{�r� ��������ԏޏ�� �A�8�J�w�n����� ����Пڟ����=� 4�F�s�j�|������� ̯֯����9�0�B� o�f�x�������ȿҿ �����5�,�>�k�b� tϡϘϪ��������� �1�(�:�g�^�pߝ� �ߦ��������� �-� $�6�c�Z�l���� ����������)� �2� _�V�h����������� ������%.[R d������� �!*WN`� �������/ /&/S/J/\/�/�/�/ �/�/�/�/�/??"? O?F?X?�?|?�?�?�? �?�?�?OOOKOBO TO�OxO�O�O�O�O�O �O___G_>_P_}_ t_�_�_�_�_�_�_o ooCo:oLoyopo�o �o�o�o�o�o	  ?6Hul~�� ������;�2� D�q�h�z�����ˏ ԏ���
�7�.�@�m� d�v�����ǟ��П�� ���3�*�<�i�`�r� ����ï��̯���� /�&�8�e�\�n����� ����ȿ�����+�"� 4�a�X�jτώϻϲ� ��������'��0�]� T�f߀ߊ߷߮����� ����#��,�Y�P�b� |����������� ��(�U�L�^�x��� ������������ $QHZt~�� ���� M DVpz���� ��/
//I/@/R/ l/v/�/�/�/�/�/�/ ???E?<?N?h?r? �?�?�?�?�?�?OO OAO8OJOdOnO�O�O �O�O�O�O_�O_=_ 4_F_`_j_�_�_�_�_ �_�_o�_o9o0oBo \ofo�o�o�o�o�o�o �o�o5,>Xb �������� �1�(�:�T�^����� ������ʏ��� �-� $�6�P�Z���~����� ��Ɵ����)� �2� L�V���z�������¯ ����%��.�H�R� �v����������� ��!��*�D�N�{�r� �ϱϨϺ�������� �&�@�J�w�n߀߭� �߶���������"� <�F�s�j�|���� ���������8�B� o�f�x����������� ��4>kb t������ 0:g^p� �����	/ // ,/6/c/Z/l/�/�/�/ �/�/�/?�/?(?2? _?V?h?�?�?�?�?�? �?O�?
O$O.O[ORO dO�O�O�O�O�O�O�O �O_ _*_W_N_`_�_ �_�_�_�_�_�_�_o o&oSoJo\o�o�o�o��o�o�o�o�o}  x.@Rd v������� ��*�<�N�`�r��� ������̏ޏ���� &�8�J�\�n������� ��ȟڟ����"�4� F�X�j�|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������>�  �� 2�D�V�h�z������� ��������
.@ Rdv����� ��*<N` r������� //&/8/J/\/n/�/ �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�? �?�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� � 2�D�V�h�z������� ԏ���
��.�@� R�d�v���������П �����*�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮��� ��������,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZl~� ������  2DVhz��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|������������� ��6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x���� ����������,�>� P�b�t����������� ����(:L^ p�������  $6HZl~ �������/  /2/D/V/h/z/�/�/ �/�/�/�/�/
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8_J_\_n_ �_�_�_�_�_�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�o�oy��$FEAT_D�EMOIN  V#t�Np�$p6t_INDEXC{Rq��6pILECOM�P x�����qQr1uzpS�ETUP2 y��u�r�  �N �qws_AP2�BCK 1z�y  �)x��{%� �$p�p�K� !u�w����*���я `������+���O�ޏ s������8�͟ߟn� ���'���4�]�쟁� �����F�ۯj���� ��5�įY�k������ ��B����x�Ϝ�1� C�ҿg����ϝ�,��� P����φ�ߪ�?��� L�u�ߙ�(߽���^� �߂��)��M���q� ����6���Z���� ��%���I�[����� ����D���h����� 3��W��d�� @��v�/A �e���*�N@�r�/�y�pP�� 2�p*.V1R /j/�*m/�/`��/�/�T PC�/|�/�FR6:�/">�/>?�+Tbpb? t?5_?�<Ep/?�?��*.FW/�?�	�3�?"L�?FO�;STMQO{O20gO�M5O�O�;H�O�O�G��O�O�OO_�:GIF Y_�_�Eo_,_>_�_�:JPG�_o�E�_�_�_Wo�*JSao�o��cxo5o%
Ja�vaScript�o�_CS�o�F�o��o %Casc�ading St�yle Shee�ts:�
ARGNAME.DTi
��@\};�a�t��j�pDISP	*���t���q�4�B��CLLB�.ZI_��@:\҅�\��Ɖ�aCo�llaboƏr�
?PANEL1�O ��s	�C��qiPen�dant PanelJ��	9�:�"��5���R�d����2 ?�(�3��ԟ�{���2ß������X�j����3G�0�3��ܯ�����3˯������`�r���4O�8�3�&�����φ�4ӿ�Ϸ���h�z��vtTPEINS.XML��=�:\)��ϥqCu�stom Too�lbarj��yPA?SSWORD����FRS7���n��Password Config�� �7���0�m���� � ����V���z��!��� E���i���
���.��� R���������AS ��w��<�` ���+�O�H ��8��n/ �'/9/�]/��// "/�/F/�/j/�/?�/ 5?�/Y?k?�/�??�? �?T?�?x?O�?�?CO �?gO�?`O�O,O�OPO �O�O�O_�O?_Q_�O u__�_(_:_�_^_�_ �_�_)o�_Mo�_qo�o o�o6o�o�olo�o %�o�o[�ox �D�h���3� �W�i�������@� R��v�����A�Џ e�􏉟��*���N�� �������=�̟ޟs� ���&���ͯ\�񯀯 �'���K�گo�������4�ɿX�j������$FILE_DG�BCK 1z������� < �)
S�UMMARY.D9G	���MD:=�}����Diag Summary~���CONSLOG@s�V�h���ߐ��sole lo����	TPACCN���\�%D߁ߌ�T�P Accoun�tin#ߋ�FR�6:IPKDMPO.ZIP�߹�
����ŝ�Excep�tion
��i�MEMCHECKw����lύ��Mem�ory Data|���:n )x�RIPE��f�x����%�� Pa?cket L"���L�$�K���ST�AT��� ��� �%)�Stat�us��F�	FTP�����|������m�ment TBD�F� >I)E?THERNE_����L�]���Eth�ern2��fig�ura)DCSVRF������  veri?fy all"��(4�DIF�F��#�9d�iff�ZL�� CHG01���)/���Q/\2��2 ///�/�N/`/��3�/�/�/1? ��/X?�&VTRNDIAG.LS]?�? ?�?��u1 O�pe�4� ��no�stic��'Ͽ)VDEVy2D�AT�?�?�?�?���Vis�1Devisce�?�;IMGy2���O&O�O"�QDI�mag]O�;UP�@ESO�OFR�S:\_B]��U�pdates L�istB_���@FLEXEVEN�КO�O�_���Q UIF Ev55���-vZ)
PS�RBWLD.CM��_��-R	oD_�P�S_ROBOWEyL;�:GIG���o�_�o��Gig�E�H�_�N�@��)�aHADOW��o�o�oO��Sh�adow Cha�nge����.dt~rRCMERRG�,>����pCFG ErrorW@�tailv MA��S�CMSGLIB���Y��b�̱�bPic ���)E�ZD�o��B��׏��ZD�`ad�y�� rNOT�I���ȏ]���N?otific����,�AG)CRSENSPK�O�����\���� C�R_ؑOR_PEAK柍�.�@��d� 翈������M��q� ����<�˯`��� ��%���̿����� ��%�J�ٿn����Ϥ� 3���W���{ύ�"߱� F�X��|�ߠ�/߱� ��e��߉��0��T� ��x����=����� �����,���=�b��� �������K���o� ����:��^p+� #�G��}� 6H�l��1 �U��� /�D/ �U/z/	/�/-/�/�/ c/�/�/?�/�/R?�/ v?�?C?�?;?�?_?�? O�?*O�?NO`O�?�O O�O7OIO�OmO__ �O8_�O\_�Om_�_!_ �_E_�_�_{_o�_4o �_�_jo�_�o�o[o�o So�owo�o�oB�o fx�+�Oa ���,��P��t� �����9�Ώ]��� ��(���L�ۏ폂�� ����s�ܟk� ���� 6�şZ��~�������C�دg�y����$�FILE_FRS�PRT  ���������'�MDONLY� 1z;��� 
 ���~�˯��� ��ؿ������ �2��� V��zό�ϰ�?��� ��u�
ߙ�.߽�;�d� �ψ�߬߾�M���q� ���<���`�r�� ��%��I������� ��8�J���n������ 3���W�������"���F��S|%�VIS�BCKY�C�h�*�.VD��; F�R:\� ION\�DATA\�^�; Vision� VD file �ASiwa� *��`��/+/ �O/�s///�/8/ �/�/�/?�/'?�/8? ]?�/�??�?�?F?�? j?�?�?�?5O�?YOkO &O�OO�OBO�O�OxO _�O1_C_�Og_�O�_�_,_�_!�LUI_�CONFIG �{;���[ $ �S^��V#o5o�GoYoko}o�i`|x �_�o�o�o�o�o|�o 0BTfx�� ������,�>� P�b�t��������Ώ ��򏉏�(�:�L�^� p��������ʟܟ� ���$�6�H�Z�l�� ������Ưدꯁ��  �2�D�V�h������� ��¿Կk��
��.� @�R��vψϚϬϾ� ��g�����*�<�N� ��r߄ߖߨߺ���c� ����&�8�J���n� �������_����� �"�4�F���j�|��� ������[����� 0��Afx��� E���,� Pbt���A� ��//(/�L/^/ p/�/�/�/=/�/�/�/  ??$?�/H?Z?l?~? �?�?9?�?�?�?�?O  O�?DOVOhOzO�O#O �O�O�O�O�O
_�O._ @_R_d_v_�__�_�_ �_�_�_o�_*o<oNo `oro�oo�o�o�o�o �o�o&8J\n ���������tRobot �Speed 100%�:�L�^�p���>�r  x������$FLUI_D�ATA |����Ł��q��RESULT� 3}Ņ� ��T�/wi�zard/gui�ded/step�s/Expert ��%�7�I�[�m����ࣟ��ǟٟ��C�ontinue �with G�ance�"�4�F�X� j�|�������į֯� ��-��Ņ�0 ��p�ǃlƁ'����ps� r���������̿޿� ��&�8����_�q� �ϕϧϹ�������� �%�7ߏuт�q'���+�=�+M�cllb��ToolSet~��g/Dist�Work@������ �%�7�I�[�m���.0��������� ����%�7�I�[�m�����w{ݐqo߁�:?�&M�rip����Num/NewFram�+=Oa s��������0x��
.@ Rdv�������p��c�/��E��M���imeUS/DST�y/�/�/ �/�/�/�/�/	??-?~�Enabl a?s?�?�?�?�?�?�?��?OO'O9O����/sO5/G/Y&24 d/�O�O�O�O_#_5_ G_Y_k_}_<?N?�_�_ �_�_�_oo1oCoUo goyo�oJO\OnO�OB�|��
�ditor�o /ASew������ Tou�ch Panel� s (reco/mmen�)�$� 6�H�Z�l�~�������Ə؏� ��o�o���o�oracces `�p���������ʟܟ�� ��$�?�Co�nnect to Netw��g�y� ��������ӯ���	��-�싘O���#���!E�pIntr�oduction 6�˿ݿ���%�7� I�[�m���u��ϰ� ��������
��.�@� R�d�v߈����]���0����Us�_#� 5�G�Y�k�}���������q1���� %�7�I�[�m�������������a
�����H������)����A��ve���{����������
0xFE/^p� ������ //$/2*�c.L/ �2D/Macro>�s/New�"_� �/�/�/??(?:?L?�^?p?�?�0x0 �?�?�?�?�?�?OO )O;OMO_OqO�OB&��]/�O�/�,�/�+�"Open�#_5_G_ Y_k_}_�_�_�_�_�? ���_oo1oCoUogo yo�o�o�o�o�o����ȶO�O��-�O�OoClos�w�����������_2+�Q�c�u������� ��Ϗ����)��o �iR���=���SetMethod.���ӟ���	���-�?�Q�c�u�8��c�[������W�n�𒼐ړ������̯ ޯ���&�8�J�\�n��� ="iqr�O�a�s���$����tr�aightOffset���,�>�P� b�tφϘϪϼ���=�X�g����g������,�>�P� b�t߆ߘߪ߼��ߍ�al�����ѿ�%�S�M�X��o��� ������������#�>.0<�'�Q�c� u���������������H)A��h ��+�=�O�Y*�� ��/ASe w6������� //+/=/O/a/s/2�DV�/z��tZ ~/?)?;?M?_?q?�?��?�?�?�?�117.762��?O O1OCOUOgOyO�O�O�O�O�/�/�$B놑%�/�/׺)�/��RotationIWW�Oo_�_�_�_�_�_��_�_�_o�?180�Ko]ooo�o�o�o �o�o�o�o�o#�OXC3�_%_7_I_onP&���� ��/�A�S�e�$o� ������я����� +�=�O�a�s�2�/�/0hz��nRz�� )�;�M�_�q���������x�-99o�� �(�:�L�^�p�����`����ʿ����´��仟�,"ݟ�tp3�Zdir/Tp3zοd�vψϚϬϾ� ���������?<�N� `�r߄ߖߨߺ����� ����ӿ��O���� +1��Meas�urement/Straigh? ����������+�=� O�a� �2ߗ������� ����'9K]�o.�@�R�d�v��/�We��Nums/New�sv' 9K]o����v�0x��� // $/6/H/Z/l/~/�/�/�/�/-`��)���#�.��Tool�Use�/l?~?�? �?�?�?�?�?�?O)j1OAOSOeOwO�O �O�O�O�O�O�O__-a
�/���/Y_?<-?�PartR?�_ �_�_�_�_o#o5oGoYoko*B2oo�o�o�o �o�o�o%7I[m,_��K_��9(�_�s/G��� r� �2�D�V�h�z�0��������� ����0�B�T�f�x� ����������{}��#�)��yPayload1Cm� b�t���������ί�������p��[�c�Ȃ��c-���L�^�p��� ������ʿܿ� ��}�ٟ�/5���3� �Y϶�����������"�4�F�X�j��10׏�ߤ߶������� ���"�4�F�X�j�՟W�A ��[���=�2O���,�>�P�b��t���������'�����5��� $6 HZl~���� ��C����}P&�����Advanced �\n���������/{�0x ��:/L/^/p/�/�/�/��/�/�/�/ ??u� ��1?u�%%���Mass/Center�1?�?�?�? �?�?	OO-O?OQOcO ҏ�O�O�O�O�O�O�O __)_;_M___v�0?`�_f?��?ss�� j_oo+o=oOoaoso �o�o�ohOzO�o�o '9K]o�����v_�_�_�_�[,��_��G.c�2�XX �^�p���������ʏ ܏� ��o�o6�H�Z� l�~�������Ɵ؟� ��������'�9�sY���į֯� ����0�B�T��%� ��������ҿ���� �,�>�P�b�!�3�E�0W�i�{���sZf�� �*�<�N�`�r߄ߖ� ��g�y�������&� 8�J�\�n����� uχϙϫ�.����p�P�\L�[�m���� ���������������� 3EWi{��� ����������0 ��$�6�rt��� ����	//-/?/ Q/"�/�/�/�/�/ �/�/??)?;?M?_?�0BTfx�rt��OO'O9OKO]O oO�O�O�Od/v/�O�O �O_#_5_G_Y_k_}_ �_�_�_r?�?�?�?����<TCPVeri�fy/2cMethod�_Vohozo�o�o��o�o�o�o�o�LD�irect Entry8J\n ����������H�_'��_�_j'o+ofyJ�����ȏ ڏ����"�4�F�X� �O|�������ğ֟� ����0�B�T��_A�`�_��[�m��fy� ��
��.�@�R�d�v� ������k�п���� �*�<�N�`�rτϖ� ��g������ϯ���ӯfy�?L�^�p߂ߔ߀�߸������� ￰117.762ǿ /�A�S�e�w���������������B�%������/mW��������������1CU�80 ÿ������ �!3EW�D��C39�G�Y�k�}�P Z�//+/=/O/a/ s/�/�/�/���/�/�/ ??'?9?K?]?o?�? �?�?d���Ϛ���yR�?IO[OmOO �O�O�O�O�O�O�O�-9m&_8_J_\_n_ �_�_�_�_�_�_�_�_��?�9´�?�?L*�O#OfyMean o�o�o�o�o�o�o0B_*gtS� �������� "�4�F�oou�3oEobJ)eowo�`axV� ���)�;�M�_�q� ����Tf˟ݟ�� �%�7�I�[�m����@��b�������K"���ˁIntroductio�o?�Q�c� u���������Ͽ�� �%�2�$�6�H�Z�l� ~ϐϢϴ��������ς� ��ѯ���B �ˀ ߇ߙ߽߫��� ������)�;�M�� q����������� ��%�7�I��6�,��>� M#a�file�2/cyclep{owƆmodeT� ����1CUg�y���#�z��b�g�X�^�[�g���� 0BTfx��Z�&e�!� ������La�uid�edȄSafety�5/G/Y/k/}/�/ �/�/�/�/�/T�?? 1?C?U?g?y?�?�?�? �?�?�?�?g�g���O�����/don ���O�O�O�O�O�O�O _ _2_D_?h_z_�_ �_�_�_�_�_�_
oo .o@o�?O#OmoGO/ȄReg,��o�o�o "4FXj|�~��EuropO �����#�5�G��Y�k�}�����abz c�o}o�oML�o �Timez}@EU ��5�G�Y�k�}�����೟şן韨wEE�T Ea rn �sa�o+�=�O�a�s� ��������ͯ߯񯰇�c`�ߏя㏡o��24���������� Ϳ߿���'�9�P_ ]�oρϓϥϷ����� �����#�5�G�^o��*�<�RO`�24/c?urrentL��� ����)�;�M�_�q�����s29-N�OV-25 17:29 �������� ��*�<�N�`�r�����_����yߋߝ�y �߿�Year�� 2DVhz��������v2025�*<N`r�������� y
����  ����-/��!��Month��/�/�/�/�/��/�/??)?;?�u11C?j?|?�?�?�? �?�?�?�?OO0OBO/' /�O�U/��DayFO�O�O�O _!_3_E_W_i_{_�_L829�_�_�_�_�_ oo*o<oNo`oro�o�oUOgHsO�o���O��Hou -?Q cu������L97��$�6�H�Z� l�~�������Ə؏�D�ogH�o)���"�o>g(inute� ������̟ޟ��� &�8��_\�n������� ��ȯگ����"�4�@���o-�;�Q Q�~��NetDonr� ѿ�����+�=�O� a�sυ��nA�ϻ��� ������'�9�K�]�o߁ߓ�W�W����� ��O"��	��-�?�Q� c�u��������� ����)�;�M�_�q��������������I� ���߽�����Xj |������� 0��Tfx� ������// ,/����!3E�/ �/�/�/�/??(?:? L?^?p?�?A�?�?�? �?�? OO$O6OHOZO lO~O�OO/a/s/�/�/ �O_ _2_D_V_h_z_ �_�_�_�_�_�?�_
o o.o@oRodovo�o�o �o�o�o�o�O�O�O�O���W�Summary�ov����� ����*��_N�`� r���������̏ޏ�� ��&�8���	-�?��RobotOp<�ʟܟ� ��$� 6�H�Z�l�~�=����� Ưد���� �2�D� V�h�z���O�O�a�諿����&��cll�bWtToolSe�tting�Off��(�:�L�^�pς���Ϧϸ����ϛ�1 ����)�;�M�_�q߀�ߕߧ߹����ߣ�
@�iͷK���%��n��{��������������/���2 3�Y�k�}��������� ������1���Q�q��.E�/��SpeedLim?it/Max�6 ��� 2DV�hz��	1000.�0����� �/!/3/E/W/i/{/�+IsDz  �gy����Val�/,?>?P?b?t?�? �?�?�?�?��OO (O:OLO^OpO�O�O�O �O�O�O�/�/�/�/����//Intro?ductioi�p_ �_�_�_�_�_�_�_ o o$o��HoZolo~o�o �o�o�o�o�o�o @2M���M'_��A_�� lectWork4�������/�A�S�e�w�6iL�ightwe�� >�qpiece���� Ϗ����)�;�M��_�q���  Er��Sew�4�/�Load�NotOHW_l��W�W�� ��.�@�R�d�v�����p����Я;d.3�? ���"�4�F�X�j�|��������Ŀֿ�OÙ>G�����ɟ7�8�����CenterMassڿ�ϘϪ� ����������(�� �?Q�c�u߇ߙ߽߫� ��������)���C���3Z5=�O�a�omml�.������� ��1�C�U�g�y�<c�EOAT w/o par����� ������
.@Rdv;xA﫟�w� �/����+=O as�����8� �//'/9/K/]/o/ �/�/�/�/�/4�X�����2��g� n?�?�?�?�?�?�?�? �?O"O�FOXOjO|O �O�O�O�O�O�O�O_�_�/�/?c_%?�/ 9?K?���_�_�_�_
o o.o@oRodovo���_ �o�o�o�o�o* <N`r�C_��y_�+�_���"� 4�F�X�j�|�������ď�h10;O��� �,�>�P�b�t�����`����Ο9_�yA Y_ �}_��~a?k�}��� ����ůׯ����� 6OC�U�g�y������� ��ӿ���	��ڟ�V_`�"�,5�G��_�� ��������*�<�N��`�r߉b�cith �o�߷���������� #�5�G�Y�k�<Ϧ���r��6��/� C�ontactSt�opInvali�dArea/�PlusZz�$�6�H� Z�l�~���������ݏ ���� 2DVh z����-ϓ�������7�����Min�v���� ���//��</N/ `/r/�/�/�/�/�/�/ �/??���b��51C�XY	�XY"?�?�?�?OO %O7OIO[OmO,/�O�O �O�O�O�O�O_!_3_ E_W_i_(?:?L?^?p?���)�?��NotHW_l�o!o3o EoWoio{o�o�o�o�o �AR��o�o&8 J\n�������P�_����_�� �_U����\�n����� ����ȏڏ�����o 4�F�X�j�|������� ğ֟��������9���� -��1SpeedLimio ��ïկ�����/� A�S�e�$��������� ѿ�����+�=�Oπa�s�2�D���h��S<����Modet�� �)�;�M�_�q߃ߕ���߹�|GDo n�ot Use (�Recommended)�� ��$� 6�H�Z�l�~����*����"���ϡ� ���\��9�K�]�o��� �������������� |�5GYk}��������yH �����7�#��� �����//*/ </N/`/�/�/�/�/ �/�/�/??&?8?J? \?-?Qcu�? �?�?O"O4OFOXOjO |O�O�O�Oq/�O�O�O __0_B_T_f_x_�_ �_�_�_?�?�?�?�? ,o>oPoboto�o�o�o �o�o�o�o�O(: L^p����� �� ���_�_�_o o~�������Ə؏� ��� �2�D�V�g� ������ԟ���
� �.�@�R�d�#���G� Y�k�Я�����*� <�N�`�r��������� ˯޿���&�8�J� \�nπϒϤ϶�u��� ������"�4�F�X�j� |ߎߠ߲��������� �˿0�B�T�f�x�� �������������� )���M��������� ��������(: L^����� �� $6HZ �{=��a�u�� �/ /2/D/V/h/z/ �/�/�/o�/�/�/
? ?.?@?R?d?v?�?�?��?k���?���/wizard/�cllb/ste�ps/Summary�?HOZOlO~O�O �O�O�O�O�O�O�/ _ 2_D_V_h_z_�_�_�_@�_�_�_�_
o�2�7��?�?�?�(O/C�onfigura�tionCompleteo�o�o�o �o�o(:L^ _�������� ��$�6�H�Z��6�#o5o�Yo�3qo/�SignalNumberAssـ�ment/SPI ރd�	��-�?�Q�c�`u�������ju1�� ٟ����!�3�E�W�@i�{��������1
�9 ��a���2ŏ׏�D�U�g�y����� ����ӿ������-� ?�Q�c�uχϙϫϽ� �������į֯�����
ߐߢߴ��� ������� �2�D�V� mz������������
��.�@�R��: ߉�{�U�������� &8J\n� ��c����� "4FXj|���?�?�������/ ./@/R/d/v/�/�/�/ �/�/�/�/�?*?<? N?`?r?�?�?�?�?�? �?�?O���GO	/ nO�O�O�O�O�O�O�O �O_"_4_F_?W_|_ �_�_�_�_�_�_�_o o0oBoToOuo7O�o [O�o�o�o�o, >Pbt����o �����(�:�L� ^�p�������eoǏ�o 돭o�$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ������ ۏ=����v������� ��п�����*�<� N��rτϖϨϺ��� ������&�8�J�	� k�-��ߡ�e������� ���"�4�F�X�j�|� ���_���������� �0�B�T�f�x����� [ߥ��������, >Pbt���� �����(:L ^p������ �������/E/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?h?z?�? �?�?�?�?�?�?
OO .O@O�/#/5/�OY/ �O�O�O�O__*_<_ N_`_r_�_�_U?�_�_ �_�_oo&o8oJo\o no�o�o�ocOuO�O�o �O"4FXj| �������_� �0�B�T�f�x����� ����ҏ����o�o�o ;��ob�t��������� Ο�����(�:�� K�p���������ʯܯ � ��$�6�H��i� +���O���ƿؿ��� � �2�D�V�h�zό� �ϯ���������
�� .�@�R�d�v߈ߚ�Y� ��}��ߡ���*�<� N�`�r������� ������&�8�J�\� n��������������� ����1����j| ������� 0B�fx�� �����//,/ >/��_/!�/�/Y�/ �/�/�/??(?:?L? ^?p?�?�?S�?�?�? �? OO$O6OHOZOlO ~O�OO/�/s/�O�O�/ _ _2_D_V_h_z_�_ �_�_�_�_�_�?
oo .o@oRodovo�o�o�o �o�o�o�O�O�O9 �O`r����� ����&�8��_\� n���������ȏڏ� ���"�4��o) ��M��ğ֟���� �0�B�T�f�x���I� ����ү�����,� >�P�b�t�����W�i� {�ݿ����(�:�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ������ߩ� ��Ϳ/��V�h�z�� �����������
�� .���?�d�v������� ��������*< ��]�C��� ��&8J\ n������� �/"/4/F/X/j/|/��/M�/q�/�+�$�FMR2_GRP� 1~�%�� �C4 w B�� 	 � �!?3<0F@ �I?@�+0G�  �q1Fg�fC�8yR}5a=?�  �?��,06�X��2��875t��5����5`+�a=Ag�  �?�;BH�4<_0E@S33!E�,!4COTM0@AjO `>TO�O�O�O�O�O�O _�O2__/_h_S_�_��#�"_CFG ;T32�_�_�_�_��YNO :�
F0.a 3`�\R�M_CHKTYP  �!� 00� ��!ROMI`_MI�NO`�#��{`��:@X� SSB�S���% �6�o�%�c�o�o�UT�P_DEF_OW�  �$3�gI�RCOMN` �$�GENOVRD_�DOpf�-}TH��0rd dJud3t_�ENB 3pRWAVC�#��g�` �A5�o�y_��a<��1J �V�qOU 0�<6aq18r15<x`��?��/�}���͏�#C��3�!���o"��!�>����Br0��49p��o�pSMT��#��y0�`��$�HOSTC�R1��9�`���0 kMC�$
�ȟ��&  27.0z�1�  e�� E�W�i�{��*3������Я������	anonymous	� 7�I�[�m�� ǟ0���������,�	� �-�?�QϘ�uχϙ� ��οh������)� ;߂��Ϧ�������� ��������Z�7�I� [�m����������� �����V�h�zߌߎ� {��ߟ���������.� /ASv���m �����*�<�N� +bO��s��� �����//8� �]/o/�/�/�/�� "$/?X5?G?Y? k?}?��?�?�?�?�? ?B/T/1OCOUOgOyO �/�/�/�O�?�O,?	_ _-_?_O�Ou_�_�_ �_�O�_O�_oo)o ;o�O�O�O�O�_�o�O �o�o�oZ_7I [m�o�_�_������|���ENT� 1�P� P!\�V�  'pD� ��p���h�ɏ��폰� ��ԏ"�G�
�k�.��� R���v�ן�����П 1���U��y�<�N��� r�ӯ�������ޯ� Q�@�u�8���\����� ɿ����ڿ;���_� "σ�Fϧ�j�|��Ϡ�����%���QUI�CC02��!1�92.168.1'.10K�@�1��^� ���D�2�߮���!��!ROUTER�"���!r�I����PCJOGr�M�/!* t�0{�=�?CAMPRT���c!r�����RT;������`� !So�ftware O�perator Panel=�oغ���NAME !~3�!ROBO�����S_CFG 1��3� ��Auto-st�artedidFTPtoI�o�t �o�����- (:]K��� ���Kn"4F#/ Z|:/k/}/�/�/h �/�/�/�/?0/�/C? U?g?y?�?�?Rodovo �o?	OP/-O?OQOcO uO<?�O�O�O�O�OO �O_)_;_M___q_�? �?�?�_�O�_$Ooo %o7o�O[omoo�o�o �_Ho�o�o�o!3 z_�_�_�_�o��_� �����o/�A�S� e�w�������я� ���N`rO���s� �������͟����� �'�9�\�]�🁯�� ����ɯ�"�4�F�H� �|�Y�k�}�����h� ſ׿����0���C� U�g�yϋϝ����� ���	�P�-�?�Q�c� u�<ϙ߽߫������� ���)�;�M�_�����_ERR ����o��PDUSIZW  �^�����>��WRD ?����  guest�ր����%�7�I���S�CD_GROUP� 3� �
�IFT��$PA��OMP�� n��_SH��ED��w $C��COM���TTP_AUTH� 1��� <!�iPendan�U�`'!KAREL:*`i{�KC���� �VISION SETy���'?:�^p���������/CT_RL ���I(��
�'FF�F9E3/��F�RS:DEFAU�LTn,FAN�UC Web Server��\!L" /����,�/�/??�,?>?}�WR_CONFIG �~����cn/�I�DL_CPU_P5C� �B����0w BH�5MIN�<���5GNR_IO�������0HMI�_EDIT ��~�
 ($IP�L_�"_SMPL�GR3 LOSEIOcon 2B��O�OPEN2Bt7H�51 FOXO22�mOO$ bktl�ead-inst�_basicpick_star^I /�O�O__;_&___�J_�_�_Z!($*?uninit�t[ �_�_�_o�_/oo,o r_wo�oto�o�o�o�o��o�o�?$INP�T_SIM_DO��6�:NSTAL�_SCRN�6 ��UzTPMODNT�OLkwT{�!RTY�Jx�1Yv3 ENB�kw��3OLNK 1���������1�C�U�g��rMASTE�0�yH"�q�SLAVE ���H D�uSRA?MCACHE����>5O_CFGǏ�s�߃UO�ۂCM�T�@� �2���YC�LƏ��� _ASG� 1�s7��
  i�������ԟ��� 
��.�@�R�d�v�q��_�NUM����
�ۂIPďևRTR�Y_CN(���gq_�UP�����q��� �ۂ���</  �0I$3��0@gr?}��� ��D�mplGrp/S�ar�e_Conf?ig.stm��������ѿ�ր��� #�5�G�Y��}Ϗϡ� ������f�����1� C�U����ϋߝ߯��� ����t�	��-�?�Q� c��߇�������� p���)�;�M�_�q�  �������������~� %7I[m�� �������! 3EWi{
�� ������//A/ S/e/w/�//�/�/�/ �/�/?�/+?=?O?a? s?�??&?�?�?�?�? OO�?9OKO]OoO�O �O"O�O�O�O�O�O_ �O�OG_Y_k_}_�_�_ 0_�_�_�_�_oo�_ CoUogoyo�o�o,o>o �o�o�o	-�oQ cu���:�� ���)���_�q� ��������H�ݏ�� �%�7�Ə[�m���� ����D�V�����!� 3�E�ԟi�{��������ïR�K�_MEMB�ERS 2�"��2� $"����^������RCA_ACC� 2���   [}}߉��*T�6�]�s�  %T�T�]g�6� T�`w��i��o���I�BUF�001 2�V�=� {�u0  �u0{����Ѫ�������|U���'�U2�=�K�U�Ud�rāĎ�U�īĹ���U������}!ī}����-��:ʲ�J��V��a�}o��{�ĉ�đH�  H�z��z��ԬԷ���zj�z	�z�z�괚!�{)�{�9�{U3�A�M�X�Uf�q�}괊��{!�ǹ2Կ�� ����������	��� ����� �%�)�%� 1�%�9�%�A�%�I�%� Q�%�Y�%�a�%�i�%� q�%�y�%��%��%� ��%��%��%��%� ��걸����������� ����������������pj������u  � ������ �%�)� %�1�%��@�%��P� %�Y���*�h���q��� B���҉��ґ��ҙ� �ҡ��ҩ��ұ��ҹ� ��"����ǹ3��� ���������	���� �'�.)�7�.9�G� .I�W�.Y�g�.i� w�.y�.��. �§�.�·�T����� ������������� �������	��T� �'�&)�7�&@� O�&#X�g���;p� ���ҏ���ҟ��� �ү���ҿ���+��~��CFG 2�V�� 4T���*T��T�<�!!�H�ISѲ�V� ��g� 2025-�11-29T� �T�;  G s#�/�/�/R�XT� U`�$h�$pr$xr$�}�$�/??T�[|�pY(8e)?^? p?�?�?�?�?�?�?�?�T���! R�x��Y"1-07-06�A?.O@OROdOR�^��s#�":�$ �$x����/�O�OP�R�X�H5O
__._@_o  T�#X�{/�p_�_�_�_�J▁H2�O�_�_
oo.o@oRoP����O�oR��QgAY"0-08-31�_�o�o�o�o
gAso0BT\f�boP�g2��o���E^��;� �"v fa#oP�&�8�Ӯ7&��C/U/g*bQdy ��G���ɏ�*!d� ��  �� ��� ��� �ԏ '�9�'?9?������� ��ɟ۟�����6邀Oh�U�g�y���yH6�  [� 8��`8� �� c�@� گ��O�OG�4�F�X�>F_8  ^]P}� h�������ѿ�_�_� �+�=�O�a�s�ao�� �ϗo�o�����'�>x9  _0�[� m��m�������ߜ��	 U@ c�p��ɯ:�L�^�@L�9$��h�z�g*�q y ��������*��� ��� ��� ��� ��� ��G�Y�G�Y��ߡ��� ��������1� ��2���z���yH��)��@6���� �lYk}k��]P ��������� ,/>/P/b/t/�/�/�� ��/����)/?(?:? L?x�/{?�?�?�?�� ���?�?OO�sra� 6B�p6B�j?_OqO�O�q�A_I_CFG� 2��� H�
Cycle T�imeqBu�sywIdl��B�Dmin{�QUp�F�A�Read�GDCow�H�O��Q�C�Count�A	N'um �B�C�{s]�pKQY�PROG��B�������(/softpa�rt/genli�nk?curre�nt=menup�age,153,��!s^�Uo�W63�1,�P le_C�onfig.st�m�Oo�MJUy�SD�T_ISOLC � ���~��OJ�23_DSP_ENB  ^j��`?INC �^ku�l`A   ?� � =���<#��
ka�i:�o ��a�o�o��o$xgOB�PC�c�E�f>q�G_GROUP �1�^k��< �tP�a�	�,?��_��!�� �(��L�^�p�����6yG_IN_OAUTOKt�i`�POSREFXvK�ANJI_MAS�K膯h��RELMON ���|_�yG�`�r��������N���S��WՃ��ʕ�քKCL_L���NUM�`��$K�EYLOGGIN�G�����*�e�PL�ANGUAGE ���f���ENGLISH lt�|�LG�A��Z�R�'��  }��H  �� �'�7  � 
����� /o=f ;���
�(UTg1:\��� � �'�9�P�]�o����� ����ɿ��(O����HQ�N_DISP ��o X��z�?LOCTOLu���Dz�Pga�a��GB?OOK ���-� �Q��-��Ԫ ������/�A�Qݑ�Sc�?�	��ԩ�q�9j�߼�Q��_B�UFF 2�^k' ��%�����>b��G Col�laborativ �%�7��v��� �����������E��<�N�{�r�����DCS ��Y�b�a`� ����E'9���IO 2��� !�@n�@�P�r� ������ $6JZl~�� �����/"/M�ER_ITM[nd ��{/�/�/�/�/�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?��P"�SEV��F�L&TYP[nj/KO]OoO��=�RST���S�CRN_FL 2�[�P����O�O�__+_=_O_�OTP�3�[o:B�NGN�AM�d��f�6�UPS_ACR�@ꏾT�DIGI�XIU�_LOADCpG �%|Z%ANI�MATIO=�RO�P\_yeMAXUA�LRM��Q��2�e
Bb�Q_P�U�P� ��a�B`CA����͜o������ddpPw 2��� �=�	:O�o+Oa D�p����� ��'�9��]�H��� d�v�����ۏƏ��� �5� �Y�<�N���z� ����ן�̟���1� �&�g�R���v����� ���Я	����?�*� c�N�����|������ Ŀֿ��;�&�_�q� TϕπϹϜϮ����� ���7�I�,�m�Xߑ��:hDBGDEF ���e��o��_L?DXDISA�P{[�KMEMO_APޣPE ?|[
 ��z��-�?�Q��c�u���B`FRQ_CFG ��gm��A z�@���|�<��d%�����t���b��k�ԯ*Q�/S� **:\�|�O�a��� |և������������� 2~ߍe[2 L�p��,(0�C ��(9^E �i����� /�/�6/8jISC 31�|YB� ���~/ ���ߔ/��/�/�/B/�T"_MSTR ��M5SCD 1�
��/c?�/�?r? �?�?�?�?�?O�?)O OMO8OqO\O�O�O�O �O�O�O�O_�O7_"_ 4_m_X_�_|_�_�_�_ �_�_o�_3ooWoBo {ofo�o�o�o�o�o�o �oA,Qwb �������� �=�(�a�L���p��� ����ߏʏ��'���K�6�o�?MK���#=�ၟ$MLT�ARM������� �����>��METPU��b����+9NDSP?_ADCOL�����CMNT.� �!�FNJ�N��FS�TLIo�`�0 �#>®���گ�!�_POSCF��Y��PRPMM���STv,�1�#; 4��#�
^�j�^�n�|� Z�|�~���ҿ��ƿ� ���>� �2�t�V�h���όϞ�����!�SI�NG_CHK  }r�$MODA����\+�����DE�V 	��	M�C:N�HSIZE���b���TASK� %��%$12�3456789 ������TRIG ;1�#; l������		�J���YP�ѣ0��EM_�INF 1�6��`)AT&F�V0E0O���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ����H�F���:�n���A�v���Y���������  ���������w*� ��������� +O�8J \���/:'/� �]//�/h/�/�/j �/����5?�Y? �/j?�?B/�?n?�?�? �?O�/�/CO�/?? �O�OP?�O�?�O�O�? _�O?_&_c_u_(O�_ LO^OpO�O�_�Oo)o `_Mo _qo,o�o�o�o|�oG�NITOR���G ?b�   	EXEC1f��r2x3x4x5�x��v7x8x9f�r�Rytrytr yt+ryt7rytCrytOr�yt[rytgrytsrys2��x2�x2�x2�x2��x2�x2�x2�x2��x2�x3�x3�x3�r�R_GRP_�SV 1��� �(j������~�l�w���o�ƥ�_Djb��ԃIO/N_DB$й(�b�_  �ސ�ސY�A���&���  
xF�y�A��`N   4�Z�&��=�-u�d1tՊ����� �P�G_JOG �Բ�ƫ
ˠ2��:��o��=���?�ˠ����*�ܞD�V�ˡm���n�0�'�ˠ+�@�����ѯN�  �ѧ��L_NAME �!�� ��!D�efault P�ersonali�ty (from� FD)Y��RM�K_ENONLY��G�R2�� 1��L�XL�< �O�l dm��� ����ѿ�����+� =�O�a�sυϗϩϻ� ������ߥ��$�6� H�Z�l�~ߐߢߴ����� "����#� 5�G�Y�k�}���� ����������1�C� U�g�y����������� ����	-?Qc u������� );M_q� ������//��<��;/M/_/q/�/ �/�/�/�/�/�/?��_E�a��*/ݟ*?_?��PN?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�Oh?z? �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �O�Oo%o7oIo[omo o�o�o�o�o�o�o�o�!o�ots���(`r}x�d����~ ���w��G{���N8�A��p .�Y� O�a�s�������׏-��Ӑ��
���	`@C�=�O�a� �3�AD�p������[� A�P̙(��q�q��"����tS|���  �tp�pE��C{   &�G�"�k�V�{�����@ů�x�qH�j�p�����p+�� �� ��� @D7�  )�?�/���?Ā1�ā@I��)���˯  ;�	�lA�	 �X  �����y� �,� � �������K��oȩ���]K���K]�K	�.��_�Z�<����@
��J���Կ��T;f�I��Y�,A��{S�ٽ�>  ?�3���Ck�j��#3��?2}H��{�bā��|S-��Ͽ�B����X�\畨� D	�����g  �  �!ֵ�?��	'� � ]��I� �  ��ٕ�:�È~��È=��͙�-�@�߯�ھ����G��-���N<}�+�  'A��|B�I��@�p�Q��V�Cj�Cn�C�Ӏ y�~�J1��|���܀ � �Nſ A 0ݹB }���|��弝���āDz��$���H�3�X��~�i���������А 4�P���ąz��؄ � �p��?��ff������� �&8j�8ĀN\
C>L����=�ݺ(Ā�P�������q��� xi�;e�m���KZ;�=g�;�4�<<�0���/���y�ɐ?fff?��?y&;�@=0M?��YH�|�6 B�ݹ1��/��u� ��	/�-//Q/�</u/�/r/�/J�zF}��/�/�/?�,? ��/_?�/�?n?�?�? �?�?�?O�?%OOIO 4OmOXO�˜O��X�? �OB?_�O_A_S_e_ z_�_&_�_�_�_�_�_o����3dՙG��Cojoo�o����ؘo�o�o�oH��"{�k�}��dD
p,��L�d��`�aUqI���!n,ȴA2=q�@��T@|j@$�?�V�^��z�Ð���=#�
>\)�?��
=�G��}�{=r ��,��C+��B�p���p}B6���C7n����?6`��(���5}G�p��Gj��F�}��G�>.E�V�D�K�����I2`�F�W��E��'E����D��;�����I+aE����G��cE�vmD�����9 ��ď���ӏ���0� �@�f�Q���u����� ҟ������,��P� ;�t�_�������ί�� �ݯ��:�%�^�I� [��������ܿǿ � ��6�!�Z�E�~�i� �ύ��ϱ������� � �D�/�h�S�xߞ߉� �߭�����
���.�� +�d�O��s�����л�����p(�q343�]����9���x!�7��U3~�mU�g�I�5Q����I�Ǔ������Q��������=+(aO�EP�P��A�O���������#\ Gl�}���� ��"//��O�OL/�/p(��/�/�/�/ �/�/�/??C?1?g?�U?w?�?�P2/�? � B�;`p�1CHpz;`�P@BoOO@+O=OOOaOrM�C�?��O�O�O�O�O�S?���C�  @�S$�P�P�aS�4�U
 �ON_`_r_�_ �_�_�_�_�_�_oop&o8o�z(Q ��}���'x#�$MR�_CABLE 2��} ��tT� �f���o�	�o wI�`q�c�ow}� 7]1g��y ������3�Y� �-�c�����u����� 珽�Ϗ��/�U���k�1{B��o����˟������������*A�** qcOM� �~i��^�6 *[��W�k%% 2345?678901~���! {�����{@�{@�15{@{A
���m�not segnt J�ӣW��TESTFE�CSALGR  eg{J�1dC�QڡY
S�� � {D�Xbp�n������� 9�UD1:\ma�intenanc?es.xml����  +Z�D?EFAULTvLqb�GRP 2�b� � �{@}6*[�V{F  �%!1�st clean�ing of c�ont. v�i�lation 56��ڏ�	P����}5+*�}J���������X�%i�mec�hp�cal ch�eck�  �BS��@]�d�}5�π�ߣߵ����(�y�roller;�M�_�����U�g�y�����(�Basic �quarterl!y���$��,D��`#�5�G�Y� �M2���{@"8��N�N���}5�����b��t�C��O��s���������&(�Overhau��6|�' x{@18}5�ew���{@$V����wI T)/;/M/_/q/��/ ��/�/�/??%? 7?�/[?�/�/�/�?�? �?�?�?:?�?!Op?O �?iO{O�O�O�O O�O �O6O_ZO/_A_S_e_ w_�O�_�O�O�_ _�_ oo+o=o�_ao�_�_ �o�_�o�o�o�oRo 'vo�o]�o��� ���<N#�r G�Y�k�}������� ��8���1�C�U� ��y�ȏڏ쏢�ӟ� ��	��j�?������� ��������ϯ���� T���x�M�_�q����� 䯹�˿��>��%� 7�I�[Ϫ��ο࿵� ��������!�p�E� �Ϧ�{��ϟ߱����� ��6��Z�l�A��e� w�������� �2� �V�+�=�O�a�s��� ����������� '9��]������� �����N#r ��k}��� j�8�\1/C/U/ g/y/��/�/��/"/ �/	??-???�/c?�/ �/�?�/�?�?�?�?O T?)Ox?�?_O�?�O�O�O�O�O@JnB	 X`�O__(_lIB IO W_UOWE__�_�_e_w_ �_�_o�_�_7oIo[o o+o�o�o�oso�o�o �o�o�oEWi'�9������|� �wA?�  @nA 5_0�B�T��nF�������lH�*ŏ** F�@ �q�vp�����!���E�W�i�{��� zOFFߏ��ϟ�󟵟 �)�;�M�������� �����������Y� k�}��m����S��� ǿٿ�1�C���3�E� W�i�+ύϟϱ������WDnA�$MR_HIST 2��u}�� 
 \B�$ 2345678901�#��Ͽ��9Ozߌ�C�u� O�����߯���.�@� R�	��i���c��� �������*���N�`� ���;�����q����� ��8��\n%��nD��SKCFM�AP  �u��q���n@���ONREL � nD�����E�XCFENB�
8��FNC�JOGOVLIM��d�^�KEY��aj_PA�N�|x�RUN�Qa	�SFSPDTYP5 ��SIGN�T1�MOTS�_�CE_GRP 1��u���@r� _/nCL/�/�s/�/k/ �/�/�/?�/?D?�/ h??a?�?U?�?�?�? �?�?O.OORO	O\O �OoO�OcO�O�O�O_��K�QZ_EDI�T���TCOM_CFG 1͹ae_w_�_ 
FQ�SI �6+����_�_��_o����O@oXT_A�RC_�@T�_MN_MODE���=Z_SPL�co#UAP_CP�L�o$NOCHE�CK ?� � �o/ ASew����������NO_?WAIT_L�;W6& NTNQϹ�Ez�Y�_ERR0!2й	����'���Ə؏��_�/�~`�O��ю�|���*/oW��<���?���v�\�� I���P�ARAM��ҹ���G�������(� = V�E�W�_� 9�����o���ɯۯ��0������C�U���y��cUM_RSPACE�i��Q������$ODRDS�P�c� OFFS?ET_CAR1P�o��DIS���S_�A~`ARK�<YO�PEN_FILE����Q<VαPTION_IOr�s��M_PRG %���%$*�Ͼ�O�WmO;��6'��Ar����:!5�����	�j�	�	 ���	���$d�ϰRG�_DSBL  Ğ� r�v��RI_ENTTO� ��C�� �A �U^�`IM_D{�����ϰVӰLCT ��c�8RҼ��d<����_PEX�`�n�RAT�g d ����UP ���b�; �{��s�|����$PAL]���c���_POS_CCH<�&���Ő2/#��L�XL���l�j�D� V�h�z����������� ����
.@Rd v����22�� ��#5GYk}������ �//%/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_k� ��_�_oo+o=oOo�aoso�o�o�o��E�a:Ҭ��o�����o	:�P�o3EW i{������ ���/�A�"w� ��������я���� �+�=�O�a�s���T� f���͟ߟ���'� 9�K�]�o���������dɯۮ��;����j�dg�8�J�/� m�{���e�������进�
�׷���	� �9�?�]������4��:�ֵ	`���x��	���:�o���'�9�K�]�f�A�C  t�и_�_��e"�x����ӿ�  �����#���C{  ο��ʿ���#� I�4�m_��Z���OU��/��/�H'����� � ����� @D�  &��?�����?���ᆟ�C4����s� � ;�	l��	 ��X � /�4�%� ��, � �xE�J��Hʪ�U�����H���Hw�zH�P����������B��  ������������>  �3���C�����c���������B���������R��f� ek�������T� D�������g  �  ���]����	'�� � 	I�� �  �<�Ռ�=���-?��@U[�����[������N<%��  '����C C C�� ��*�/�a�`��$�z�� Nq� A 0��B%Ѕ%$ё%0d�l�%��DzV��/�/�/�/?*?��݀A2��I2�� 4PI"Z5���z��^�|���l ?�ff���?�?�/? ���?�;��8���?J>LO~ ����(��6EP?HZ9<�`3�7�C1 x���;e�m�B�KZ�;�=g;�4�<<�m��O�?������%Bq�?ff�f?l?&�@��@�=0�E?�� U�Y$��A�����=_ ��\_�G!��?�_|_�_ �_�_�_�_�_!o3oo Woio@o�oxo�o(_J_ L_�o�o/S> wbt����� ����H����o ���o��z������� �O&�8�ҏk�V���z���ş��"�ߔ}���C�����:�%�?Ƀ�D�K���o���E�� %�~�D���د�^��^�]��@�I�͞,ȴA�2=q@��T@�|j@$�?��VT��z������=#�
>�\)?��
=��GH���{�=@�,��C+��Bp��[��B6��C7n����?���(��5�G�p�Gj���F�}�G�>.�E�VD�K������I2`��F�W�E��'�E���D��;������I+a�E�G��c�E�vmD��� ��:��7�p�[ϔ�� �ϣ����������6� !�Z�E�~�iߢߍߟ� �������� ��D�/� T�z�e�������� ��
����@�+�d�O� ��s����������� ��*N9r]o ������� $J5nY�}� ����/�4//�X/C/|/g/�/�/m�(�m�34�]�/mA����%�%�/�/U3~��m??�"�5Q8-???�"��Y?k?Q����=�9�?@�?�?�?O�<n�P�B	P?N^�[�hO�/tO�O�O�O�I���� �O�O_�O_>_)_b_ M_�_q_�_�_�_�_�F`P�R��_.oh�1o ;oqo_o�o�o�o�o�o��o�o#Is02<�_t  B�琾���qCH��z�s0@ ������t�cH�Z�l�~���fs3?���=@ @s3�5ts0s08�8��[ts5
 ���� ��0�B�T�f�x����������ҟ�c�ԁ ���);�'x#��$PARAM_M�ENU ?�5��  �DEFPUL�SE�	WAI�TTMOUTH��RCV[� S�HELL_WRK�.$CUR_ST�YLF���OP9T�q��PTB�����C��R_DECSNS�0E�\���!�J� E�W�i���������ڿ�տ���"��SSR�EL_ID  �5YA�1�USE_PROG %,�q%σ�2�CCR_��C�YA4���_HOSoT !,�!���ϐ�TP@���û������0ߏ�_TIM�E]�Cƫ��GD�EBUGA�,�2�G�INP_FLMS�KY߈�TR�߈�P+GA�� x�7����CH�߇�TYPE
)�5���M�v� q���������� ��%�N�I�[�m��� ��������������& !3Eni{��������WOR�D ?	,�
 �	RS���CP�NS�E��:JO�ɡ�BTE�D�COL�E����LV_� �0�s0ȫ��dm�TRACEC�TL 1ׅ5�6� =@ �*=@7@��D/T Q؅5 ��D � i�� ' 	+$
�+$+$+$�0-"�+$+$C�-"+$*+$+$+$+!/C�/WA-"��-"Ѐ�-"��-"Ȁ-"Ā-" +$*/</N/`/r/�/�/ �/�/�/�/ ??$?6? H?Z?l?~?�?�?�?�? �?�?�?O O2ODOVO hOzO�O�O�O�O�O�O �O
__._@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�o �o�o�o�o�o&�8J\n��� #!�%k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w���g��������� ���!�3�E�W�i�{� �������������� /ASew�� �����+ =Oas���� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgOyO�O �O�O�O�O���O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ m������ ��!�3�E�W�i�{� ������ÏՏ���� �/�A�S�e�w����� ����џ�����+� =�O�a�s����������ͯ߯�����$�PGTRACEL�EN  �  �����3�_UP �/���b�j�N��c�3�_CFG7 �b�L��
c����������|E���  ����w�DEFSPD �ۂ��E���3�H_CONFI�G �b�J� U��d)��B� �,�PôƱH����3�INz�T�RL ނ���8lõ]�PE����b���(���3�WLID{����	�ɿLLB 1��� �I�B8�B94Ӵ� I�!���LŶ� << �?�K�j�K� b߄߲ߘߺ����� � ���8�f�L�n����4��������M����<�/�A�r���GRoP 1������@A!���4I���A �Cu��C�OCj+VFx����-�Ʊ0����(�(����q�C���´B$BE lL6H�l���&�B34�����`�j 4MJ�n� �,����%//  DzJ#S/��:/ {/*/�/�/�/�/�/�/ �/??A?,?>?w?b?Л?�?�?�:)�1
�V7.10bet�a1��+�@��*�@�) @��+A )�?���
?fff>�����1B33A�ж�0
CB(���A���AK�� �9AD	AVOhOzO�O��O��p���8�@�@>K��@A���?��ff?�@�������Mb�������?��? �,_>_(_b_L_�_�1)�l��u)A�Zb� �_��_o���1EE�A6�S BڰB�:o,eSBHbc�T���MdI���T��Q�
�Tx�dxo�o o�o�o�o l���2��- ?s)WM_	t����KNOW_M  �������SV ��?�Y�i/� � ��_D�/�A�z�������M���� ��B	��6� I��^��Z���Oo
�b�T�@ڱ��1ڰ$� �2����MR��鯍T�_^+������~�OADBA�NFWD���ST^��1 1�b��p�4EOAT �w/o part��B�����=LQ� 0�B���f�x������� �ү�)���,�>� P�b���������ܿR���2򜻁4ڿ  G�</���3�+�=�O��4l�~ϐ����5���������A6�$�6�H��7e�w߉ߛ��8�����߬���MAҐ�����OVLD  ��ޏz��PARNUM  ��p��#���SCH]� k�
�������UPD���^�>�_CMP_��`�����p'ޕv�ER�_CHK����`ޑǂ������RSq��՟�q_MOҟ��_���
�_RES_G
���
ROʽ_d ������� 7*[N`3�@P�5k��� �7����/7� /</A/7d�\/{/�/ 7�Л/�/�/7
��/x�/�/7V 1��f|ې��@`h���THR_INRq��bፂޕdm6MASmSz? Z�7MNy?��3MON_QUEUE ���ޖ V�@ 
�N{�U��qN�6�8�3ENDAIEXE*OE@��BE)@O�3OPT�IOG(�0PROGRAM %�:�%�08?���2TA�SK_I_�qNOCFG ��?���O^PDATA���[`a��2ƅu_�_ �_�_�_h_�_�_oo�)o�_Mo_oqo�o6_IWNFO���S]��4 ?o�o�o $6H Zl~����� ��� �2�D��g�d��S\ nQ��DIT �_����>TWERFLKH`3��CRGADJ M�A���? `��1��1
P�a�_�?���z��NcQ<@����f% �`r�وn!�MQ2�/�V�b	H�0lA7_2�<�>�����t]$�*�/� **:�� ��d���6�1����;���a�C2[�)��� 9�K�y�o��������� �ۯ�g��#�Q�G� Y�ӿ}�������ſ?� ���)��1ϫ�U�g� �ϋϝ��������� 	߃�-�?�m�c�u��� �߫�������[��� E�;�M���q���� ��3�������%��� I�[���������� ������w!3aW i������O �9/A�ew���X6	"_F/ۀ 4/m/X$㙏/�[/�/�W/�/�/���*S�YSTEM�V9.40107 2�7/23/202?1 A%݀
7���#�PREF_�TLA( $GR�ID@ES  �$BARcB]2SoTYLE]1 ?0�OTOENTJ0�  $P_7NAMs0!�0{2�]1z1XY(�J1 �� $LIST�_PORT]2�3E�NB�8SRV�0)��4�6DIRECTS_1�2�42�93�9U4�95�96�97�9�8�1  �PF_�HRK0  Q0VA�LUEv�S0OU�Pv�$AXIS�zA��YA�4� !$ENABr0� �1G�3�%$CUR��wERcAN�C�Bn0AR�0�YPoA$TOTAL_TI�Ar@�C�PWRpBIC1�DR�EGEN�JRpBE3XE\A�A$]C�A�^1REe0�EMON�TR_R)Q�2�A_�Sx@WWP:SV_L�IM�0tV@�1EG�RE�CG0?PHzBO�VERU0�TV_H�d0DAYSV�QS�_Y�A$MAX�SIZ9SSUMM�AR�P2 $�CONFIG_S�ET�CUP�2{AL�A�0RUQ=QC_�o6$CMPR�4� cDEV�@�P/bI��@Z c�S]1�BE�NHANCE�A | 
�E*a�@TTN�QINT�0QM(�|^1��_MASKj3PD_OVRD�3�GE2IX�0JPAX�yPZ5OVCyQ�TB�UqR�CF5 4 �S?e71[o6�PS�LG�P�A \ �$PS_�V=pMO�P^1�AS�0ra3aU<q�fTv�SDbtAU�A-p80P�A (0Q�Ar�JvOPCrFI�L_McS�qVELL:S�0TQLP�3N�0�.PCPSUL�P _ 	$V�{C��P_�po@�M'�V�1&�V14�2C�2�4�3C�34�4C�44��A�0 ��@��ܿ0��MINщVI#B1+0��2�*1T����3��3��4��4���@�L��@@���@̇Ʌ݅ɅPLUS_TORQnAp؅����+pSAVba�	d $MC_FOLDER`	$SLđÑse��@M�pIsc��LO}A�`  $��2cΐKEEP_H�NADDّ!�R�#�CCOMi0`;�{1ڒ=p<�OP ��b�ؑ_0<�xg<�REMS�;��A�2x�ԏ���U�4e;�HP�WD  �S�BM�a�0COLLCABLt�@>p�AE�a��@ITSa��r�$NO�FCAL(c�CDONrb�qÒܚa�0
 ,Q0FL�ANGoA$SY�NҐI�M�0Cb�~�@UP_DLY�1=C�DELA{��A�k2YPAD�Q$TABTP_R���QSKIP:�g Ĵ0�PORk������P_�Pʰι �@J��b�}Q���Q�� @��@��+@��8@���E@��R@��9�a�R=A�3 X�P�B��gMBa�NFLIyC�3��REQU�0<�cqwNO_H��r��,`�_SWITC�H�2RA_PAR�AMG�q ��_0mhUSE_WJ�[r
��SscNGRL�T{�O�q$WA�RNWpYp(c�STb�@J1���rAP#`�WEIGH�3J43CH�01�OR�11���bOO�@;RATI�O/�J�@D�0�bS�A��&e�ӓ�OBO��Du1W@J2���1��bEXD_RTQTD_IT�C��@0�����a��@RDC|�A=� � �`d�`��R݀��TH?Q�����RGEAPRIO��8�W�G `Y��?PER���SPC����UM_�бs2�TH2N�a���� �1 (�ED�{1�2  D �liX�LVL2_P���Sgq�QP�L10_CA�q�'���a  h :q�0��j�0(S��q J�H��М�Ձ�b 񩓁�@�Bb�zApW@��`�� P��DESIG"���1
�1�����10���_DS�q���E�FPOS11�1 l�B�ZrH��C��SATq����pU��EIND�`�1= �=0���HOME(g0�2/�ASew�3 ������L04);M_q�5���P����6/�#/5/G/Y/k/��7�/�/�/�/�/�/
�'8??/?A?�S?e?��Sߠ1  �QP����я�ЎB T0��D�FCIO�q=I�I�0bO�_OP�IEaC�B��POW=EӁ @H�r�/��D C�ޘB$DSB?pGNA���v�C�����S232#E  ��9��5H�3`ICE���SPE���Q��I9T�Q qOPB��RoFLOW�PTR1�4�Q��U�SCUPi��a�UXT�a�Q�`EORFACT��U%P���SCHca! t�Ր_	P`^��$FREEFROM�PPsAq�(�A`�ۑUPD�)��PT�0&eEXذ�X�S!��FA�p2b| �@yPdPca"� �
�5�AL�q�9P��EX`PIQb�P1PY8e�B_�r��4aQSf#WR�a�?�9DP�wf�P��6FRIEND<:�p$UF��t޴`TOOL�fMY�HՐ�bLENGT_H_VTE�dI�q��c��$ �`�hU�FINV_ y��ARGI�q6�IT�I��gX���g=vG2=gG1Ga^P��WrhwPRE_�b���D���a�����S�cEQ�ӀC��b�q�v �8��lS~Q# @.@P� Q꒬zWhjU�jU����B��P�T$�X �M�PCTQcH��YhP�/U)d�S%G��WI`m�҂�	D��a@Kq���ʰ�ؒ����$�v C2#�qa wi1�h�r`2uk2�3uk3 �j։-��i�I��60`��0`!�$V�
rV>uV!�
q��q�rP%7�kV��ߡO��v�CR�����b�Z���E�e��	s���5$AG���PR����p�S!�PR��"�R&A�& ����+�ˀ$�В�ˀ%π�P�p^P�β
@�S�A' �ؠ�R��7A\�/@U�NN�@AX%Q�pA�`L�ar´�THI�C��G���@�^PF�ERENZ���IF'_CHkc��Iug���6��G1���0$�t�
p<�_JFE�sPRL�_��RVW��A~Q(  $�X�;Q  ^�VAL"E� ��j�:�)�Bn��  2( �S�,�0*
  �$�_���a�����γqT�Ь�γDSP�&��LILSpE
��A0��šȳ��AX��UV=K�P_MIR�!�2�pMD�B�AP2� ��E/`b�AԶ�SYS�8�R��PGw�BRYK�r�VNC��I�1  ��vc��в���AD;Aγ;�BSO�Cٶ3@N��DUM�MY166�bSV�\�DEfASFSP�D_OVR��^�f��LD��OR��0N���F�֫�OV�SFTڥ�W��Fp�Q%Ås���a�lCCHDLY�R�ECOV��pT�W��M�����������r
�_��\� @���,pVEz@�1OFS2,pC���cWD8���`4����2[���TR5Q�	A��E_FDO>[�MB_CMKAF�B BL��@�hⰑ+�VlQ�R�PY�ƳP�Gi�|�AMz�\��P�������_M��NRMŰ9B��T$(���Q>�3T$HBK�Qg��IOue�YA��PPA�?�$�O�7����YB��DVC_DB/s��h��B����2�"��1�����3����/ATIO1�]Q,���Uzc�8FCAB 
�tb�s=����0���Q�T�_RPg�SUBCPU���Si��@R� ��P�Sp���B�?$HW_C<Pȭ����Akq���$/UNIT��� � ATTRIj����CYCLcNEC�A��L�FLTR_2_FI��H��F��QLP�����_S�CT�sF_�F_�8�
FS�A��CHA�a y��CRxRSD�зB��գ찡Y@_T��PROX��@�9PEM�0_��r��Tfw� f̀��DI`i�RAOILAC���rM��#LO���c��7�b␰�������PR��S��qπW!Ct��@	���FUNC���RIN�ps�o` w$8Q3RA� �b �#8
@	��#WAR5���#BL�q�'�$A�+��(�(DA���!8�#�%LD�PЅ�33�2�!�33TI�S5�ɱ��$�PRIA��QRAFD P0��~3�Є5󀘂��MsOI� C�DF_�`؇ӸQ;PLM��FA���HRDYPdORG80H��ao`0�5MULSE�`j�S*���J�J6�K��F�FAN_ALMsLV5SRAWRNYEHARD���V`�p��P� 2QAQƱ��_,��g�AUmPRkOR?TO_SBRv�E���J� v�!�CMPINF����D)1n�CREGvfNV�P�!c��DA�`R�FL��$M0��RGd�ࠠ`HgUCM�uN��Y�#NONI� �NE�PYBjRs&���8I�๱+ ���a�$Aa$Z$q�������,$ ��o�EG�γ��QAR�����23#e� �|�AXE�ROB.�RED�W�a��_]m��SY��8a��:fS�gWRI��f� STR䵼@��*�%E���d8�A"�B�`���f9'#���OTOQ����ARY�r!!������FI��,�$LI�NK�1��'qc�_�c����3O��`Oq�XYZwBYz�jsO�FF��&rNrBxpB�l"�t���p �sFI� �ww��4��l"��_J���@(�3s���@�d�j3p����TB�qB5�CL� k�DU���32�.7"TURT@XZ3n��q�BX�`���FL�m���`��pu�i3z9�
� 1+��%K
�Mg�\�54%S8�S%�ORQ�� �##���␂�1��0��<�j��#QQ�OVEX���M,0��Sr��S r��Rq��@o�p��  o�B�q ,�0��Y�9� ����0�j�Y�v����S������ER��!	B8"E��|�D#9�A����u�%�w11AX�ӆ�1� � (r�����A��ƀ�� 쀞�����3 ���`���`��1fp���0���0 ���0���0˩�0۩�0 ��0���0��0�8��,�� �2~�DEBU}$x!�C���JrAB'�8�R�V�| 
©�� /�m;�e�;�Ɓ;�� ;���;�3!;��a;��a��4:��2ϒ�sLAB��r�y ��GROh� �}L��B_�  ��d1ӽp�@����8ձA �ANDڀ8 @.���Su1��A]� �စQ�`q�1��� RpNqTd@�ӣ�VEL� ͔��!���r�0ҭs#NA��phbC�T��`s3#,��b  �S�ERVE���P- q$�p� ��!)�SPOJ�� _�T9P�!�P��1�P.�  $M�TREQ��
L�hbV�/Z�Ƅ22.k�b0 _ �0 lT�AERR�ra�I���͔N��TOQ͔ʐL<`P���b���G+�%<q�"�V`0 1 �,'�o��/ёRA~� 20 d0��f��b� 2�P$f���0���P�M�OC1x�3 � ��COUNT��aZ�Z�SFZN�_CFGU�4 4� %V�T"z���<���� �n��^�S5 �,�M��+B��pɓo��F!Aq0ؕ6XX`- 	���Ga,�� Xa9PzB�PHELAP��6 5�pB�_BAS"RSR$V` RcS<L1� �1�� 2�
3�
4��
5�
6�
7�
8��RO�� �-pQp3NL�Q@�AB8�
 n� ACK�IN^�T_UUU�@	@�AL�_PUX�~Be2OU:�P� %Xy��@�`�y�TPFWD_KcAR��-Q��RE7���0P#p1� QUE�$Yf�Y�I���~@�AI U@�yOp���VOq�SEM�q?&E��0AnSTY[SO* P�DIg�@��!x��1_TM9SMANsRQ�&OpENDN��$KEYSWI�TCH��z!$H}EI�BEATM�PE(`LE��� �J�(U�F.$�S$�DO_HOM�0OlzAOEF9�PR�qP��ja�`UUC
0O�1<���OV_M��pE�pOCM;�'E���RzHK�Q7 �DLq&W��U��"M�`�K�<�FORC.*SWARձD�x�OM` 8 @����s�@U�cP`1(FgPD3F4�А��Sc�O�L�29<�%XUNLO���mZDED�A  �P+0��: <NP�1y�}�MSUPGN���ACALC_PLkAN�C1�pAY��a�zB��; � 	�@9�PA�$�MQ{A@ϵ�·`���%Md0����r�F�Td��RSC��M�P�ѱ� �<Q���p�OTYWZZWZE!U AR㐡PTaՈR��P�V�2NPX_A�S��< 0� AD�D����$SIZ�eA$VA���M_ULTIP<�S�@A�1= � �$��P>2�p6bS���aC��"fFRI	Fa�^�S�IB4`{NF�$ODBU�``��#efcai7�CM�!$�ձ������Ƃ�k� !�> � ��P��TE��
��$�SGL�aT5r��&���c���`�`STMyT��sPSEG8"� qBWY��dSHO�Wub�BAN�@TP�p���,��7��l�V+�_G��? �$PC��_�+�֏�FB�1P�xSPb Af�u�VD�p~��@� ���A00���q@�w@��w)@�w3@�w5�y6��y7�y8�y9�yA �y�@�w @�w���v�@B�wF�x+����y1�y��`���1$�11�1�>�1K�1X�1e�1�r�1�1��1��1P��:�x��y2�y2
�U2�2$�21�2>�U2K�2X�2e�2r�U2�2��2��2��U3�y3�y3�y3
�3�3$�31��H��K�3X�3e�3r�3��3��3��3��4��y4�y4�y4
�4��4$�41�4>�4�K�4X�4e�4r�4��4��4��4��5��y5�y5�y5
�5��5$�51�5>�5�K�5X�5e�5r�5��5��5��5��6��y6�y6�y6
�6��64�6A�6>�6�K�6h�6e�6r�6��6��6��6��7��y7�y7�y7
�7��74�7A�7>�7�K�7h�7e�7r�7*�7��7��7��H�VP_UPD�qAs Z��C 
:@�V\b�qB x �$TOR��`  �7SO�� l ��Q_w�RE�r��'��`��S��C1����_�U;`��wBYSLO>�C � �Udb ��Qd�W$05�0�RVALU��q���zR�F
�ID_L�#�z�HIu�I�2$F�ILE_����q$?3���SAV�q�D h����E_B�LCK���q��D_CPU���P���P�u������� �R �E � PW��`.I`XLAq�SR��]ngRUN�@G�\�g�  ��\�gH�s�� g�1T2�_L}I�2F  '�G_O:"�P_�EDI2�@T2SPD�G�PIDxq`��DCSy �Gi�H � 
�$JPCw�s� S�PCOC^$M�DLQ$u0~T�CP�UF� S�COB� � N�;�r�pI�0M�\��Oz�aT�ABUI_<�pJ<�B< HD"R�I$2#A�S�`LLB_AVAI2���1$�qK �$� SEL� NE\s� RG_� N�`ؔAq2#SC�0LS �o!B@TB��q� _M�@�pM 1\��PFo1L_���&)M�b-@G�pUy2]t]6ZrPS_XbP�`� �P,5Ew"�TB;C2�EN ��`�@l�@�B$�FT@pqag4"PZ�TDC�e�� �0�P;c�5{7THDX`�1�4��7R�{$�PERVEn3��4{3�4�aF2_AC��0 OX -$A�@n3D{3@� rPI`aPLOW�'F1A��2HG*P���`3C\`ERTIA�5T��pI��@�KDE|�EXaLACEM��CCcC��V2�P�F8�E�G�ATCV�L�A�GTRQ�LUZ�r �C�q:U�C�qJQ��DQZ�Ja��p�E�Q
�EA2�9p*!@l�C�0JK�VVK|q �Q�1�Q�a�PJpq�Q��SJJ�SJJ�SAAL�S�P�S�P�V�a2�R5�3)PN1\)`��K�@uD�!_qq`����G1CF�"P =`��GROU`��a�ZB�qN^0CpS�`R�EQUIR�2>�E�BU3�1�� �2O�a�0�fG1S�GL5Q�  AP�PRPCw ��
$:� N�hCLO-yaS�5y�E0 BC� ]AR �d0M�0p�@P�2Wt_MG��apC�p��kx�0lw�BRKjyNOLD�jvSHORTMO���z�}[uJ�!3CP �T�@�S�@�S�@c�@Pc�@#1�r7�u8�1���1M4S� ��b(Bn1G��1U�PATHQ�j�`�j�-Hhf�Gp�`R��NT� aA%�w�b`qIN B�UCt@[A��C?PU%MɈYJ@��iPЁ�~��1늣0��P�P�AYLOA�wJ2�Lf�R_A� *�L�Y 6�2�&�B�kuR_?F2LSHR�4o�LO7���p�̓~�̓ACR��������r�2HS�uB$Hkr^ޒFLEX�c;BJK6T P�b\?�n?�?�?Z@@qJ EU :OF�@p����"O�1�@+O=OOLF1��ե�^OpO�O�O�O�O�E�O�O�O�O 
__._@_R_��TW ��T���s_�_�_���ZTa��X��gQ�U \�D��U�ŗ��_�_�_ �P�Ue�Ueo1oCo�Ui�BJhdV ��W0uo�o�oZ�g�AT��a^PELp��"��j�hJ�`U�`JE�p'CTRw"��N������gHAND_VB����_�M4W� hQ@kv�4M�SW��� ZG0EvX� $$MT�Xy���q���q�쳰��r��A@��#�[v����d}Au|C��zA�{A�{��v{T �zD�{D�{P��Go m�ST�wu�yu�N�xDY� �`kv ����4�@f���f���@%��WDį����uP�u��u�
���%�.��9[�M4Y w�\��O� *�s)qA'SYM��P`�`���XR`������_SH \b��؄�}�H�����*�J1��pC�c�Yb��_VI+���)s�V_UNI�3���n�J�U� �������&��^P@���pß՟f%��딴�D2E�pCHh Z ��dO�[TO��PPD�V�3(�$�5��R��P�q�� Xq� �$�!� _u�����0�%�!����PROoG_NA�$Tj�$LAST�qR�C�AN���3� XYZ_SP���$X7�� ��l6S� 05q1EN�p14CUR�(z��`oHR_T�b[A�D�1y3N��pS�O�48X��0�\ ����I�A�$�� A���C�����r��0 �] � Y�M�EX���)Bc"�T�0PTFe�q�QAU`�Yd�(VHqAeIT�GZa $DU�MMY1��$P�S_ �RF   tq��F�FLAj`�YPR��BYC$GLB_T���5�EQ@��&@LIFh^1�E��f�@OW+@O�.UVOL�a� 0Q_2Ɂ�D2.��@�p`P�6R�00S�@TC�?$BAUD��S�ST6�B��@AR�ITYpSD_WA��TAIUYC��r�O�Uv��Q�YTLAcNS�@�[��SZ\C'�BUF_�RL���x�X�0�YCHK_0�CESɡ��JO�G@E�AQ!4hRUBYT:�KiH�Kd�r n�nf`�Q��!��fH�q�>���1_ X
����aSTY���S{BRU M21_� ��T$SV_ER�R�e�cCL�@�bA�q�O�"�0GL�E�Wh` 4 $�[A$�Q$�Q�$W3sy��!U�#0R�ɂe�qUua �b�"4$GI�{}$q `&@8qLphb L$pnv�}$FEvvN�EARR�?2$F�yO�TG1/� �uJ0R�� cw�$JOINT��z�tMSEThd  kwE�ur����S���1�q��he��  ��UX�?����LOCK_FOx��`��0BGLV��GLg�TE:0XM��&�EMP�pz�8���BR�$UP�rF{ 2a��Ls��b|�h\�W���`�aCEo�|sҀ $KAR��}M�3TPDRAp��qVEC�� ��pkIU��c��HEY�OTOOLɣ%�VȤ;RE�IS3H�E��6/��!CH�� d&�1ONWE�D3Wc;��I�"6P@$RAI�L_BOXE{!���ROB0��?�~�aHOWWARp!x���@m�ROLM�B Ǖd�j�ؒ��6P�;�O_F��!��HTML5x1K3��Pࠥ�� r_�hf�~�#��� W�hg�r����q��v�Phh 	t�Э�`NA�Ҵ�R�V��PO[�1IS0��NP�;���_����|2��!ORDEDW��� Q��pXT��%1)��3��O@ i 7D �@OB��� W� �C�@���wSYS�ADR���0Q@� �� j 9,b�V$A^�!5�\�=5%APVWV�A,Ak � �0r�5PR�"�$EDI1��VS�HWR������I1S�p�Q`ND;@wc<س�cHEAD+` 4�;��KE�Q�@sCPi0�JMP��L�5C�TRAC�E�4l��Q�Ij��S��C%�NE.�<���TICK/���M�1�02�HN�am @��O��7�C7�P�6���@ST�Y�"k�LO�AS� (0ě�ns�
0 6S%$��"4=��SW�!$�{ @A�Ear�EP� �6SQU��RLO�B�TER�CU@Z� S�o up�`�׭ s�������OV@ICU IZ�D"1�E�A%a�B����A�PP�R��_DO�?2[�X�PS�1�3AXI�Q����3E�� T���P�REQ_�,�ET-�*P33J���F���A���D9BX�0 �"�SRdplmз����s��
����VJ1��h���A ���q��@��A8��� I���� ��D+��PH?���C��,�C=��%7ID�TSS}C�@ q hu�cDS�����@SP� &AT*�J2�ь��[BADDR)c�$�P� IF3��_'2CH+�/`O����m �TU�`I�� r�rCU�PN�1V<�I�2sM�t�.T�C�
��
;�Vj�����0t \�`��� �����@0�C^���Q��
���b��TX_SCREE�u�0_P��INAs|pL�"4-�.�.Pv TA��`�B,��a���`��+��ҕ��RRB`��q+���D��UE�7�w ���!a�@S�q,�RSM����U`۠W��6!�0S_Fs�#&��!&)A'��.�CxL��� 2vGUE��x�2�bf&~1MTN_FLj���1�`���q^�BB�L_o�W�@�0y �����"O@q�"L�E^�#����$RI�GH�TRD�dTC'KGR�@5Tܠ
7>1WIDTHBSͰ�B���A+bZ�UI���EY���z d�$p
�Ɛ��6P��B�ACK���B~5q�4@FOɡ�7LAB���?(4@I-�P�$UR���0�pW0:@�H� { 8 $�0T_�l�2;@R�PR�GSu��A�pR�1Oe�`|��w��PU� /CR`�ґL�UM/C�N ERVȊ�pW0P�p^4} 7� b�GE�2�q�Y���LP�EW�ET���)�G��H��HTY��I5�K6�K7�K MP�@RҚӸ��pDU�1Y�=`A |�V1USRt~ �<�`�0Urr�rrF�O� rrPRIj�mxy��рPTRIP��m�UNDO6�ipЙP�չ�������+�` q��2KP$aG ��aT���m�ROSr���VR1��S+��!��"4s;~b��fA��U�A�!�o.o<#�B��N�SOFF��� � %DcO�`���u��dZ�d�u�GU&�P�a��r�c���gk1SUB��� ��E_EXeE6�V���SWO�� �c`�W�WQA��KPq��J V_DB-sEp;�KP	T`�䅖��q��;#sORo�uuRAUD "vtT�yD�[q_��7��� |��D�OW�N��s$SRC���0�D���u��M�PFI����-�ESP�є�d=�^CޱZG�K�C�u���� `�e`rs��2�COMP�$���P_�p`x�o�k�v�7rCT3�q)�qK���DCS�ŐPL��4 C3OM\PZ�Q�{�@xҏ��}�HcCq�a���o�VT�Qg`
�bY�Zޱr`K�F�� �ѷSB$�>�r���_�M*�e��gDIC_�AY�.��PEE0T�1��#VRq��$������0C�� <������W���~ Gg5�vsA0�4������ �~�SHADOW��Q
�_UNSCA̤��OW���DG�DE_LEGAC�i���VC��C>\c�� ��%������R�w�0�w��@Cr@w�DRIV��8��C�!��h��� ܂ MY_UBY+T���c��1� d)��0�̱_ ����&�L��BM�!$nZ�DEYI�EX� ,��o�MU&�X=�l�� US*��{P_R@bobpPc��paG_�PACINj��RG�q����zc��9c��K#o�RE�2ba�bq\���� � � 
a�G��P/���P]�	R`� �f0(@�L1��b	n���RE=�SMW��_A���`k���OAQ-1Ao�s¨��E��U��ϒ ��P]�HK�%@���EП�o����EA�N��prpr�`]�MwRCV�!� �z@GORG�Б�#	�8�c���REF�'$� ���a�k@[�I�PPڀZ��Z�)�|�ֱ�_ �p�ʲ�����SP���ˣڅ�]��$� ���?�Q\QХ�O�U�؛� ����2�� Mq�jP�-��F� N �UL_ �.�CO��i��\�Y�NT )��䩂��A��8Q��e�L)���0���A��8Q�VIAv�� �pHDw v0�$JOP�"��$Z_UP���Z_LOW5��d��1x�"���$EPY� �S�Y%��@G\FG �
�q��� m5-PA81 -oCACHf�LONр����]���C1���CJ��I_F����T�������$HOrps��Á���O� 3��L2���q}A��VPx�� 0�_SIZf��Zd��5�7q3�MP�
FAI��G�V���AD�	o�McRE���GP �R��py�ASYNB;UF�RTD-9��3OLE_2D�_tcUW9c����U�K���Q��ECCU�VEMհ�����VIRC�M5�9_~�j�P�P��AGIR_�XYZE -#_�W/�(L�$dk1�Tb�L�IM��L�C0��GRABqBa<�{�LER��9CN�{�F_D(���.V50�()��%B ԛ��O`�2LAqS902ћ�_GE��� ����q�O�%�T���b�/�9R�I�4����BG_L3EV�1��PK���,�Q�GI� N�0t�%��0����k��P���S� ��N�4��L
q����σcAO�*SbD�QDEY��q�8��8B�W�
a��p
�b�WP�:ڄ0T8S*��Q�DtQ�ParPuTĂUfq� $&qIT�RyP�1��ΖbVSFd��� a �Po���_�UR�ƛSM�U��R�xAcDJ]@���ZD�Fg� DHV�AL?�x� t U�PERI�"$MSG_QM$���7r��gp���RzG�Q^�c��X�VR�T��"�PT_����2
�ZABCBbu�RڃC�
�!��AACTVSg� � � $�U<3 
SCTIV�1G�IO���SB��ITlU���DV�
���Y0���q `P	Sݑ�r ��rGސaGLST��G��M�\f_S����R��CH�r� L mq�c�U���j�D���� GNAET`��G��_FUN?�G �!7ZIP�t�TRQ��$LˢA�u1ZMPCFbu��Bp�R��qڡLNK��
�q ct� �$@��tCMCM��Cx�Cb�Zq0��P�Q $JxsrtDv~r�r�w����u��rw�ԍr�wU9X!uUXEq��v !�u�u�u�q�q�y�q�wpFTF��~s8�n2��Z�e�� ��J�dPQ�Y^�D�g  � 8��R�� U�$HEI3GH��zH?(a�gV�B���R�� �c �D/ѱP$Be�x����SHIF�HRV��FPC����PC�srhqx�@�� �3p�#9�kDI�b`�CE�PV��Q�S�PHER�� �� ,a���������y@GNp�)�  ��������8`8`
8` ���IORITY �P��ʒ����$`SP�@�����ԕ��;���8�ˑגODU��x�����W�5��G�GL�H�1�H�IBHQO���TO�E�1D�  _(!AF��E ��ӯާ!tcp|ޯ�!ud��~.�!icm��V�5�XY�� ��� �ԑ)�� *������8`� ��Ϳ��������� �S�:�w�^ϛϭϔϐ�ϸ����*4�p�����%+�=�O�a� o>��/c�	�=/�� **:��哈9߮�����ض�A}��,  �ΐ�����*��`���Z��m�������ENHANCOE (���A>��d�����  �1�����ѓ����QTkR�8`���>RTREP�w�g�SKST�`㖡�wSLGu ������ԑUnothing�����  ��CUgY���TEMP D��xz�4 _a_s_eiban�	Š ����2V Azew���� ��//@/R/=/v/ a/�/�/�/�/�/�/�/ ??<?'?`?K?�?o? �?�?�?�?�?O�?&O OJO5OGO�OkO�O�O �O�O�O�O_"__F_ 1_j_U_�_y_�_�_�_<�_��VERS׀A��` dis�able��]SA�VE 	D�	�2670H700�X�_po!��ro�o/��o 	�h*�|��o�e�o�e;M_qz*|�o�9�\/gƁ 1
��]`�p'��5���'�.��URGh�Bu���h�WFA������/��W̠b�K�f�WRU�P_DELAY �����_HOT %3�,�����s�R_NORMA�LňL�Տ*���SE�MI	�/�n�֑QS�KIP�s3��sx �_���_ן�����3� "�0��P�b�t�:��� ����ί�򯸯�� :�L�^�$�n������� ʿܿ�� ���6�H� Z� �~�lϢϴ��όπ������ �2�D�3���$RACFG �����|��b�_�PARAM��3 @��@`\��|�2C���|�M��Cg�G�BbЏBTIF����b�C_VTMOU������b�DCR�s��� �ʑ=�t�B8*B�(^P@���@-�S;����￟��}վ-��T3�
�̟��ޗ�;e�m��K�Z;�=g;�4�<<���J���� �:�L� ^�p���������������� }�RDIO_?TYPE  7��u���
EDPROT-_f���C�|��BHg�E��X��2�h ���B� �Я�
������ +�\[���� ߴ����"// F/T'rw/��>/�/�/ �/�/�/�/�/�/?B? d/i?�/�?$?�?�?�? �?�?O�?,ON?SOr? $O�O O�O�O�O�O�O _�O(_JOO_nO0_
_ p_�_�_�_�_�_�_o 4_9oKo
oloo�o~o �o�o�o�o�o0o5 TohV�z�� ���@1���X?INT 2ȉ�=�q�G;� o������祐j�f�0  Ǐً����	��� S�A�w�]�������џ ����۟�+��O�=� s���k�����ͯ��� ��'��K�9�o��� g�����ɿ��ٿ����#��G�T�EFPO�S1 1'	  x���t�� �ϩ����ȈϚ���5�  �Y���}�ߡ�<ߞ� ��r��ߖ���C�U� ���<�����\��� ��	����?���c��� ��"�����X�j��� ��)��M��qn �B�f��% ��mX�,� P�t�/�3/� W/�{/�/(/:/t/�/ �/�/�/?�/A?�/>? w??�?6?�?Z?�?�? �?�?�?=O(OaO�?�O  O�ODO�O�OzO_�O '_�OK_]_�O
_D_�_ �_�_d_�_�_o�_o Go�_koo�o*o�o�o `oro�o�o1�oU �oyv�J�n ���-����u� `���4���X��|�ޏ ���;�֏_������� 0�B�|�ݟȟ���%����I��F���k�2 1w�!�3�m�� ֯��3�ίW��T� ��(���L�տp����� �����S�>�w�ϛ� 6Ͽ�Zϼ��ϐ�ߴ� =���a���� �Z߻� ����z���'���$� ]��߁���@���d� v����#��G���k� ���*�����`����� ��1������*� v�J�n��� -�Q�u�4 FX���/�;/ �_/�\/�/0/�/T/ �/x/?�/�/�/�/[? F???�?>?�?b?�? �?�?!O�?EO�?iOO O(ObO�O�O�O�O_ �O/_�O,_e_ _�_$_ �_H_�_l_~_�_�_+o oOo�_soo�o2o�o �oho�o�o�o9�o �o�o2�~�R� v���5��Y���}��������3 1��N�`�����<� B�`����������U� ޟy����&���ӟ� ���k���?�ȯc�� ���"���F��j�� ��)�;�M����ӿ� ��0�˿T��Qϊ�%� ��I���m��ϑϣϵ� ��P�;�t�ߘ�3߼� W߹��ߍ���:��� ^�����W����� w� ���$���!�Z��� ~����=���a�s��� �� D��h� '��]��
� .���'�s� G�k���*/� N/�r//�/1/C/U/ �/�/�/?�/8?�/\? �/Y?�?-?�?Q?�?u? �?�?�?�?�?XOCO|O O�O;O�O_O�O�O�O _�OB_�Of___%_ __�_�_�__o�_,o �_)obo�_�o!o�oEox�o��Ƅ4 1я {o�o�oE0ioo� (�L����� /��S�� ��L��� ��яl��������� O��s����2���V� h�z���� �9�ԟ]� �����~���R�ۯv� ����#���Я��}� h���<�ſ`�鿄�� Ϻ�C�޿g�ϋ�&� 8�Jτ�����	ߤ�-� ��Q���N߇�"߫�F� ��j��ߎߠ߲���M� 8�q���0��T�� ������7���[��� ��T�������t��� ��!��W��{ �:�^p�� A�e �$� �Z�~/�+/� ��$/�/p/�/D/�/ h/�/�/�/'?�/K?�/ o?
?�?.?@?R?�?�? �?O�?5O�?YO�?VO �O*O�ONO�OrO�O�o�d5 1�o�O�O �Or_]_�_�O�_U_�_ y_�_o�_8o�_\o�_ �oo-o?oyo�o�o�o �o"�oF�oC| �;�_���� �B�-�f����%��� I��������,�Ǐ P�����I�����Ο i�򟍟����L�� p����/���S�e�w� �����6�ѯZ���~� �{���O�ؿs�����  ϻ�Ϳ߿�z�eϞ� 9���]��ρ���߷� @���d��ψ�#�5�G� ��������*���N� ��K����C���g� �������J�5�n� 	���-���Q������� ��4��X�� Q���q�� �T�x�7 �[m�//>/ �b/��/!/�/�/W/��/{/?�/(?_ T6 1+_�/�/!?�? �?�?�/�?�?O�?O AO�?eO O�O$O�OHO ZOlO�O_�O+_�OO_ �Os__p_�_D_�_h_ �_�_o�_�_�_ooo Zo�o.o�oRo�ovo�o �o5�oY�o} *<v����� �C��@�y����8� ��\�叀�����ޏ?� *�c�����"���F��� �|����)�ğM�� ���F�����˯f�� ������I��m�� ��,���P�b�t���� ��3�οW��{��x� ��L���p��ϔ�߸� �����w�bߛ�6߿� Z���~�����=��� a��߅� �2�D�~��� �����'���K���H� �����@���d����� ������G2k� *�N�����1�U;?M47 1X?N��� �/�8/�5/n/	/ �/-/�/Q/�/u/�/�/ �/4??X?�/|??�? ;?�?�?q?�?�?O�? BO�?�?O;O�O�O�O [O�OO_�O_>_�O b_�O�_!_�_E_W_i_ �_o�_(o�_Lo�_po omo�oAo�oeo�o�o �o�o�olW� +�O�s��� 2��V��z��'�9� s�ԏ���������@� ۏ=�v����5���Y� �}�����۟<�'�`� �������C���ޯy� ���&���J����	� C�����ȿc�쿇�� ���F��j�ώ�)� ��M�_�qϫ����0� ��T���x��u߮�I� ��m��ߑ������� �t�_��3��W��� {������:���^���x��hz8 1� /�A�{�����#�A ��e b�6�Z �~��� a L� �D�h� /�'/�K/�o/
/ /./h/�/�/�/�/? �/5?�/2?k??�?*? �?N?�?r?�?�?�?1O OUO�?yOO�O8O�O �OnO�O�O_�O?_�O �O�O8_�_�_�_X_�_ |_o�_o;o�__o�_ �oo�oBoTofo�o �o%�oI�omj �>�b���� ���i�T���(��� L�Տp�ҏ���/�ʏ S��w��$�6�p�џ ���������=�؟:� s����2���V�߯z� ����د9�$�]����� ���@���ۿv����� #Ͼ�G�����@ϡ� ����`��τ�ߨ�
� C���g�ߋ�&߯ߕ����MASK 1����������XNO  �� ��?MOTE  "���X�_CFG �_��Tԓ��PL_RANG[�WѶ�����OWER ������SM_�DRYPRG �%���%\����T?ART ���UME_PRO�����v���_EXEC_ENB  ����GSPDO���;��TDB�����RM����INGV�ERSION �#�e���I_A�IRPUR�� pW�0�l��MT_���T��]����OB�OT_ISOLC� ��h ����N�AME�-��OB_CATEG ���1�$�8@O�RD_NUM ?���eH?700  T�{�����PC_TI�MEOUT�� x���S232x�1 �#��� LT�EACH PEN�DAN�tד�$�[�Y����� ���� c�e ConsT��/-&"'/U�мֳ e-W//K�?No Us�/�/8�/�NPO)��������C7H_LR�!����	F1?!UD�1:l??R��VA�IL\�T ����PACE1 2="#�
?���,zӑ��U i)L�< ��0?� �;PO�?0O�O�O~O�O �G�?�?OO�O>O`O V_w_6_�_�_�]#�#� �]�O�O__�_B_d_ Zo{o:o�o�o�o�o�O �_oo,o�oPoroh �o�����o�o (�Lnd���D� ������Џ� ��$� 6�H�Z�|�r�@����� ɟ������ �2�� V�x�n���N���ů�� گ��
��.��R�d� j���J����������� ��*�<��`���x� ��HϺ��϶����� &�8���\ώ�t���T�@���ߢ���;�12�<� �?�*�<��� `ߒߕ���u���������3�'�9�K�]� ������������"#�46�H�Z�l� ~�0������.CD5Wi{ ��Q���>� ./O/&/d/e6x� ���r/�/?_/@�/O?p?G?�?�/7�/ �/�/�/�/�??7?:O��?OpO�OhO�O�?8 �?�?�?�?O�O&OXO [_�O;_�_�_�_�_�O�G &�K t�_�
(` o  �EHoZolo~o�o �o�o�CX�m_�_�o�_2�dHp-o?om ������o�o �n�z!�3�P�CU� ������ˏݏ��� 	��=�O�p�c�u��� ��ǟٟ������p)�;�]�o� `�_ @Ш�������������� ����*�l�~���R��� ƿؿ�������2��� ��JόϞϼ�rϤ� �����������R���"�
֯���_MODE  �IR��/S '�K��L��J�/_ү��M�r�	�m��+�CWORK�_AD����n�-�R  �K��@������_INT'VAL��T��C��OPTION� ��N V_DA�TA_GRP 2Y)(��AD��P�� o���~��������� ����,<>P �t������ (L:p^� ������/ / 6/$/Z/H/j/�/~/�/ �/�/�/�/�/?? ? V?D?z?h?�?�?�?�? �?�?�?O
O@O.OdO ROtOvO�O�O�O�O�O _�O*__:_`_N_�_����$SAF_D?O_PULS�����/�c�Q�PCAN_GTIM�ў�0��Q�R */䈿0���&`&b,��AA�cK��Q�� �� 6oHoZolo~o�oo�o��o�o�o�o��o��b27t�Q�Qd�Cx:qJq���Sy ��������fyz� \��t��_ ��  T�����#�5�B�T D��B�k�}�������ŏ ׏�����1�C�U��g�y����&�xz���ڟ쟱�  }@�;�o���
�K�p���
�t��Dik�a7�  � ��b��e �Q��F���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ���������� �2�D�N���r߄� �ߨߺ��������Q� %u.�@�R�d�v���@���������0�r \�S�h���!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������\�/ '/9/K/]/o/�/�/�/ �/"��/�/�/?#?5? G?Y?k?�����b�? �?�?�?�?OO)O;O MO_OqOI�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxoM�衟Q��o�o�o�o �o,>Pbt��������zp�o�$�.����2���	123�45678s�h�!B!�� +
F��`���� ����ʏ܏� ��$� *��oM�_�q������� ��˟ݟ���%�7� I�[�m�~�<�����ů ׯ�����1�C�U� g�y������������� ��	��-�?�Q�c�u� �ϙϫϽ�������� �ֿ;�M�_�q߃ߕ� �߹���������%� 7�I�[�m�,ߑ��� ���������!�3�E� W�i�{����������� ����/ASe w������� ��=Oas� ������// '/9/K/]/o/.�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�?����?�?�5�/O�1OCO_�Cz  �A��j   ���h2�}� >OF
�G�  	��2�?�O�OH�O�O\�oL��O R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o7_�o�o�o &8J\n� ���������"�4�B�A�A�B<�_� U��A  �o���sCu@�l��A�At  �v@��ŏ�@(ۃ `�Rl����iMu@0\��$SCR_GRP� 1,0+�04� � �ވB |E	 �`�� h�y�r��^�~E����������ڟRM��@גD�#\���כ0\CRX-�10iA 012�34567890J�@N� \��@N�30 k��A
X����	���K �� h��W���W�0S^�בv�����	�����*�<�N�^���#H����l�W��������ſ׿���o�A ��Ϯ�?�XG0�w�\C�h_@,[}xx � �䄑B�  CBƊψ¡Ą�Av@���  @�@�ń�@9����� ?��Ǆ��H��߳ʄ�F@ F�`+�3�*�W� B�{�fߋ߱ߜ����� �ߤ�������$��!�3�E�B�S��ߙ�� �����������;� &�_�J�����/^�ß����|G�@���@I���e@M B�bX������?�TA�������� 0Q��A ����/�pDPb1 (�@�(����{��� /)L����='�£�7�ECLVL�  Q   ���Ǣ� Q@P!L_D?EFAULTX$L!_��@l#?HOTSTRx-���"MIPOWER�FW ZE�%�$W7FDOy& �%6��ERVENT 1�-_!_!�# L!�DUM_EIP�/8�j!AF�_INEx =?T!'FT?l>3?�?9!���? �?�?�!RPC_MAIN�?�8��?(O�3'VIS�?�9�OtO!OPCUAuO�JcO�O!TMP�@PU�O&9d�O�_!
PMON_�PROXY_)6e �OX_�B&_"=fG_�_�!RDM_SR�V�_&9g�_�_!�R��o'8h�_<o!%
�0Mo_#<i+o�o�!RLSYNC̉o�i8wo�o!gROS?�l�4�o� !
CE�@MT'COM!)6kl{!	5rCONSm�(7l[�!5rWOASRC�_)6m�v�!5rUSB��'8n�P�!STM� j�%:o?����?����S����#ICE�_KL ?%�+� (%SVCPGRG1�1��21�D6� �3Y�^� �4��D�� �5���� �6џ֟ �7���� �y�A�<�9I�N��ov�  �#��� �K�Ư �s� � ���� �ß>� � �f� ���� �;���  �c�޿H����H��� .�H�ܯV�H��~�H� ,���H�T���H�|��� H����H�̿F�H��� n�p��� � ��� ����@��&��J�5� n�Y��}������� �����4��X�C�j� ��y������������� 0T?xc� ������ >)bM���� ���/�(//:/�^/I/�/�_DEV� �)�U�T1:�'4��~�$GRP 21�%�� �bx 	_� 
 ,� �/ ?�"�/.??R?9?K? �?o?�?�?�?�?�?O �?*O<O#O`OGO�O�O �/�OqO�O�O�O_�O 8_J_1_n_U_�_y_�_ �_�_�_�_o"o	oFo �O;o|o3o�o�o�o�o �o�o�o0T; x�q����� �_o,�>�%�b�I��� m��������Ǐ�� ��:�!�^�p�W���{� ��ʟ!���$�� H�/�l�~�e�����Ư ������� ��D�V� =�z�џo���g�Կ�� ��
��.��R�d�K� ��oϬϾϥ������ ����<ߓ�`�r�Yߖ� }ߺߡ߳�������� 8�J�1�n�U���� �������U�"���F� X�?�|�c��������� ��������0T; x�q����� �,>%bI� ������/��:/!/3/p/�#d Խ&	^/�/�/�/�/0�/�/?";%�"?G?�#���`11`5 p?~7h?�?�?�?�?�? �94?O\9�?FO4OjO XOzO|O�O�OO�O*O �O__B_0_f_T_v_ �O�O�__�_�_�_o o>o,obo�_�o�_Ro �oNo�o�o�o: |oa�o*���� ����T9�x� l�Z���~�����ď� ,��P�ڏD�2�h�V� ��z����ן韠� ��
�@�.�d�R���ʟ ���x��Я���� <�*�`�����ƯP��� ��޿̿���8�z� _Ϟ�(ϒπ϶Ϥ��� ����@�f�7�v��j� Xߎ�|߲ߠ������ <���0���@�f�T�� x����������� ,��<�b�P������ ��v�������( 8^�����N�� �� �$fK] 6~���� �>#/b�V/D/f/ h/z/�/�/�//�/:/ �/.??R?@?b?d?v? �?�/�??�?O�?*O ONO<O^O�?�?�O�? �O�O�O_�O&__J_ �Oq_�O:_�_6_�_�_ �_�_�_"od_Io�_o |ojo�o�o�o�o�o�o <o!`o�oTBxf �����8� ,��P�>�t�b���� ��я�������(�� L�:�p�����֏`�ʟ ��ڟܟ�$��H��� o���8�����Ư��֯ د� �b�G����z� h�����¿��ҿ(�N� �^���R�@�v�dϚ� �Ͼ� ���$Ϯ�ߪ� (�N�<�r�`ߖ��Ͻ� �φ�������$�J� 8�n�ߕ���^���� ������� �F���m� ��6������������� N�3E����f �����&J �>,NPb�� ���"�//:/ (/J/L/^/�/��/� �/�/�/? ?6?$?F? �/�/�?�/l?�?�?�? �?O�?2Ot?YO�?"O �OO�O�O�O�O�O
_ LO1_pO�Od_R_�_v_ �_�_�_�_$_	oH_�_ <o*o`oNo�oro�o�o �_�o o�o8& \J��o��p� l���4�"�X�� ��H�����ď֏ ���0�r�W��� ��� x���������ҟ�J� /�n���b�P���t��� �����6��F��:� (�^�L���p����Ϳ ��� ϒ��6�$�Z� H�~������n����� �����2� �Vߘ�}� ��F߰ߞ��������� �.�p�U����v� ��������6��-� �����N���r����� �����2���&6 8J�n����
 ���"24F |���l��� �//./��{/� T/�/�/�/�/�/�/? \/A?�/
?t??�?�? �?�?�?�?4?OX?�? LO:OpO^O�O�O�O�O O�O0O�O$__H_6_ l_Z_|_�_�O�__�_ �_�_ ooDo2oho�_ �o�oXozoTo�o�o�o 
@�og�o0� �������Z ?�~�r�`������� ������2��V���J� 8�n�\���������� �.�ȟ"��F�4�j� X���П����~��z� ����B�0�f����� ̯V������ҿ��� �>π�eϤ�.Ϙφ� �Ϫ��������X�=� |��p�^ߔ߂߸ߦ� �����������6� l�Z��~������� ������ �2�h�V� �������|�����
 ��.d����� T����� l�c�<��� ���/D)/h� \/�l/�/�/�/�/�/ /?@/�/4?"?X?F? h?�?|?�?�/�??�? O�?0OOTOBOdO�O �?�O�?zO�O�O_�O ,__P_�Ow_�_@_b_ <_�_�_�_o�_(oj_ Oo�_o�opo�o�o�o �o�o Bo'fo�oZ H~l���� �>�2� �V�D�z� h�����׏���
� ��.��R�@�v����� ܏f�Пb������*� �N���u���>����� ̯��ܯ��&�h�M� �����n�����ȿ�� ؿ��@�%�d��X�F� |�jϠώ�������� ���ϰ��T�B�x�f� ������ߌ������ ��P�>�t�ߛ��� d����������� L���s���<������� ��������T�z�K�� $~l����� ,P�D�Tz h����(� /
/@/./P/v/d/�/ ��/ /�/�/�/?? <?*?L?r?�/�?�/b? �?�?�?�?OO8Oz? _OqO(OJO$O�O�O�O��O�O_RO7_vO�A��$SERV_MA_IL  �EvP��\XOUTPUT�kX�@@�`TRV 22 V  yP (QF_�_�`TSAVE�\zYTOP10 23�Y d |O2oDo Vohozo�o�o�o�o�o �o�o
.@Rd v������� ��*�<�N�`�r��� ������̏ޏ�����&� UeYP�_]SF�ZN_CFG 4 UyS{D�Q��Uf�GRP 25�p��Q ,B  � A���AD;� �B���  B4~&cRB21�VoHELLi�6 U��V�P�_���(�%RSR(�)�;�t� _����������˯ݯ ��:�%�^�I���������  ��Q%��Կ濡�������@����zG��2�@d���ۖ�HK 17� ϚϕϧϹ����� ���*�%�7�I�r�m߀ߑߺߵ�����՜OMM 8�)�ڒ�FTOV_ENB�kT�Q�YHOW_R�EG_UII�^RIMIOFWDL��9~�WAIT�F�Ɉ���Pj�ܳT��TIMj������VAjP��~�_�UNITE���YL]Cc�TRYj��U-`PMEi�:���Q�	���f�;r� �������<�����X�@Đ `	P?�  �����_'�P@6��V�VMON_AL�IAS ?e��Phe1_���� �
�%7�[ m��N��� �/�3/E/W/i/{/ &/�/�/�/�/�/�/? ?/?A?�/e?w?�?�? �?X?�?�?�?OO�? =OOOaOsO�O0O�O�O �O�O�O__'_9_K_ �Oo_�_�_�_�_b_�_ �_�_o#o�_GoYoko }o(o�o�o�o�o�o�o 1CU y� ���l��	�� -��Q�c�u���2��� ��Ϗ�󏞏�)�;� M�_�
���������˟ v����%�П6�[� m����<���ǯٯ� ����!�3�E�W�i�� ������ÿտ����� �/�ڿS�e�wωϛ� FϿ�������߲�+� =�O�a�s�ߗߩ߻� ��x�����'�9��� ]�o����P����� �������5�G�Y�k� }�(������������� 1C��gy����Z�$SMO�N_DEFPRO�G &����� &�*SYSTEM*����RECAL�L ?}�	 (� �}4xcop�y fra:\*�.* virt:�\tmpback�?=>192.1�68.56.1:?11320 fm���}86s:�orderfil.datCUk��/ /}/6mdb:@�g�v/�/�/�35>Pbi/�/ ??�4�/�/�/{? �?�?��M/h/�?O O0/�?T/�?wO�O�O �/A?S?�/�O__,?��O�Ob?s_�_�_�77�5Fhome.tpCUemp\�TU_k_ �_oo�?�?MO�_yo �o�o0OKoTOfo�o	 �OA_S_�Ou�� ,_=Ob_���*g�\�d:ipl_f�anuc_smp�lgrp_close.ls�Y=�O� ����3oEo�o�rn� ܏��o�oя�o�Q� �"�4�Xj�|��� ��ß���s�X������tpdisc 0}��pR�d�v�������tpconn 0 ��Я��� ���*���=�O�a�s� ��ϩ���D�ߏ�� ��'�9�T�]�oρ�� ����J�۟��V�!�#� 5�F�ٿk��ߏ� ﳯ ſ?�������1�7�1}�O�a�s���)� ;���_�������Ϲ� T���o���%�7��� [���V!�ߵ�F�� k�� 3�E���i ����L��gy �//��e�	/ �/�>/P/�u/�/?�+�95�anima�tion_pick�\�/�p�/?�?%?7=dropK?�?o?@�?O%7I�? �? \O�O��QO�lO�O��O!^�$SNPX�_ASG 2<����@Q�� P 0 '�%R[1]@g1.1!_kY?�-�%k_�_z_�_�_�_�_ �_�_'o
oKo.o@o�o do�o�o�o�o�o�o �oG*kN`� �������1� �;�g�J���n����� ��ˏ��ڏ����Q� 4�[���j�������� ğ����;��0�q� T�{�����˯����� ��7��[�>�P��� t���ǿ���ο�!� �+�W�:�{�^�pϱ� �ϻ�������� �A� $�K�w�Zߛ�~ߐ��� �������+�� �a� D�k��z������ ����'�
�K�.�@��� d������������� ��G*kN`� �������1 ;gJ�n�� ����/�/Q/ 4/[/�/j/�/�/�/�/ �/�/?�/;??0?q? T?{?�?�?�?�?�?O��?O7OD3TPAR�AM =@U�JQ �	�;JP��D�@�H�D�� ��3POFT�_KB_CFG � zCFU0SOPI�N_SIM  @[�F�O�O_�@Q@�RVNORDY_�DO  �E�E�%RQSTP_DS�B�N�Bi_uHQ@S�R >�I �� & IPL_�FANUC_SM�PLGRP_OPENu]yD�@Q@�TO�PN_ERR�2_OB�QPTN ��E
`�D��RRING_PR�M�_DRVCNT_�GP 2?�E�A�@x 	e_do|@Ro��ovo�o�WVD9`ROP 1@`I�@�a �I�g�o�o 2Y Vhz����� ����.�@�R�d� v������������ ��*�<�N�`�r��� ������̟ޟ��� &�8�J�q�n������� ��ȯگ����7�4� F�X�j�|�������Ŀ ֿ������0�B�T� f�xϊϜ��������� ����,�>�P�b߉� �ߘߪ߼�������� �(�O�L�^�p��� �����������$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@gd�v�����bPRG_COUNT�Fs�
b�ENBo��M#�D/_UP�D 1A�[T  
�{Bf/x/�/�/ �/�/�/�/�/??C? >?P?b?�?�?�?�?�? �?�?�?OO(O:OcO ^OpO�O�O�O�O�O�O �O __;_6_H_Z_�_ ~_�_�_�_�_�_�_o o o2o[oVohozo�o �o�o�o�o�o�o
3 .@R{v��� ������*�S� N�`�r���������� ޏ���+�&�8�J�s� n���������ȟڟ������_INFO� 1BT%: \�	 3�w�b������?*&�?����>Y�L=��n-�����h>F��d9��]/������>�@ ?�ݸ)�<@� �D&t�����D)�´ �²E�³���*�<��YSDE�BUG�U �*�d�=)e�SP_PAS�S�B?w�LO�G CQ�^! � *�#�0�  ��9!*�UD1�:\��7���_MPAC��T%%�7�T!��U� T!�SAV D��!��̱�$���SV��TE�M_TIME 1�E��_  0 7 L(��#�����ù�MEMBK  T%9!̰̿9߼K�[�X|: � �'��}ߢ߲��v�������r� ��@���,�>�P�Àh�z�������� �������0�B�T�f�x����e������ ����*<N` r���������SK���`$�Tfxl�n*�EX�2�߷#� ��p)�����������</N/`/7.e�*�� ��/�$���/�/8�/���2�?;? M?_?q?�?*�U�?�? ���?'���?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_@��T1SVGUNS�PD�� 'w���HP2MODE_LIM F��{�DT�2QPqQG��CUA�BUI_DCS J7w�F�'�_ �$�$G�6_�\o�WG�o*���9a 
?`H�9o'�Sh��Sc�ɼ�UEDIT �K�_�XSCRN������R�G �M�[�U�:�eSK_OPTIONl���{��b_DI��ENB  �%w��a�BC2_GRP 2N�Y���o��0�C��s<\BCCF2�`P]{�� ����v`�����!� G�2�k�V���z����� ׏ԏ���1��U� @�y�d�������ӟ�� �����?�Q�g^� p�������0�ٯį� ���3�a�N��#�V� |�j�����Ŀ���ֿ �����B�0�f�Tϊ� xϮϜϾ�������� ,��P�>�`�b�tߪ� �؆`������ ��� 6�$�F�l�Z���� ���������� ��0� 2�D�z�h��������� ������
@.d R�v����� ��0N`r� ������// �8/&/\/J/�/n/�/ �/�/�/�/�/�/"?? F?4?V?|?j?�?�?�? �?�?�?�?�?OBO0O fO~O�O�O�O�OPO �O�O_,__P_b_t_ B_�_�_�_�_�_�_�_ �_o:o(o^oLo�opo �o�o�o�o�o �o$ H6XZl�� �|O��� �2�� V�D�f���z���ԏ ������
�@�.�P� R�d����������П ����<�*�`�N��� r���������̯�� &��>�P�n������ ����ƿ�ڿ�"�4� �X�F�|�jϠώϰ� ����������B�0� f�T�vߜߊ��߮��� �������,�b�P� ��<����������p� ��&�L�:�p����� b��������� �� $ZH~l�� ����� D 2hVxz��� ����/./@/R/� v/d/�/�/�/�/�&� ��$TBCSG_�GRP 2Q�%��  ���! 
 ?�  ?+??O?9?s?]?�o?�?�?�?�;�"�#S~ <d�HA�?�!	 HA�����5>���>��=q?�\�5AT��A 2HOTH�J�ff?aG��?L G>BpTOVN��t@#E� @wA� 6J���O�M@��RjI>G�33*A�5�ABCO��O�H�BPOQY�,_.^��HBY�ArBU�PB�t_.^�H�6 �H�U�_�_�_ o=oo�oho�o�kjh��a	�V3.002	Ocrx�c�`*�`p�d�"8T�O ?�S2� Hqji p�mn  �3C�oXY`s�!J2�#T =�`lxCFG -V�%
1 0�z+��r,r��x����� � E�0�i�T���x����� Տ��ҏ���/��S� >�w�b�������џ�� ������=�(�:�s� ^�������ͯ2+ د �����/��?�e�P� ��t�����ѿ���� ¿+��O�:�_υ��! �/�϶/�ϼ������ (��L�:�p�^߀ߦ� ���߸������ �"� $�6�l�Z��~��� ���������2� �V� h�(/����<������� ����
@.Pv ��X����� *<Nr`� ������// 8/&/\/J/l/�/�/�/ �/�/�/�/�/??"? X?F?|?j?�?�?�?�? �?�?��O$O6O�?fO TOvOxO�O�O�O�O�O __,_>_�Ob_P_�_ t_�_�_�_�_�_�_o o:o(o^oLo�opo�o �o�o�o�o �o$ H6X~l��� ������D�2� h�V�����HO��ȏ�� ��
���.��R�@�b� d�v�����П����� ��*��N�`�r���>� ����̯��ܯ��&� �J�8�n�\�~����� ȿ���ڿ���4�"� D�j�Xώ�|ϲϠ��� ��������0ߪ�H�Z� l�ߜߊ߬������� ����>�P�b�t�2� ����������� ����L�:�p�^����� ���������� 6 $ZHjl~�� ���� 0V Dzh����~� ���ߺ@/./d/R/ �/v/�/�/�/�/�/? �/�/<?*?`?N?�?�? �?�?t?�?�?�?�?O 8O&O\OJO�OnO�O�O �O�O�O�O�O"__F_ 4_V_X_j_�_�_�_�_ �_�_o�_oBo0ofo �/�o�oLozo�o�o �o,P>t� ��h����� (�:�L�^����p��� ��ʏ��ڏ܏�$�� H�6�l�Z���~���Ɵ ���؟���2� �B� D�V���z�����ԯ¯ ��
��o"�4�F��v� d�������������� �*�<�N��r�`ϖ�8�ϺϤ�  ����� �������$�TBJOP_GR�P 2W����  ?�/��C��	���Y�����X  ���Y� �,� � �x���� @��?}�	 ߐA��͔�C��  D�ǌь�>~0�>\?�����aG�:�o���;ߴAT�ͰՌ�A��Ӭ����ߦ�>�я\)�?��D�8Q�|�Ѵ�L��>���^��;iG�Ҍz��Ap�Љ� ��A�ff��0��m�����^��:VM��ҹR�����)���@��RD�Cр��щ�i��e�H�Q��ff��:w�6/D�33��B   �����D��V�h�Q�Q�x���:�cS���}�,B�6<?Q@��Hd���r����d�=m�<#��
���0�;/�e�d���B�� ���ٰ��"�� :kF ��� �����/4//�,/Z/�/��C��Ɛ��!��	V3.0=05�crx�#� �*� i�������*� C�  E$�` E�h E��� F� F3�� FV4 Fx�� F�� F�� F�X F��0�� F�F �F�� Gs �G G� Gk G&�#��� Y? E@ �E�� E�� �E� F� �F2 FN� �Fj� F�� �F�� F� �F�H F�| �Fʰ 9�IR$�1t,H�5 *���?*�2���3?����`-�ED_TCH� Z��(�#�2���h���d$�(�O�O��� �TES�TPARS  ���SC�HR�@AB�LE 1[� A@��fւҞG�:
�G�H�H�����G	�H
�H�HU��U�H�H�H�F'RDI�O(�__ %_7_I_[U�TO�_�[@�_�_oo/n�BS�_&� �Z�o&8 J\n����� ����"�4�F�� �`�o'� W��po�o�o �oR_d_v_�_�_�X�B~m�NUM  �ū(�p��� ��@�P�B_CFG �\V����@�IMEBF_TT�At��PE��VER�S�fѮ���R 1]��K 8zO��d��� ����  � ��)�;�M�_�q��� ������˯ݯ��� %�7���[�m������� ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/�x�S� e߮߉ߛ߱߿����ߐ���:Bۑ_P�Ŗ@�ϕ<@LIF M^V��0ʑ������"��( 0
�:�@��@� d��W�MI_CHAN��� ϕ ��DBGL�VL��PF��ET�HERAD ?�E����0��7��I���ROUT�!HJ!}�����SNMASK�ϓ$�255.���#��������#<@OOLOFS_DI�@R0�����ORQCTRL� _�K;c�?yT h������	 -?Qcu�� ���g��/9C�PE_DETAI���>
PGL_CONFIG eV��f���/cel�l/$CID$/grp1/�/�/�/�/�/6c�d�??%? 7?I?[?�/?�?�?�? �?�?h?�?O!O3OEO WO�?�?�O�O�O�O�O �OvO__/_A_S_e_ �O�_�_�_�_�_�_r_ �_o+o=oOoaoso��}o�o�o�o�o�o�/+
}�o`r ����o��� �&�8��\�n����� ����ȏW�����"� 4�F�Տj�|������� ğS������0�B� T��x���������ү a�����,�>�P�߯ t���������ο�o� ��(�:�L�^��� �Ϧϸ�����k� ���$�6�H�Z�l�g ��User Vi�ew |)}}12�34567890 �߯�����������2�,}������2���� a�s������,���3D�	��-�?�Q�c����2�4����������v�82�5 ��q�����*�2�6`%7I[ m��2�7� ��/!/3/�T/2�8��/�/�/�/�/�/�F/?2 lCamera�� �/M?_?q?�?�?�?�bE@?�?�?�>��O!O`3OEOWOiO_	  '6 C�<?�O�O�O�O__ �?7_I_[_�O_�_�_�_�_�_ ?�'6��p_ %o7oIo[omoo&_�o �o�oo�o�o!3 E�_�W���o��� ����o�!�3�~ W�i�{�������X�W �KJ����#�5�G�Y�  �}������şן� ����Ə(5��i� {�������ïj���� �V�/�A�S�e�w��� 0��W� �տ���� �/�֯S�e�w�¿�� �Ͽ������Ϝ��W{) ��A�S�e�w߉ߛ�B� ������.���+�=�O�a���9�ߢ�� ����������2�D� ��U�z�����������
c*	)50Z�!3 EWi����X� ���/���� .00;������ ��//*/uN/`/ r/�/�/�/O)5�K?/ �/??*?<?N?�r? �?�?�/�?�?�?�?O O�/��k�?`OrO�O �O�O�Oa?�O�O_MO &_8_J_\_n_�_'O9E t{_�_�_�_oo&o �OJo\ono�_�o�o�o �o�o�o�_9E���o8 J\n��9o�� �%��"�4�F�X� �o9EL������ȏڏ ����"�4�F���j��|�������ğk�  o����)�;��M�_�q��������� �  ə?fffB�Pߡk�����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h� zߌߞ߰����������
��.���
k�( � ��( 	 ;�q�_����� ���������7�%�[��I����� � �������[�0 BTfm������ ����� 2y Vhz����� ��?/./@/�d/ v/�/�/�/�///�/ ??_/<?N?`?r?�? �?�/�?�?�?%?OO &O8OJO\O�?�O�O�O �?�O�O�O�O_"_iO {OX_j_|_�O�_�_�_ �_�_�_A_o0oBo�_ foxo�o�o�o�oo�o �oOo,>Pbt ��o�o���'� �(�:�L�^������ ���ʏ܏� ��$� k�H�Z�l��������� Ɵ؟�1�C� �2�D� ��h�z�������¯	� ���
�Q�.�@�R�d� v���ϯ����п������*�<�Nϕ�u�@� p�}Ϗϡ�p��w�[��� frh�:\tpgl\r�obots\cr�x��10ia.xml]���� �2�D��V�h�zߌߞ߰�  ����������� � 2�D�V�h�z���� ��������
��.�@� R�d�v���������� ����*<N` r�������� &8J\n� �������/ "/4/F/X/j/|/�/� �/�/�/�/�/??0? B?T?f?x?�?�/�?�? �?�?�?OO,O>OPO�bOtO�O�N���� w���<< �� ?��K�O�O �O�O#_	_+_Y_?_q_ �_u_�_�_�_�_�_o �_%oCo)o;o]o�o�����(�$TPG�L_OUTPUT� h�����` �jfffB4  �a���o
 .@Rdv�� �������*��<�N�`�r����� ���`cell/f�loor/wal�l rite 3�456789012��ʏ܏� ���� �`�/�A�S�e�w�� !�����џ������}�6�H�Z�l�~�� (���Ưد������ �D�V�h�z���$��� ¿Կ���
Ϣ���@� R�d�vψϚ�2Ϩ��� �����߰�&�N�`� r߄ߖ�.�@������� ��&��4�\�n�� ���<��������� "�����X�j�|����� ��J�������0 ��>fx���F~�b $$zb ����:,^ P�t����� �//6/(/Z/L/~/ p/�/�/�/�/�/�/?}�A(?:?L?^?p?�?=@�O�?�?�J ( 	 ?�?�? "OOFO4OjOXOzO|O �O�O�O�O�O_�O0_ _@_f_T_�_x_�_�_ �_�_�_�_�_,ooPo����  <<?�o�o�`to�o�o �o�o��qo7I�o UYk��%� ���3�E��i�{� �c���K������ӏ �/����e�w���� �������A�S��+� ş3�a�;�M������ ͯ߯y�˯���K� ]���e���-��ɿۿ �����o���G�Y�� }Ϗ�iϗ���#ϭ��� ߧ�1�C��/�y��� �ϯ���[��������� -�?��C�u��a�� �������Q���)��� �_�q�K�������� ������%��1[ ������=��� �!EW�C��gy��gb)�WGL1.XML��?
-�$TPOF?F_LIM l`�0�ha�&Nw_SV    �4�2*P_MON �ide4$�0��02)STRTC�HK jde2&�%?"VTCOMP�ATG(�!6&VWV_AR kg-�(.K$ �/ ?�0�z"!_DEFPROG %�)�%IPL_F�ANUC_SMP�LGRP_CLO�SE�/?0ISPL�AY' �.<2INST_MSK  �<� x:INUSsER�/~4LCK�<��;QUICKMEyN�?~4SCRE@�de�"tpsc~4�1.@3I2"D@�_HIST�*2)RA�CE_CFG Ulg)�$0	4�
?��HHNL C2mK:D`�A�+ !2 �O�O__/_A_S_e_�wZ�EITEM 2�n�K �%$1�23456789y0�_�U  =<�_x�_�_c  !
ok0�_Wo3�_xo �_�o�oo�o6oHo lo,�o<b�o�o�o �o �D��(� �L����N���� ʏ܏@��d�v���� Z���~���􏜟�*� �N��r�2�D���Z� ̟����¯&�ү�� 
�n��������0�گ ������"��F�X�j� �Ϡ�`�r�ֿ~��� ���0���T��&ߊ� <߮��ω��Ϥ�ߴ� ��`�P�b�tߎߘ�� ��h������(�:� L���p��B�T���`� ���� �����6��� l�����k����� �� �D�z :�Jp���
 .�R�$/6/� Z/���f/~//�/ �/N/�/r/�/M?�/h? �/�?�??�?&?8?OʍDS�Bo�OJ�g  �RJ �A]OT9
 jO�OwO��O5JUD1:\��L��AR_GR�P 1p�[� 	 @�@_[�_>_,_b_P_�_t^� �P�_�Z�Q�O�_�_	o�U?�  $o6k o VoDozoho�o�o�o�o �o�o�o
@.dRt�	�5��~CSCB 2q"K o��0�B��T�f�x�����LUT�ORIAL r�"K�O�GV_CONFIG s"M�AZO�OF���OUT?PUT t"I7���R������� ̟ޟ���&�8�J� \�n�4���������̯ ޯ���&�8�J�\� n��������ȿڿ� ���"�4�F�X�j�{� �Ϡϲ���������� �0�B�T�f�x߉Ϝ� ������������,� >�P�b�t�ߘ��� ��������(�:�L� ^�p������������ �� $6HZl ~��������  2DVhz� ������
// ./@/R/d/v/��/�/ �/�/�/�/??*?<? N?`?r?�? �2����? �?�?�?
OO.O@ORO dOvO�O�O�/�O�O�O �O__*_<_N_`_r_ �_�_�O�_�_�_�_o o&o8oJo\ono�o�o �o�_�o�o�o�o" 4FXj|���o ������0�B� T�f�x��������ҏ �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@�R��d�v߈ߚ߬ߏ8��������Ѷ�� �?,�>�P�b�t��� ������������(� :�L�^�p��������� ������ #�6H Zl~����� ��2DVh z������� 
/./@/R/d/v/�/ �/�/�/�/�/�/?? )/<?N?`?r?�?�?�? �?�?�?�?OO%?8O JO\OnO�O�O�O�O�O �O�O�O_!O4_F_X_ j_|_�_�_�_�_�_�_ �_oo/_BoTofoxo �o�o�o�o�o�o�o +o>Pbt�� �������%���$TX_SCR�EEN 1u����М}�ipnl/Y�gen.htm%�x���𜏮���/pPa�nel setupČ}�ď��)�;�M�_��鏖��� ��̟ޟ�g����8� J�\�n�����	��ȯ گ����"���ǯ�� j�|�������Ŀ;�� _���0�B�T�f�ݿ ￜϮ���������m� �ϑ�>�P�b�t߆ߘ� ߼�3�������(��:��(�UALRM_MSG ?E��R� S�(z��� �����������;��A�r�e�������n�S�EV  |����l�ECFG �wE�O�  �(u@�  A �  B�(t
  ��/sE�Oas�� �������GRP 2x; 0(v	 9[�n�I_BBL_N�OTE y
T��l/r�J�/q nDEF�PROx�%|� (%���2p���  //D///h/S/y/�/��/�/�/�/dFKE�YDATA 1z<E�Ep (vHK?]?4?�?�?j:�,(�?�?(t([ INST ]�?��>  ��� ��Z���?�>:OLO�E�һ�� eσb�vRO�:[EDCMD�?�O8@���� Əڂ����O,O�O�O�O #_
_G_Y_@_}_d_�_��_�_�_�_�_f>���/frh/gu�i/whitehome.pngo`Io[omoo�o�"finst4o�o�o�o��o�g  FRH�/FCGTP/wzcancel�o N`r��%s��������%nex�oS�e�w������d}"fedcmdC� F�ڏ����"�-�#earwrgB�Y�k� }������şן��� ����C�U�g�y��� ����>�ӯ���	�� -���Q�c�u������� :�Ͽ����)�;� ʿ_�qσϕϧϹ�H� ������%�7�o�� m�ߑߣߵ������� ���!�3�E���i�{� ��������d���� �/�A�S���w����� ������`���+ =Oa������ ��n'9K ]������� �|/#/5/G/Y/k/ ��/�/�/�/�/�/x/ ??1?C?U?g?y?? �?�?�?�?�?�?�?O@-O?OQOcOuOl�K��`�����O�O�M�O�O_�F, �_5_�_Y_@_}_�_v_ �_�_�_�_�_o�_1o Co*ogoNo�o�o�o�o �o�o�o	?& cuTߙ���� �O�)�;�M�_�q� �������ˏݏ�� ��%�7�I�[�m��� ����ǟٟ������ 3�E�W�i�{������ ïկ������/�A� S�e�w�����*���ѿ ����Ϩ�=�O�a� sυϗ�&ϻ������� ��'߶�K�]�o߁� �ߥ�4���������� #��G�Y�k�}��� ����������1� 8�U�g�y��������� P�����	-?�� cu����L� �);M�q �����Z�/ /%/7/I/�m//�/ �/�/�/�/h/�/?!? 3?E?W?�/{?�?�?�? �?�?d?�?OO/OAO SOeO�?�O�O�O�O�O �OrO__+_=_O_a_ �O�_�_�_�_�_�_�_����[������o.o@mobotoNf,`�oX�o�o �o�o�o#
GY@ }d������ ��1��U�<�y��� r�����ӏ���	�� -�?�Q�c�r_������ ��ϟ�󟂟�)�;� M�_�q� �������˯ ݯ�~��%�7�I�[� m�������ǿٿ� ����!�3�E�W�i�{� 
ϟϱ���������� ��/�A�S�e�w߉�� �߿���������+� =�O�a�s���&�� ����������9�K� ]�o�����"������� ����#��GYk }�������� 1�Ugy� ��>���	// -/�Q/c/u/�/�/�/ �/L/�/�/??)?;? �/_?q?�?�?�?�?H? �?�?OO%O7OIO�? mOO�O�O�O�OVO�O �O_!_3_E_�Oi_{_ �_�_�_�_�_d_�_o o/oAoSo�_wo�o�o �o�o�o`o�o+�=Oa8 c{�>8 ����� �}����v,Џ� ȏ9� �]�o�V���z� ��ɏ���ԏ�#�
� G�.�k�}�d�����ş ��������C�U� 4y���������ӯ�o ��	��-�?�Q�c�� ��������Ͽ�p�� �)�;�M�_�ϕ� �Ϲ�������~��%� 7�I�[�m��ϑߣߵ� ������z��!�3�E� W�i�{�
������� ������/�A�S�e� w�������������� ��+=Oas� ������ '9K]o��j� �����/5/ G/Y/k/}/�/�/0/�/ �/�/�/??�/C?U? g?y?�?�?,?�?�?�? �?	OO-O�?QOcOuO �O�O�O:O�O�O�O_ _)_�OM___q_�_�_ �_�_H_�_�_oo%o 7o�_[omoo�o�o�o Do�o�o�o!3E �oi{����R ����/�A��e��w���������я��Ӌ�������� ���B�T�.�,@���8�����͟ߟ Ɵ��'�9� �]�D� ����z�����ۯ�ԯ ���5��Y�k�R��� v���ſ������ 1�C�R�g�yϋϝϯ� ����b���	��-�?� Q���u߇ߙ߽߫��� ^�����)�;�M�_� �߃��������l� ��%�7�I�[���� ������������z� !3EWi���� ����v/ ASew��� ����/+/=/O/ a/s//�/�/�/�/�/ �/?ڿ'?9?K?]?o? �?�/�?�?�?�?�?�? O�?5OGOYOkO}O�O O�O�O�O�O�O_�O 1_C_U_g_y_�_�_,_ �_�_�_�_	oo�_?o Qocouo�o�o(o�o�o �o�o)�oM_ q���6��� ��%��I�[�m�� ������D�ُ���� !�3�W�i�{����� ��@�՟�����/��A�0C��0���l�~���h���į��,�������  �=�O�6�s�Z����� ��Ϳ�����'�� K�]�Dρ�hϥό��� ��������#�5�?Y� k�}ߏߡ߳����� ����1�C���g�y� ������P�����	� �-�?���c�u����� ������^���) ;M��q���� �Z�%7I [������ h�/!/3/E/W/� {/�/�/�/�/�/�/v/ ??/?A?S?e?�/�? �?�?�?�?�?r?OO +O=OOOaOsOJߗO�O �O�O�O�O�?_'_9_ K_]_o_�__�_�_�_ �_�_�_�_#o5oGoYo ko}oo�o�o�o�o�o �o�o1CUgy ������	� �-�?�Q�c�u����� (���Ϗ������ ;�M�_�q�����$��� ˟ݟ���%���I� [�m������2�ǯٯ ����!���E�W�i��{��������@��}��@���ܿ@� �ؿ"�4��, � e�߉�pϭϿϦ��� ���� �=�$�a�s� Zߗ�~߻��ߴ����� ���9�K�2�o�V�� ��O���������#� 2�G�Y�k�}������� B�������1�� Ugy���>� ��	-?�c u����L�� //)/;/�_/q/�/ �/�/�/�/Z/�/?? %?7?I?�/m??�?�? �?�?V?�?�?O!O3O EOWO�?{O�O�O�O�O �OdO�O__/_A_S_ �Ow_�_�_�_�_�_�_ ��oo+o=oOoaoh_ �o�o�o�o�o�o�o�o '9K]o�o� �����|�#� 5�G�Y�k�}������ ŏ׏������1�C� U�g�y��������ӟ ���	���-�?�Q�c� u��������ϯ�� ���)�;�M�_�q��� ��$���˿ݿ��� ��7�I�[�m�ϑ� � �����������!��P�#���P���L�^�p�Hߒߤ�~�,���߈������ /��S�:�w��p�� �����������+�=� $�a�H���l������� �����_9K] o���Ϸ��� �#�GYk} ��0����/ /�C/U/g/y/�/�/ �/>/�/�/�/	??-? �/Q?c?u?�?�?�?:? �?�?�?OO)O;O�? _OqO�O�O�O�OHO�O �O__%_7_�O[_m_ _�_�_�_�_V_�_�_ o!o3oEo�_io{o�o �o�o�oRo�o�o /AS*w��� ���o���+�=� O�a����������͏ ߏn���'�9�K�]� 쏁�������ɟ۟� |��#�5�G�Y�k��� ������ůׯ�x�� �1�C�U�g�y���� ����ӿ������-� ?�Q�c�u�ϙϫϽ� ������ߔ�)�;�M� _�q߃�ߧ߹����� ����%�7�I�[�m�h��hp���hp���������������, E��� i�P������������� ����AS:w ^������� +O6s�d �����/�'/ 9/K/]/o/�/�/"/�/ �/�/�/�/?�/5?G? Y?k?}?�??�?�?�? �?�?OO�?COUOgO yO�O�O,O�O�O�O�O 	__�O?_Q_c_u_�_ �_�_:_�_�_�_oo )o�_Mo_oqo�o�o�o 6o�o�o�o%7 �o[m���D ����!�3��W� i�{�������Ï�� ����/�A�H�e�w� ��������џ`���� �+�=�O�ޟs����� ����ͯ\����'� 9�K�]�쯁������� ɿۿj����#�5�G� Y��}Ϗϡϳ����� ��x���1�C�U�g� �ϋߝ߯�������t� 	��-�?�Q�c�u�� ������������ )�;�M�_�q� ��������������$U�I_INUSER  ���"��  �_MENH�IST 1{"�  (�/ ڀ)/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,1133,1A��$��({�5�5�GYk��'�8 %����~��2$5�B/T/f/�,/�71�6w/�/��/�/��,�/�ed�it�DEFAU{LT�PICK��Q?c?u?��z ?HO;ME@0ON_<?�?��?�?��<�?!>IP�L_FANUC_�SMPLGRP_CLOS�1SOeOwO�L����v�A�O�O �O�O�O�O_ �O6_ H_Z_l_~_�__�_�_ �_�_�_o�_2oDoVo hozo�o�o-o�o�o�o �o
�o@Rdv ��)����� �*��N�`�r����� ���Ȍޏ����&� 8�;�\�n��������� E�ڟ����"�4�ß X�j�|�������įS� �����0�B�ѯf� x���������O���� ��,�>�P�߿tφ� �Ϫϼ��Ϲ����� (�:�L�^�aςߔߦ� ������k� ��$�6� H�Z���k������ ����y�� �2�D�V� h�������������� u���.@Rdv �������� �*<N`r�� �����/�&/ 8/J/\/n/�/�/!/�/ �/�/�/�/?�/4?F? X?j?|?�??�?�?�? �?�?OO�?BOTOfO xO�O�O+O�O�O�O�O�__�$UI_�PANEDATA 1}���KQ�  	��}  ttp://127.0hP�1:3080/f�rh/jcgtp�/flexdev�.stm?_wi�dth=0 &_�lines=15�&_column�s=40&_fo�nt=24&_p�age=whol�e�P'_)  r3im�_�_  \P
o o.o@oRodo�_vo�o �o�o�o�o�o�o�o <N5rY������ � � �p%#t\ o	��-�?�Q�c�� ���_����Ϗ��� l�)�;�"�_�F����� |�����ݟ�֟��� 7�I�0�m��y��MS ������ѯ����Z� +���O�a�s������� �Ϳ߿ƿ��'�9�  �]�Dρ�hϥϷϞ� ������߄���G�Y� k�}ߏߡ�����8��� ����1�C�U��y� `������������ �-��Q�8�u���n� ���0�����) ;��_q�ߕ�� ���V�7I 0mT����� ���!//E/���� ��/�/�/�/�/�/:/ ?~/?A?S?e?w?�? �/�?�?�?�?�?OO  O=O$OaOHO�O�O~O �O�O�O�Od/v/'_9_ K_]_o_�_�O�_?�_ �_�_�_o#o5o�_Yo @o}odo�o�o�o�o�o �o�o1UgN ��O_����	� �n?�Q��_u����� ����Ϗ6��ڏ�)� �M�4�q���j����� ˟ݟğ��%���}�6�o���������ɯ)]��a�ݯ�,� >�P�b�t�ۯ����� �����ٿ���:�L� 3�p�WϔϦύ���Z���s�{�$UI_P�OSTYPE  ��u� �	 ��-���QU�ICKMEN  ���0���RE�STORE 1~��u  '���a��ߴ���a�m������1� C���g�y����R� ������	����(�:� L������������r� ��);M��q ����d���� \%7I[m� ����|�/!/ 3/E/��d/v/��/ �/�/�/�/?�//?A? S?e?w??�?�?�?�? �?�/�?OO�?OOaO sO�O�O:O�O�O�O�O __�O9_K_]_o_�_�;�SCREK�?�P�u1sc���u2�T3�T4��T5�T6�T7�T8ܼQ�STAT�� �_Ӵu��USERx�P�_�RTPSC�SSks�SWd4Wd5Wd�6Wd7Wd8Wa��N�DO_CFG ��F�E���OP_CRM5  A���f��PD�Q9i�None>��0`_INFO 2Հ�up]�0% �_Z�
K.o� d���������5�G�*�k�4��aO�FFSET ��qx�"S��*_�� Ώ�����(�U�L� ^���b��������ܟ ���$�6���`߂�p���
��ʯV�a�aWORK ��m�������z�/`U�FRAME�o�R�TOL_ABRT8i��c��ENB��{�?GRP 1���\�Cz  A�� ޱ"Q޿���&�8�!B�T�y�J�U���a~��MSK  ���q��Nf�%�i��%R��ϛ�_EVNĉ����f֑b3�
 h�aU�EV��!td:�\event_u�ser\��M�C7�Rߧ��`F׭F�SP�K�P�spotw�eld��!C6 �߈ߚ߾P��!��a� �T��ו��C�1�� ��g�y��������� ��^�	���-�?�u��� ����������6%Z �;��q�@�� ��
"�W�33�:i��8�� r����/ �'/9//]/o/J/�/ �/�/�/�/�/�/?�/�5?G?"?X?}?�?�$�VALD_CPC� 2��� 8k?�?�a O��Q�<�*�O7OIO��"S&BdpJm@j��IlD[ �OV�?�O�?�?_O /_A_S_bOtO�O�O�_ �O�_�O�O(_oo=o Oo^_p_�_�_�_�_�o �o�_ o$o9K�o lo~o�o�o]�o��o �o� �G�Y�hz ����׏b��
� �.�C�U�d�v����� ����Џ����*� +�Q�c�r��������� ̟����)�8�M� _�n���������˿گ ����%�4�I�[�m� |�����Fϴ�ֿ���� ��3�B�W�i�xϊ� �Ϯ����������� /�>�S�e�w�ߘߪ� �߾�������L�=� ,�a�s�������� �����$�9H�] o����������� � �D6k} �������� .C/Rg/y/�� ����/�	?/*/ ?N/O?u?�?�/�/�/ �/�?�/O?&?8?MO \?qO�O�?�?�?�?�? �O�?_"O4OI_XOm_ _�_�O�O�Oj_�_�O o_0_B_Wof_{o�o �_�_�_�_�_�oo ,o>oSbow���o �o�o�o��(: pa�P�������� �� ��'�6�H�]� l�����*���Ə؏� ���#�2�D���h�Z� ������ԟ����
� ���@�R�g�v����� ����Я���	��-� <�N�5�r�sϙϫϺ� ̿޿����)�8�J� \�q߀ϕߧ߶����� �����"�7�F�X�m� |ߑ��������ߎ� ���3�B�T�f�{��� ������������� ,�AP�b�w���� �������(= L^��t��� �� $&/K/Z l�/��/�/N/�� �/�/2/G?V/h/"? �/~?�?�?�/�/�/?�?.;�$VARS�_CONFIG ��i0PA�  FP53��4LCMR_GR�P 2�PK��8�1	a0\@  %�1: SC13?0EF2 *�O�@�54�.5i0��8�0��5`0`1?�  �A@�@p
@�.N &OX_.8<_�N_{_�Av_�_UA)��@�Q�52�_�_�52 B��� �Q51�U�_ og_Doo hoSo�owo�o�o�o�o =o�oRov��<DIA_WOR�K �PE�p<z0�6,		j1PE|��wG�P ��p�Y9�qRTSYNC�SET  PI��PA�WINURLg ?�b0���X�j�|��������vSIONTMOU��53<� �ʅ_�CFG �S����S۵P~Z@ FR:\̃�\DATA\�� ��� UD1��LOG�  �1�EX=�51' B@ ����P�=?��P���ş.7� � n6  ���.6|��<����A  =�����54�Q�TRAI�Nf���&� 
�7!p��v�]4#��:|B�PK (?qg� ��7y����ӯ���-� �Q�?�Y�c�u�����\��Ĉ_GE�PK7�``0�
z0x2,�c�RE���PE�.8HLEX�PLa0�1-e��VMPH?ASE  PE�3��P=CRTD_F�ILTER 2�.PK ��E�_�� ������,�>�P�b� t�.7�Ϣߴ����������� �2�D�7ISH�IFTMENU {1�PK
 <k<1%����݂����� ����������K�"� 4�Z���j�|������������	LIVE�/SNA`C%v�sflive��+̃ �U`@4menuJO������r`��5�Y�M�O�Q��@@@Z�D��.�51<Y���P�$WAITDINEND׈`1�>HOK  �Ic�Պ~S�eTIM.ׅ���GO� q+�����cRELE|�'�Hxҏ�J_ACT' �(�qc_� ���y�%�?9F�"R�DIS`@�.�$�XVR��Q���$ZABC{B1�N+ ,Y�Bu2?�2M!� VSPT ��Q͚E�
�
��?�
�?O�7�DCSCHG ���{�@�04GBph0I-P$�+A�O��O�O�:MPCF_OG 1��IA�0��X�7_�OMPn3��I��p���?o_=���  3~�� �w�?�?��vԿ�P�R����~�lD&�t����D�)��?^U���=��Q�w@t_�_ �_�_�_�_�_#`d2u�Vo<o^_�o�ei´� ²E�³#��o�h�h�`�o �o&P{�_�_o� b0&o8od4�@�����O�t_CYLINuD����K �}f ,(  *��&���O�6�s�Z� �o����͎���_� ����J���n����� Տ��Q�7��ӟ��� e�F�X��|����G�! �_�����3�o�ܯǯ �婓�0�姖�J�A��tSPHE_RE 2��}̪� ����������(�;� �(Ϥ�L��ѿ��i� �ύ�������5�G�$� ��H�/�A�~��Ϣߴ�l��h0ZZ�& ��