��   ��A��*SYST�EM*��V9.4�0107 7/�23/2021 A 
  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41p� d =R��&�J_  4 �$(F3IDX���_ICIfM_IX_BG-y�
_NAMc M3ODc_USd��IFY_TI� ��MKR-  $LINc �  "_SI�Zc�� �. �h $USE_FLC 3!�:&iF*SIMA7#QC#zQBn'SCAN�[AX�+IN�*I���_COUNrRO�( ��!_TMR_cVA�g#h >�ia �'` ��p��1�+WAR�K$�H�!�#N33CH�PE�$O�!PR�'Ioq7i�OqfOoATH�- P $E�NABL+��0BTf�$$C�LASS  ����A��5��5��0VERS�G�  XKAIRTU� O@�'/ @E5��������-@{FA@A�E��%A�O����O�O����QEI2\K �O;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo�O)�W?"Hg@ ����j@�o�o�i�ܧ � 2\I � 4%Xo�� }A�A�o;_qP ������@�A� ���8��)�n�M��A@�c$"+ �k�K-@b��ń�AЄX}A @A-@�N��
��.�@� R�d�v���������П ���F�A偍A��(� :�L�^�p���������`ʯܯ�DxLsWn� 2�l� O�a�s���������Ϳ ߿���'��A�Z� l�~ϐϢϴ������� ��� �2�=�V�h�z� �ߞ߰���������
� �.�@�K�d�v��� �����������*� <�G�Y�r��������� ������&8J U�n������ ��"4FXc |������� //0/B/T/_q�/ �/�/�/�/�/�/?? ,?>?P?b?ah�4�0�� �?�p