��   g�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����BIN_CF�G_TX 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG���DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST��NSS�* 8�D�FACE_NUM? �$DBG_LE�VEL�OM_N�AM� !� FTޒ @� LOsG_8	,CMO>�$DNLD_F�ILTER�SUBDIRCAPCp��8 . 4� �H{ADDRT�YP�H NGT1H����z +�LSq D $ROBOTIG ��PEER�� MwASK�MRU~;OMGDEV���PINFO. �  $$$�TI &�R�CM+T �A$( /�QSI�Z�!S� TAT�US_%$MAI�LSERV $�PLAN� <$�LIN<$CLyU��<$TO�oP$CC�&FR�&�YJEC|!Z%E�NB � ALA5R:!B�TP,�#�,V8 S��$VkAR�)M�ON�&����&APPL�&P�A� �%��'POR��Y#_�!�"ALE�RT�&i2URL �}Z3ATTA�C��0ERR_T7HROU3US�9H!��8� CH- c%�4M�AX?WS_|1;��1MOD��1AI�  �1o (�1�PWD  � LAط�0�ND�1TR=YFDELA-C�0<G'AERSI��1vQ'ROBICLK_HqM 0Q'� XML+ �3SGFRMU3T̑ !OUU3 G_�-COP1�F33�A�Q'C[2�%�B_AU��� 9 R�!UP=Db&PCOU{!�C�FO 3 
�$V*W�@c%AC�C_HYQSNA�U�MMY1oW2?���RDM* ? $DIS��{SM	 l5�o!�"%Q7�IZP��%� �VR�0�UP�� _DLVSPA}R�  �SN,
3 �_�R!�_WI�CTZ_I�NDE�3^`OFF,� ~URmiD�)c��   t 9Z!`MON��c�D��bHOUU#E�%A�f�a�f�a�fLOsCA� #$NS0oH_HE���@�I�/  d8`A�RPH&�_IPFF�W_* O�F``�QFAsD90�VHcO_� 5R42PSWq�?�TEL� �P���90W�ORAXQE� L�V�[R2�IC�E��p� �$cs ? ����q��%
��
�p�PS�A�wo# XK	�Iz0AL��' V�
���F�����!�p�i��$� 2Q�$a����� ���� Q���!�q�����$� _FLT�R  �\� *����������d$Q�2��7rSH`�D 1Q� P㏙�f���ş��� ���П1���=��f� ��N���r�ӯ������ �ޯ�Q��u�8��� \�������󿶿�ڿ ;���_�"�XϕτϹ� |��Ϡ�������6� [���Bߣ�f��ߊ� �߮���!���E��i� ,��P�b������� ���/���(�e�T����L�����z _LUA1}�x!1.��0��p���1��p��255.0��r�	�n���2����d %7I[3e���  ����[4���@T'9[5U����{���[6 ���D �//)/s���QȁMA���MA�P������ Q�	 ��u.<�/?&?�/�J?\?n?A?�?�?m�P �?�?�?�?�?O.O@O@ROOvO�O�Ou.kO�l�q��O�L
ZD�T Status�ZO�O5_G_Y_n�}�iRConnec�t: irc{T/?/alert^�_ �_�_�_mW#_oo,oP>oPobot�^�P~2g���go�o�o�o�o �o�o	-?Qc�ul�$$c962�b37a-1ac�0-eb2a-f�1c7-8c6e�b56401a8  (�_�_��H�"�p�1!W��(��"S��JE�� X��C� ��,$���W��� ��ˏ���֏��%�� I�0�m��f�����ǟ��������!��u��R����� DM_�!����SMT�P_CTRL 	����%����D F���ۯt�ʯ��'�d�Lz�N�� 
j���y�q�u�����Ԙ��#L�UST�OM j���̜��  ���$TCWPIPd�j��HX�%�"�EL����z�!���H!T�b�<�n�rj3_�tpd7� ��i�!KCLG�L�i�|��5�!CRT�������"u�!C�ONS��M�[�i?b_smon����