��  
��A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1zTU4QRP�ARx1�R� � $TIT91� ��� ��Td�T0�ThP�T5��V6�V7�V8�V9�W0�W�WOQ�U�WgQT�U�W1�W1�W1�W�1�W2�R�SBN�_CF�!@�$<!J� ; ;2�1_�CMNT�$F�LAGS]�CH�EK"$�b_OP�TJB � ELLS�ETUP  �`@HO8@9 PR�1%�c#�aREP	R�hu0D+�@��bl{uHM9 MN�yB;16 UTOBJ �U�0 �49DEVIC�ST	I/@�� �@b3�r4pB�d�"VAL�#ISP_UNI��tp_DOcv7�yFR_F�@|%u13�x�A0s�C_WA�t�,q�zOFF_T@N.�DEL�Lw0dq8�1�Vr?^q�F#S?�o`Q"U�t#�*�QTB�����MO� �E �� [M�����R;EV�BIL����XI� v�R � !D�`��/$NOc`M�|���ɂ/#ǆ� �ԅ���1X�@Ded� p E RD_�E��h�$FSS�B6�`KBD_S�E�uAG� G�2BQ"_��2b�� V!��k5p`(��C 0q_E�D� � � �t2�$!S�p-D%$$� �#�B�ʀ�_OK1��0] P_�C� ʑ0t��U �`LACI�!�a�Y�<� �qCOMM� # $D
� ��@����J_\R��IGALL;OW� (Ku2:-B�@VAR���!�A��BL�@� �� ,K�q���`S�p�@M_O]˥���CCFS_U	T��0 "�A�Cp'���+pXG��b�0 =4� IMCM ��#�S�p�9���i �_D�"t�b��M�1� h$�IMPEE_F�s��s��0� t����D_���J��D��F��%�q_����0 T@L��L�DI�s@G�^� �P��$I�'�����CFed X@G�RU@��Mb�NF�LI�\Ì@UIR�E�i42� SWIYTn$`0_N�`S 2�CF�0M� 	�#u�D��!��v`(����`J�tV��[ �E��.p�`�ʗELBOF� �շ �p`0���3����� F�2T��A`�rq1�J1��z _To!@��p��g���G�� �r0WARNM�p#tC�v`�ç` �� COR-UrF�LTR��TRAT�9 T%p� $AC�CVq��� ��r$�ORI�_&�RT���S<���HG�0I����TW��A�I�'�T��1D���� �202�a1��HSDR�2��2�2J; �S���3��4��5���6��7��8��9�KD׀
 �2 @.� TRQ�$vf��4'�1�<�_U<�G�����COec  <� P�b�t�53>B^_�LLEC��!~�MULTI�4�"u��Q;2�CHILD���;1���@T� "'�STY92	r��=��)2�������ec# |r056$J ђ��`���u�TO���E^	EX�Tt����2��2�2"y����$`@`D	�`&��p���� ��(p�"��`%�ak�� ���s�����&'�E��Au��Mw�9 �%� ��TR�� ' L@U#9 ��z�At�$JOB�����P��}IG��( dp������^'�#j�~�L�pOR��) t$�FL��
RNG%Q@�TBAΰ �v&r�*`1t(@��0 �x!�0�+P�pX�%���*��͐�U��q�!�;2J�_)R��>�C<J�8*&<J D`5CF9��`�x"�@?��P_p��7p+ \@RO0"pF�0��IT�s�0NOM��>Ҹ4s�2��� @U<PPgў�P�8,|Pn��0�P�9�͗ RA���l�8?C�� �
$TͰt�MD3�0T��pU(�`�΀+AHlr>�T1�JE�1\�J����PQ��\Q��hQCYN�T�P��PDBGDd̰�0-���PU6$`$Po�|�u�AX�܆��TAI�sBUqF,��E�1. ���l�F�`PI|�-@PvWMuXM�Y�@�V�FvWSIMQST}O�q$KEE�SPA��  ?B�B>C�B�z�P��/�`��M�ARG�u2�FAyCq�>�SLEW*1�!0����
� �1M�CW$0'���pJqB�Ї�qDECj��exs�V%1 �Ħ�CHNR�MP�s�$G_@�gD�_x�@s��1_FP�5�@TC�fFӓC�Й���qC��+�VK�*��"�*�JRx���SEG�FR$`IOh!�0S�TN�LIN>�csPIVZ��1_�A�D2�� ��r 2��hr�r�A��?3` +^?�� �եq�`��q|`����p�t��|aSIZ#�!� �T�_@%�I��qRS�*s��2y {�Ip{�pTpLF�@��`��CRC����CCTѲ�Ipڈ�a���b��MIN��a1�T����D<iC �C/����!uc�OP4�n j�E�Vj���F��_!uF��N����|a��=h?KeNLA�C2�AOVSCA�@A�(�R�@�4�  c�SF�$�;�Ir P�4�@�05��	D -Oo%g��,,m�����ޟ��BRC�6� n���sυ�Uz��R�0HANC���$LG��ɑDQ$ft�NDɖ��AR۰�N��aqg��ѫ�X�M�E��^�Y�[PS�RAg�X�AZ�П���rEOB�FCT��A��`��2t!Sh`0ADI��O��y�s"y�n!�� �����~#C�G3t!N��BMPmt@�Y�3�afAES$������W_;�BAS#X�YZWPR��*��m!��	 c`R_L\
 � 7 ���C��/�(zJ�LB�$��3����5�FOsRC��_AV;�'MOM*�)�SԫBP�H�1�HB�ɀE��F���PYLOAD&$ER��t&3�2��Xrp�!�rz�R_�FD�� 8 T"`I�Y3��E�&���Ct��MS�PU�
$(kpD��7��b�9�B�	EVI��
�!e�X   $I��B@X���X<&�SY5�; �R_HOPe��: �pALARaML�2W�rxR_�0; hb P�q�`yM\qJ@$PL`AB��M����0�E���	���V��0�~qU��PM3�U��<�T[ITu�
%�!�[q�Z_;��3= ŔB pQk��6NO?_HEADE^az� �}ѯ��`􂳃���d@F�ق�t� n��>����@��uCIRTRH�`��ڈL��D�CB@64�RJ��p�[Q��ƽ�?�2>���ORĭr��OK��T`UN3_OO�Ҁ$���P�T��Ъ�I�VaC�np��DBPXWO�Y���@�$SK�ADR�DBT�T+RL��Az�րfp0bDs���6�DJj4 �_�DQ5�AP5L�qwbWA��^"WcD�Ak�A=�2>CUMMY9��C10������B��[QPR�� 
���D�����C l�Y1$�a$8�/
�L�D����7����0E������PC�1F/_cPWENEA@Tf�G=/����RECOR>"HH @��oC$L�#D$��PR���+jp��nq�_yD$�qPROSS��
���
�r� -�$T�RIG� �&PAU�S�#ltETURN��"�MR��U� �Ł� EW����SI�GNALA�QR$L�A�0O5�1E$P�D�F$Pİ�AG�c0�A�C~4�3��D�O��D��"�!&G�O_AWAY�"M�OZq�Z�CS�G�CSCBg�I qԻa#�<�ERIL0�Nn�T�`$�������3�2L�@	BGAG~@R�P���44BD�/ACD�OF�qF� YF�'C�CMA� X'C��$FRCINI_��5#Ӑ@��$NE��@�F�4L��� J� ���<����R�/���P\ OVR�10���$Ҡ�$�ESC_�`uDSBIOX��(Te���VIB�� `szLZp��LV��pSSW��L����VLP�:�Lk� ZX���ѣ�QP���USC�P��A���A��MP1�U�C�P��Rt`�S5QeU����S g�Cg�Sd���dc�C��g.���AUT�O$�a҃oac�SB ����T���C/B���2�f$VOLTr�g��A� �� �1D���a���@���ORQҀr�$DH_THE� �PRp� )t&wALPAH&t��o�Jw�  p���.�R��{s�5 c`r��A��ED�S\ %F�!M�q�sV�r�v��ûvL�R�tk�����BTHR����T(`����zVɖ�L��Q�DE7 ��1K�2P�C�X�C�f�F�� #�g��QT,0Т�p� ��f�d����g�����N~��s2>�Y0IwNHB��ILT�  ɡ�T?��3��/�఩3��P)Q0Q�T)PeŖ0Y�AF5�OM�r�o� �z���o�)Pڳ|���`o�P��͘o�PL?�xx��o�TMOUXc |��o�� w�+��1H�H��A��g�Io������DI~���'�S#TI�󍣣�O��� Hҽ�ANǥ�Q`�S8��b͑�h$kЈ����/�_Ig�yPR	AOP�P.C��kӦGMCNQe�E�L�VERSe��bP'PI/�F{������-G�DN��G����Bo�F�2��ӷo�MԺ��F��_ԴM�D ��䧭�ed��3�ea���DO� ��U��2�j�ʹDI��e�۴��� �������/�F0�����ON���ȅQI�VALȤCR�_�SIZJ���A&�REQ�R���2���D�CH)���ʹ��z�`D��ō��&�S_��>X��/WFLG�����/U$CV�iM8�@VQ��FLX��"`�B��-䯤��ALJP��C��� �bT^�W�^� gRxc� cQ�NGDMS�m�K�C�{P_M�  �STW`.������h�AL�P Y�YQk����V��e�IAG�'�d7��J�T�A�P� R� �A^��]� `]�	`]�6[�q_D��g��c ����YP����r�"8=Tc� ?����@�1��T�ۡ���LH�?��! �0��LDĀ��U0JFRI�0 �P��I\15�jIV1U�s1IUP�PZ�Q��C�LW���
�P�L�C��S��CWC �	/�� �IZ!Fů��T�Q�g��?���g���~�
�P�5R�SMI�T��0  bb *�sd2AWda�_T
p5��0NS_PEA��;����ܢSAV�����7%8I��CAR؀�P0�!<$f�E"CR������T[#El@I�\"STD;�[!F�`'�x'�QOF7�k%B�"RCO҇&RC��v(����1�R�'=�G%��WMEA�Q_naI��AQ��(�a$2F�-4I�*7�I>R99/Q97��k8M��H!C�`Rp  �tp�2F��SDNXX�Va��  �G2�AK P $M!� �s�S�17��3nc%j9�f��4[�RA�D�0CY_ L L!IG10'1BV�1@�07H2�NOà���޻CDEVIP �M�0$�RBT��FSPc3�C-T�DB�Y4�A�G3�3HNwDGD�1N H�0�GRP�HE�!XL�<Uj�SDF02��4L�` O�Bp��U�sFBQ\�FEN�@��uSV��3 �1P �d�@DO���PMCS�?P��?PuRN�HOTSW24�DpELE�1�U0\�P�RQ T�@I�[r@ � f�o`OL�GHA8F#��c:�4й3�A��0R � $M{DLb 2Q��EXȃqn6�q� �i�c�e�cJ]�	�e���#��n�d�g]PTOa�ت tb���3SL�AV� S  n�INP���F��By��1_��ENU�1T; $
�PC_eq�2� �RLvw�0�2bpS{HO�� U ���A�a�q�2rr�v�u��v�^rCF\ ?V` ,�xr�OG�W�p�%�q ��Yp�rI��!�M�AX��q0 AY�vW�A (�NTV���rV�E�0�uSKIg�T��`�}�2S���JsX!��C��s��f���_SV��`XCL�UL� �p�ONLdB�߃Y�T��OT�U�HI_V�!��AP7PLY��HI�P�v��_ML�� $VRFY�����=M3IOC_�Z�" 1��l���O�@��LS/"@$DUMMY4x𛐒�_C= L_TPJ�T�8#Cc�1CNF�Օ@_E��j@�1���D#�Q_������PCP�B���R S��k�����u �� W ���� RT_�@`�[uNOC�R X;r��TEL������rzDG��x`Y D���P_BA`L#c��!�ȥ_Ѐ�ҬHУ6Tb�E�� �Znp�R�SAR�GI�!$���`Y�n�SGN�1[ �8�`ЎIGNQ�G�,J����VJ�d�>[�ANNUN��ޕ���_E�'wATCH������Ķ���u\ <�0�@����S$ah�����������1EF I�� �] @�0F��I}T�	$TOT! @�C�����-�M�@NIva^,B�����A�q��DAY�3LOAD�D�&������ �EFV��XI@R_\���I�O���a �AD�J_R_!x``���� 2�"�������`_��PI�cѝD���AG����1a �0��\�=� \��䇡��U! ���CTsRLN p b;��TRA��#IDLE_PW��G�XԮQ���V�GV_WЉ`a� �'��Ax`c�� 1$k��P�STAC�#M��Q���R2 A�e����SW��A�����Չ``f�OHα(OPP��#IR9O� �"BRK�Ө#AB��o�㾢��@�  ��F�Չ`b��x�"@�RQDW��MS��6X�'2�?IFECALƳ� 10tND��M���`B��� ���CP¢ʱN� Y���FL�A#��OV Y�H�EO��"SUPPOd���gL�p��Q�R�"Xт��Y��Z��W�����P����Bт�XZbq�$Y2@C	O@P�S��2
報`�bD!���"��*pyI�0�sd `�@/CACH�5�Vc�S��+0LA SU7FFI���p7�Yq���6���RM�SW�e 8vK�EYIMAG�TM@S��&�""@r|�27QOCVIEN��6�f ^aBGL[�F��?����0R�j�g���PST��!�b�������x����EMAI�`�N��E���FAUD� 7�h^�Yq��Z�U�3)qq 5�i�< $#�US�Wи�ITߓBUF�����DN��H�SUB-$�DC���"��p"SAVx%:"#�@_q�X��'󀤶P$N�UORDO�P_- �^%=��(OTT��_�P���0LM$��$g�F�'AX�3.�U�X- ����#_GD�
z@Y�N_��7�j�D��E��M����Tʬ�FQ�a��DI.BEDT�0Ch�6�Ik;r�GN!�&E�D$`���QvP��FP� l (�pSV � �Tć�[����1��?m� <�n����#C_RYIK Q�#B\� D3pRE���1DSP6BP�`hIIMx#]C�A���1A�U:G��8!CM�IP\�C��~ \DCTH^ oSPB��T\��]CHS�3?CBSCi�m ��V�dVP�#�T_D*cCONV�ˁG*cT^ ZF- F�D�A�d?C�0"1R�SqC��DeCMER�T>�1FBCMP�S�0�ET�S nFMU��DU! ���6ђCDSI�@� �O �EO���oӈG�QR�Q�U=�MAS��Z-��P�T�2��P[�A�1p� �"��Q�4$ZO�0+�q�$�U��ޔ�ePM��eCN�$��l<�l�iGROU�W��2��S� �MN�ku �eu�ep
||�i�c�H�p!�ez��0CYC��shw�c��:�z�DE�_D���RO�aP��qf��gv3�O���vO��w�tU��B��u��8�p�ALA �1q��1z�Г0��PB��J�QR�T7��Rr ,�0>��%�>�G1LR1q �
H0��NOՑ�1s �����Ų���Pv���EC����U�A�I����0V`tH *��L���	��V° ��12�b�2���2����2���2��2�7/�8B/�9/�D�1�;�1H�U1U�1b�1o�1|�U1��1��1��2���2;�H�2U�2b�2�o�2|�2��2��2*��3��3;�3H�U�U3b�3o�3|�3���3��3��4���2X	T�ѡ1u��\0xf�\0�Ug0}�@eK�F{DR��vT VE���!G�RG��RE��FG�SOV�M6C�A�TRO�V�DT� 
�MX��IN깅�	���IND(�*�
Tȑ0E0Z0G-1����PM�3�9D��RIV�Pyb�SGEAR6AIO*�KڲQN�0��1��(��P�0�aSZ_M�CM8 G񨰰�UR�Rw���P!?� ��]p?&�C�?&�E
�.��:!\�P��x ��Pq���RI���;"E�TUP2_ y b�9#TD�@
�7%�T�`>є׎�Fռ�C�Q2z T�:"�4)��:%�PBW�(�I+FIf�W M������PTP�FLU=I�{ иqd UR��!��B�18P0 �sEMP�pC2u$b�S�?xn�qJ��� �#VRT^���0x$SHOc�L)��ASSP�!s��@��BG_;�������U���b���o�FOcRC�T �Qd|�KFU�1�2�2�1p�� �^ (�} |d�7NAV_a�b�����ְS�yc$VgISI��ۂSC4CSELЮ�� �rV�pOg�$b�ְ�b��$r�I���@��FMR2��~ ���P{r���0 ���������������ڲ_ɡ��LIM�IT_���TC_L�MƤ϶�DGCL�F_Å�DY�LD�>т�5��yϋħ�Mԝ��SJ-	 �T�FS� �T� �Pl�	�3E0$E#X_	 	1!0YP�ba	3B5B�G�'Q��� �d��RS�Wa%ONZP�EBcUG��ߵGR�`�g@U{SBK�aO1n� C�PO ����P��Mt�O�t`SMu�E�"n�up�F�y`_E �� �0i�TE�RM%�%o�ORiI�1 �)SMp	Os� �%�S`Z(}�f&��UP�p �� -E�Fyb�b�)#� �x�yG�*� ELTO7��p�0BPFI*c�1���a�@$�$�$UFR��$���!0L�UH OT7BPT�aܻ�#3NST�pPA�T�q74PTHJ��a�PE�P�3ap�!ARTi �%� i 12�"�REL{:�1SHF�T�B�!?1m8_��R(�P�SX& c $r'�0��h����]s\1�0IԞ0eU�R �pPA�YLO�@nqDYN_#�O��R?14�Ʌ�@ERV:�
AX�8^� 7�p{2ס�eE���RCN�ɅASYM�FLTRɅ�!WJ�'^�Z�E^�i1�IX��QU�D�pAm5� YF5PFP$CFQ�6OR��pM��h!������>0� Ea s�Hs��T� �%2X���POC�!�>��$OP����rc��ֱ��jbRE�PR�#\1��q?3eH�R=5�U�X�1>��e$PWR���u�=@R_�Sb4d�t��#UD^ҧ�WQ�" ����$H��!^L`ADDRxfH!AGA2eaZaSan�R���� Hl�SSC �ף�e壒eU��eb��SE��� HSC=D��� $N�zPE_�p_��2�bPE��D�:�HTTP_���H�� (��OcBJ�pSb��$^f�LE03:`qt� G� n�Q�p�_U��T�arSKP��2�K9R�gHIT���� zP��Par��^��P��PSS����JQ�UERY_FLA��!_qB_WEBS;OC���HW���!����`�@INCPUVd�O �vq:��7��d8��d8�b���IHMI_ED] �T �7RH��?$d�FAV@ �}��b�OLN�ґ 8�l�R���0$SL�!R$INPUTM_��$�P��P��w ��SLAz ��������|C��|B�0���`F_�AS����$L��5w�ѿ1��b�!`;ࢃ���@HY|�pl�E�SQ �UOP�� `1���^f8�\�8�c����PP�3�P���Αc�ےĖo�IP_sME��m�� X1��IPZ`V�_NETV�pd�R|�+��qWDSP��p��F��BGV}`g�MgA�m�� l:�3TA4"B<pA�TIԕ�E��� ���0PS��BU ID�r�����P��
qd���10�D�v�������N	�| 
��IRCA̰�!� � �Sy6�CY�`EAT�K�@}�P�8��3h�]�RY0x�A���ADAY_w���NTVA7�Ԡ��p܂]5����SCA@��CL��w�TQ��z��m����^2�'�N_�PC�)�Ţ��n����C�\�0rw���`��� 2�W�c���m���ғ�0r��LAB11�� �ǗUNI
���C ICTY��e�^eԂR�������?�R_UR�LF��$AL��EAN�`�e�t �sTh��T_U]�ABKY9_2�2DIS�������J�m���$`ҙE��R����O �A�灋�Jh��F�L+]������Ѭ
��UJR��� �SpF3�7��'��Q����J7��O�B$J8�7`��
���7����83� �AP�HI� Q�P�D�J7J8�2i�L�_KE��  ��KZ�LM� 7� <�XR$�-��C�WATCH_V�A��'@��,vFIE�L�Pcy����� D '1V0@@���C�T���%� ��LG ��� �$=�LG_SIZ�[t�2�� 1�(�1�FD<�I0�G��>�/�  I�;�.�S7���  ��(���^�� ���A4�� _CM32

F�A..�r�T(-��29�S� S(�S^�_I Ri�S k].�RS��N0  MZ�IPDU~��LN��r����p2@�O���c�KPLn�DAU!EA�`0Z�nT7-GHoR(��4�BOO�a�g� CK��IT�s�k^`G�REk��ScCR; �sL�DIF��S� �`RGI"$D�̆?��T��t4�	SAs3�W�4�?��JGM'MNCHL�s4�FN{�&K?'�-�=)UFK(�0K(F�WDK(HL�)STPK*VK(��K(rK(�RS�)HPg+<�C�T�#�B?��`�9U �a_$�� %��T�R"G/)�0POV7�*�`�#5$W�M)EX;�TUI=%I��B�G����Ar�3#�3; ��$Sű�	ᰟ�0v�NO�6ANA4�{Q²AI4�Zt�EDCS���cQC�cQBOWHOcGS=ӁBnH9SzH�IGNG�Ű�Y�<!�k�ZDDEV6�'LLu�Y��eФ���TU$p=���(�A����B�Qdѥ���P��3�\�sPOS1IU2IU�3IQ���2R@eЦ �S{FP,D���������a�uq0��VST��R8Y$��0�P� �$E�VC �[ep�`�Vf
q�4d�� L
�Z���o�0� �SxpO��t�`id���^�_ ���W��q޳��c �MC��� ���CL�DP��s�TRQLaI��u��i�dFL\��b���c�D���g��LD�e�d�eORG�{��! r��RESE�RV;�LtG�LtR� ��c��� � 	`�e�%�d�e��PT�`ұ�	0q�t�vRCLMC�tL^�y]�D�q� MI�#�������$DEBUGMCAS]�������U��T7@��E��ޠM�FRQ��� �� "�HRS_R%U�aa^�Al�#5�FREQ8 t$<�00�OVER��Y��&��V��PT!EFI�̠%Fa_��QX�yt� \
Ќ���$U�P\�?L�pűPSHP��	��AC@�s����sU��$�?(��`IS�C�ծ d��QR5Q��	I�TB�̠c ���1��AXs��������EXCES�"�_�Mj���۠�t�s�'Qc�SC�P O� HY���_���~��������M�K Ա���%�B�_�FLICAdB��QUIRE�#MEOs�O���V�Lc`M�Ų �`z��h�a��r�aND������Q�#���D|O�INAUT��O�RSM����@N��r��3����PS�TL�� 4�L�OC�VRI���UEX��ANG-B-�qq�ODA\��p����Ю�MF�e�����Ybb�0le�� #�S�UPhe	�FX��I�GG~ � � �pbc��E�bc	6bd�� ݂�R4��PD��PS�4�0s3/�W�TI��<p�V���M~��� tV��MD��IA)��W@���q��H�����GDIA8��Ñ�W����/Q�1��D?)$�L���Ӧ��� �CUG�VОp-��
�O�_�=ѹ ���ДS������i�{�P{�� ���P�z�KE2��H-$qB: n֤�ND2�r�����2_TXkdX�TRAWC���r�M8Ԁ4q�`�P.�}X0���P�d�SB)`�U/SWCS;�Tf����V�PULS����N�S��n�
u�JOIN�� u�6`"��r=b��cb���P�r�����cb��o�TA�8�{����� �E&r�SC��PJ��
��R�PL	� ��&��LO9>л�m�&� l���Bҍ����|aMRR2g��O 1}�A�q/ d$G�I����GEA��2���p ;EPRINE��w<$R��SW0�t��sABCŸD_�J��z�-���_J3:D
>1SP���-�P>e3dG�8`
-��J�s�mr�q�O�AI��qCSKAP�j�3�3��J@L�Q������_AZ�r�6ELx�A��qOCMP���q���RTD�a�c1���m��P1��t�0�Z�SMG� ���tJG�`SCL<ɐ��SPH_�@L����-���RT�ER ����A_D@�!ڰA�@�SL��$DIL�23U��DFԐ5!LWn;(VEL�aINwb�0^ _BLW@-�f$ ��qV$k'�'|%�s΢ ECHR�tTS�A_Ԑ���E5`���B��%�BS��!:5`_S� ��%�"&%TR�%��9,'�L�DHɐ��=��8P$V�����1�$�������$��A�`R5�>��H �$BEL.�|m��_ACCEl!��7�q�0IRC_4 ��?pNT��SO$PSɐ�bLԐ ��5�c���63�F@�6 �ѩ9G�3G3�2S�̑_FQs2P@VA��7�n�1_MG|�DDsA"��FW�`Q�3�Eؿ3�2�HDE�KPP�ABN�7�SPEEfBJQ�O�`�JQ����1�!$USE_tG��PP#�CTRT�Y�@�0�q �YN�f�A=V� ��=QM9�M�o�m@OX AjTINC'Ԓ��B�D��8�W��ENCF���-��1�2���0INP�O	�I�2�U���N�TV#}%NT23_9"��cLOJ ��`��Iנ�!f? �#���g`�U"�C� �VMOSIxA;�Z�VA���L�PERCH  >c��� �g���ck� $b�tk�\T'U-@U@�A�2�eLT�6����U�$jv:fTRK�сAY���c� Oq�2^uSs��g��R��MOM)ҍ��M!P���C��jsAC�R��DU��KBS_�BCKLSH_C �2�u9�_f��ES,� ��R
�TQ�CLAL�M�Tl�p%0<�CH�K� ����GLRTYo����T���Q��NTd_UM���C��p�A����@LMTa �_Lq0O����ˇE ō�؋Ā�5��8v `�qYQ�`'��hPC�a��hH���wE��CMqC�Ձ@�GCN_��1N�ӆ��SF�1�iV'R���W�[��bʕn_�CAT��SH� ��D�V��q�V~��1�~����PA���R_	P��ys_� �Vv���fsx�i�JGŰT��v��y�z�TOR�QUPgRcoy�@O�UW�jb{�@ݢ_W �uOt�t1��e3��k3���I�I�Ik3F���P��}@VC"�00
Q�tp�1w�u@8��v䀳JRKw���,��pDB�Ms�p�MC? DLe1�bGRV���e3��k3ܱ�H_��ڳ"@)�CO1S6�i6�LN��Y� z�`�e0[ɮ[�-��ʈ��K�׵ZT�jfܱM�Yb���B���J���T�HET0*eNK2a3k3 �_3c�CB%�kCB_3C��AS{ �I�-�X�e3X�%�SB8e3v�0�GTS��ACzR��A���ڔ�$DUf�w����(m%��|%Q�a_;��Q��0�3�Kv�s(R��A�A�J�(�3�3��LPH6���U�S z���Œ���Ƽ�(����R�Vc�VX�U0�{�V��V��V��V���V��V��V��H�c�|��z�������H���H��H��H��H*��OT�Oc�O	y�UO��O��O��O��UO��O��O��F��Eѡ	�ŦV�SPBALANCE_����LE��H_�S�P�!v�������PFULC�$$���*1�uUTOy_a�i�T1T2e�22NH��2�P��@�q&��2�3�qTp�O90�1�INSE9G�2CaREV�C`��QDIF9u91�l�,"1�B�OB�,�öw2Ǡ�PS��?LCHWAR�B�2ABH��u�#C`��(\Q�%��X\qP
�{&8:�F2Z� 
|"ڡܞ1�UROB��CR��b�%p�@��C�1_�d�T � x $WEIGHYPF�P$T��#{�IYQ�`IFQ�@LAG�JR)�SJR�JRBI�L05OD�pF`2S	T�02P�,�0�1(��!� �� 
�P�2<KQ�1  2�Qd6/DEBU3L@_2=��MMY9�5�qN2��4�P$DAƛa$�0v�� ]� DO_�0A�!� <� y6o%�KQ�7�BI2A0N�SH_�(`KP�f2O9� _�� %��T�P��Q��T��4�0TI�CK 34 T1�0%qC�pz@N��TC��R�pKQD"�ED"�E�0_PROMPYSE6�? $IR��IQpo��B�`RMAI�h�Q[R�E_*0�C��eq]PR�COD�~3FUQP6ID_��.U��B� G_SwUFF-� $34@Q�A�BDO�G��EC0�FGR*3D"lT �CxTD"�UD"�U��lT��4�0�� H _F�I}19�SORDfI1 � �236���RIQ�0$ZDT�5U�`f1�5�4 =*�L_NA%Az@|<b�EDEF_ILh <b�FXd�EP2�FZ4�F0�c�E�e�FISྐ Ap�D�c�CVdё"�44��!�Z2DX�r�t~3D��O� BLOCKE2�fS�O�O0�G�alRfPUMkU<b lT�clT�elT�bxRns wUgcxT�dxRX6�v�a �SO e��U<b�U�c�S�w�hX?@P �dO@��a��0WMxL�Cs��(`TE7��4��( $1LOMB�_f���02VIS���ITY2Av�O>J3A_FRIU��F SI�a��	Rw@H҇�@҇3�32W��!W��찰���_��QEAS3�R������p�Bӆ4Љ5Љ6�3ORMULA_uI2�E�THR2 �G,g�� Ч<�8�5COEFF_AO^A�Ԕ^A��G
�23S0�2CA&�?b�3$H�3'dGR�� � � $hCp�BXN@TM6w�N�CudBKsh�CER��T,t+d�0�  �NLL�TpS6�_�SVt����p��0ȸ�����0� @�SwETU�cMEA�@�KPi�0f1�R� � g�  ��  �0���'�$�'�q2�AbHz@q7qt����Rb��Ap�apn�t�� PREC�Q:,�9ASK_� 4��� P�!1_USER�"��3 �����VELe���3 ��ܵD!I`��M�T?ACFG��� � |@�Oj"N�ORE� $@'��S�I�!��w6M"UX��P�A�DE�� $KEY_�3}�$JOGu��SV����Ñ!Y�5�SWj"�aaӍ�T4�GIY� 4 �?� 4  �e'2k!XYZ�S����3k  ��_ERR���� � ��=AP��Є1��{�$BkUFf�XX� T�wMOR4�� H� CU�$Ak!j��Aax����Q$� r��aW�	 ����G6�� � �$SI��Y�İVOxY���OBJE�Z�ADJU�2\�EGLAY`��%��D
�OU�P��j�JQ�R=i�T�9��8��2DIR=�E����� DYN��"��	TY�"R��O@I0�"�OPWORK����,�0SYSB9U1�Y�SOP��?�$����U���PCp���PAð,���f"Y�+OP�PU!��!zM�$�IMAG/�1� 1�Z2IMz�M��IN��J�RGO�VRDv���İ'�P )�I� ���s��k"�LApBЗ�'�PMGC_E`?ѭ1N1 M��1�21�2d0v��SL��� � ?$OVSL��cň�a�`c�2j"��_ v�#�Pw�#�P-B=�2bC� >`��q�?w�_ZER7���Z�$Gd�ю����� @����%MO6PRI\�� 
��P�	����PL����  $FWREE�E����T���L���e�Tg �^0ATUS��TRGC_Ta�N�MBR� W@+��c�1,`���� D�1%�fÌ�L����"���QJ ����X�EQ3������� � PUPa��`�aCPX�@w"�43��^��PG�ڻ�$SUB?�%�q�?�JMPWAI�T�2W%LO��F<eA�RCVF�A}@�R"Z!RV�R"AC�Ct R��pB�'IG�NR_PL�DB�TB^0P�aS!BW�P�$/�U1@�%IG��@I��TNLND�&�"R��<r�N�@���PEED�HADOW^0��/����EK4")!W`SP]D0!� L<A2�pX`k0��y3UNI*��{w0�R�|LY�`� IS�PH_�PK����RETRIE�3�)���0v�@FI��� ��P��0�4 2��D�BGLV�#LOGgSIZ]��aKTw!�U��0DD�#� _T���M��C��R�V@�?MRPC5���CHE3CK� ���P�0!%�#��9a�L#Y�NPA*pT�2����@P1 � h $AR#B!R���S�a��O�P��ATT���"��#FV@2��aS�3UX��B��PLI�"0!� $<���ITCHR"�-W��AS�'aQS�LLB0!�� /$BA��DsY��BAM� f�Y�F�PJ5u�	��R6�V>zQ_KNOW�C�Rv�Ud�AD�X�v0�DðiPAYLOA,��p#c_O�,g��,gZ)cL�q��L=_�� !�ebP�Q��rd���fF�iAC��`j+�cd��I`h!R��`g;�|dB>��љJQ��a_Jja۱��AND:�|�tjb�~a)�PL� AL_ �^Pv0���QT��Ce�D(cEd���J3p1v� T�@PDCK��>���>�_ALPHAs�s�BE��z�AS|����!�� � �\�"oD_1)j2SdD�AR���u�� ���TIA4/�5:/�6e�MOM|�;��[�H�[�U��Bn A�D;��H��U�PUB��R`���H���U� ���1p��1 �ف2a� �2RQ����� e$PI ��1�s̱.g$�kHi*$�I0�I>�IL�� }�!}�!��}rpr�b��/3HIGmS /3o%h4Ɩh4o%� V��Ɩ��՘�!䙥!o%SAMP�o�8�Ɨ9�8o%�Ps ��h� �� ��w� ��h0�p �� ������8���-p2U�H 0��INǬ-p �Ψ�Ťo"Ъ�礼�0�GAMM��SSԨ ET��K����D�t��
$4pIB�R�2I�$HIB��_f�O�����E��b��A��ϰ��LW�� ��Ϲ����r��0:jqC�%CHK��� o v~I_� ����,r�x,q��z�s����y�1s �$cx 1��I�� RCH_D�!Ɣ RN3��#��LE@Uࡒ���x���0�MSWFL�$ہS;CR(100;�,@v�37B[֝��`;���xo�h0~�PI3A�METHOB���%V��AX �X20���2ERI��8�3�d�R�0�e	��pFHU�9�}�⌣��&�L��9�;�OOP�}���Qጡ��APP�3F��@U�v�a�&��RT��0�Oph0�.ŧ��턱 1��#��k ��L���RA��@MG$�B �S�V��P�CU9RA��GRO50��S_SA�Q��3��NO�pC���t3� ���4oFoR�����x���R���� �DOg1A ��bAw�qڪ����Aϗ��A��1-��ic�VM��� � �YQL"��a����S�b4�7B�I���a�Ô��a_��CѣM_Wb��A���=�M� ��`�0q|$AJ�R1I�"�PM$��� �A{ ��YWC�$��L1Q VaC�tA�tA�tAUt� ͰN�P��dS��J-pX�0O�s,qZ���Py �� ���M��x�u���������`2������@�qPL�q_XR� |tq�3� [��&H��&U�3�4��' �&N�sQ}�KP�Rq"
��KPW`q$P�A�PMON_QU=�� � 8�@QCsOU���@QTH]�sHO|80HYSP3ES�R80UE#0)��@OVT�  �0P�!��T�RUN_T�O��@O���� P`�5C�|A��INDE��ROG�RA� HP� 2A�N�E_NO�4�5ITx��0e0INFO�1�� `Q�:�1��sCH�1�2� (��SLEQ�� A�� @��6�e0S_EDI�T�1� �P�K�ށ����E��NU�pGjHAUTO�mECOPYށ���L��[��M��N�@�KK�PRkUT� �BNF�0UlR$G�2�D�"�RGADJ�1� -htpX_� I���(#V�#VW!XP!X��#VϓP��Np_C�YCo>RGN�S_h3�q 	�L�GOXã�NYQ_/FREQÂW֠:�N�QSIZB��L^`�r�P!QV�֠��CR1E����Y�IF>��3�NAA�%�T_G>��STATUt ��w7MAIL?��q=a<�34LAST=a�qކTELEM�Q� ��qNABot�EASI|a1l�� XЀkb��<�f�ҳ���I �0�īR4Q;1� ��b�ABS1SpE�0ӐV_a�fBAS]r�e���āU񐳐H�$,qwRM�R�c�� ��:s�𐠲Xat	0��T��| 	�b 2� ���� �v(r�w]r ���(r8�w� �DOU�3��^p��$$CX`S0O����c�c�3 �pY�SI9��w�XK��IRTU����A�� _WRK 2 �@� 0  �5��w���t��� ���	ɀ��ݏc�A��ˏ�����,�8��ȁ>�s�����Q�BS�SA� 1"�� <a�ҟ� ����,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D� V�h�zߌߞ߰�������ߝ�CC�@XLM�T0�����  �d��IN����P.�`EXE'�S�6��^0-r ��@�Q�DVʗ�Svp@�S�%�select_macro�߫��|�IOCNV�cV	� ��P��Up�(㲗��0V 1.^�P $N���H�B�E�A�?���� h� z��������������� 
.@Rdv� ������ *<N`r��� ����//&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6H Zl~����� ��� �2�D�V�h� z�������ԏ��� 
��.�@�R�d�v��� ������П������*�<�N���LARM�RECOV ����6�!�LMDG� 1�<���~��_IF 1���d  YST-�324 Over� Payload� change �distance� P) d ou�t tion f?or BWD��7� ?��S�e�w�������?, 
 ��ҿ�M�>IPL_FA�NUC_SMPL�G>  LINE� 0 �AUTO� ABORTED���JOINT 100 %׿:�!��$�RP_CL�O�@��k�E�S�BN-060 I�nvalid a�ttribute� syntax data����������NGTOL  �j� 	 A �  1�C���PPI�NFO ��� ��v߈ߚ߬��  �����ߕ���� ��)��%�_�I��m����O�������� 	��-�?�Q�c�u����������PPLI�CATION ?}������LR Ha�ndlingTo�ol� 
V9.40P/17B�~��
8834��F0F3170�2 
'7D�F5 ���Non}e��FRA��� 6c��_A�CTIVi�]�  ���*�  ��M�ODi���(��CHGAPONL{ +OUPL��;1	ة� hl�~��CUREQw 1
ث  T���	���� $�����//'/�9/�/]/��Κ� �$H��k�*HTTHSKY�/���$\~/ �/>??r/,?J?P?b? t?�?�?�?�?�?�?:O OO(OFOLO^OpO�O �O�O�O�O�O6_ __ $_B_H_Z_l_~_�_�_ �_�_�_2o�_o o>o DoVohozo�o�o�o�o �o.�o
:@R dv�����*� ���6�<�N�`�r� ��������̏&���� �2�8�J�\�n����� ����ȟ"�����.� 4�F�X�j�|������� į�����*�0�B� T�f�x����������L俬TO����DO_CLEAN�8�o�NM   � ����������ߠDSPDR3YRv��HI��@��q߃ߕߧ߹��� ������%�7�I��MAX��V���G�g�XV�fcf�PLUGGVW�cWPRC(�B����`�R���O��1�C�/SEGF/K�� *�ϩ�q�����������$�LAPN�a��# 1CUgy�������*TO�TAL���KUSWENUN�[ <��@鲬RGDIS�PMMC-�!1CL5�y�@@C�[OL��n�9�W_STR�ING 1'
_�M S�
�
�_ITEM1�  n��� //*/</N/`/r/�/ �/�/�/�/�/�/??�&?8?I/O �SIGNAL��
�ײ����������޼��ƭ�خ���ޮ����5���9��������� = 10�0������������۸���� ��1�2�t3�5�3ʰ���ް� t�M?H �װ��A����??=??OQO cOuO�O�O�O�O�O�R��R���O,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^opo�OWOR-���a _�o�o�o�o* <N`r����������&�P	O�e	L��k5�o� ��������ɏۏ��� �#�5�G�Y�k�}���p����şG�DEVO� �c�ݟ�)�;�M�_� q���������˯ݯ﯀��%�7�I�[�m�PALT]���on� ��ο����(�:� L�^�pςϔϦϸ���p���� ߂�GRIl� �8Ѭ��`�r߄ߖ� �ߺ���������&� 8�J�\�n����&�R]��P߶��� (�:�L�^�p������� �������� $6<H��PREG���  ��Z����� &8J\n��������N=�$�ARG_�`D ?�	���/!��  	�$N6	[C(]�C'�N7d)" SBN_CONFIG�0�/+�1�2�!|!C�II_SAVE � N4�!�#" TC�ELLSETUP� /*%  O�ME_ION=N<%?MOV_H� �/�?REP��M?*U�TOBACK� �/)�!FRwA:\n X?,n� '`�0n�8�� �;�  �20/07/�31 12:49:12ne(nO0 OMODO�<��mO�O@�O�O�O�O�On��O _._@_R_d_v__�_ �_�_�_�_�_o�_*o <oNo`oro�oo�o�o��o�o�o��� � �1_p3_\AT�BCKCTL.TM;�Sew��b;INI���5�&j3?MESSAG� �q�!7 �#�!�qODE�_D� �&�%�xOx��j3PAUS`�� !�/+ , 	�e /%d�r�,		\������� ������ڏ��� �J��4�n�X�z���7�A�TSK  G��?��m0UPDT�p�wd���XWZD_�ENB�t�*�ST�A�u/!�!!XIS>� UNT 2ǖ�!�� � 	 ���l�J�7C� ��� ]�� �n
�|������!"��
����,��Я�|��G�P �b �u�+ %M> ?A8R ��N'ȯ�)��M�+^�METV��2j��� P{��B95@�-�A�B4@���A/�yB"�v�7�>�8=�&��=�Q�<�I_=?�*��7_��SCRDCFG �1/%�1 	��%�"E��+�=� O�a�sϚ?n
Q�)� ���������߄�A� ��e�w߉ߛ߭߿�&�`�'p1GRc��%����6pNA0.+	�p4��_ED�p1��� 
 �%{-<pEDT-��0*:|����Y�$0Q-p3o�n
e"cOx6h��  ���2�);��l�*���:�@�������"�
�3�� M�*q���q����`��
�4��= ���=��,�
�5u��	���	/ Pb��
�6A/� �/���j/�//./�/R/
�7?}/Z?�/���6?�?�/�/�??
�8�?��&O��]��OmO �?�?\O�?
�9�OO�O9O`���O9_�O�O(_�O
�CR�H?�_ �_~=�_oJ_\_�_�_���K�NO_DEL�
��GE_UNU�SE��IGAL�LOW 1.��   (*S�YSTEM*4��	$SERV_GqRE{�`A�REG�e�$�c4��`NUMx�js�mPMUi`>4�LAYu�4��PMPAL|�p?uCYC10Jn�]~GpK~�sULS�U=�m_rA��cL���tBOXORI��eCUR_�p�m�PMCNV9v�p10s~%�T4D�LI%���i	*P�ROGRA�dPG_MIK~u����ALU���~���B����n$FLUI_RESUcw��o��!�MR�n�`l o,�e�w��������� џ�����+�=�O� a�s���������ͯ߯ ���'�9�K�]�o����\bLAL_OU�T �k���W?D_ABORdp�n����ITR_RT/N  T��i�?NONSTOB��� ��CCFS_UTIL .����CC_AUXA�XIS 3N� h���Ϧϸ������CE_RIA_IL�`�Кa@�FCFG N��Y�M�
�_LIMv�b2U� �P7� 	��B\��T�P
���Y�Z�U�Y������Թ�� ��Q��&$��v�X
_���"�9�PÀGP 1r�#��k�P}���`�C�`C�@�C7��J��]��p�������� C����������๪�����������ߪ�����������;L���pCk�������U����������������������� D� D�K�K�K�K� m�V?�>�HE8`�ONFI-��m�G�_P�1r� Uerŷ����������#5m�KPAU�S�q1r��  sr7}r�k��� ���9I oU����?��Aii�?�M�NFoO 1H�$Ї �]�9/T^���h>F�d9���]/�A/�� D�&t����D�)�´ ��E�³��z/4�'@�O� �*�~�!LLECT_�a!H���>��$ENU�pŕb�Ҳ!NDE�#�#H�Y�1�234567890I7R�a$�G?Y6��	H��S)�?�?�\�? �?�?�[�?�?BOOO 1O�OUOgOyO�O�O�O �O_�O�O	_b_-_?_ Q_�_u_�_�_�_�_�_��_:oo#6B�$�+� �-'2IO &29��k#Ƽo�o��o�o�gTR?�2'�nm(�؈2o ~x��(�m*z-��&_MO-RS�3)r͌a��u ]ѳy��������r:�q*r�,}�?$f�f�f���Kp���J?�P,2,�/.�e� ��Ώ������󒰊8uk)@o,�k# � ja�(�PDB.0.ʼ)dcpmidbg]������ʓ:�n��p�����Ȗ  �"n��A��X�!��럊���f�mgz�ӯ�� �f¯��| �-`ud1:@��i�+ꂑDEF Y-��c)T�cy�buf.txtt�Pu���=�/nm�Տ>����a�MMC�r20��|cdC�,$Òs212ͤ!�q��k&CzkЎ1^�A���hAӡ�A׿�B5O�����C4 y�H+C3/��C%;]C���D}�C����D�F-Ev��@F?�UE��fE�v�E�_F��n�?�����<�23nlD(�)h1��!��2�ӧ�k���
&pxc�������  D4�q��λG��  E�%q�F�� E�p͟�F-F�P� E��fF�3H ��G�M����_�>�33H��i�G�nc�G�@�G5����G�Ai��k$=L��<#�{u�`V��c:���RSMOFST �+����P_Tu1�4nmA g����MODE 5����`��3q�w!;�-�O�I�?��ߚ<�MܾTEKST��2����R�"a6�/y�uƦ� Al�k(�� b���mC�0B���CE������:d�{s +���*!�����^�T_��PR_OG %G�%ӿ�L[��`NUSER��`KEY_TBOL  G�!$"��	
�� �!"#$%&'()*+,-./R7�:;<=>?@A�BC��GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������&���͓���������������������������������耇����������������������  LCKjp�a�j STAT�\�X1_AL-�p1}�_AUTO_DO�6o�#FDR �38��2hk)U ;`/r/�/�$O/�/ H�-�k��/5����)�/ �/�/<?>O?5�\�J� N/�?�?�?�/�?!Oe� T���8ObOh3fOPO�O �OnO�O�O�O
]�?/_ A_S_�?d_�_4O�_�_ �O�_�_�_�_�_o(o ^opo_�o�o�of_�o �o�_*o,X f<z����o� �#��o4�Y�z�t� �������Ώ����� .�@��g�y���6��� ��l��ܟ�����(� 6��J�`�����V�ϯ �󯞟�)�ԟJ�D� b�d�V�����t���ȿ ��Ͼ�7�I�[��l� ��<��Ϭ�ʿ�Ͼ��� ����0�f�x�&ϟ� ����n����ߤ��� 2�4�&�`�n�D��� �������+���<� a���|�������� ������ 6H��o ��>���t��� �0>Rh ��^����/ 1/�R/L/jl/^/�/ �/|/�/�/??�?? Q?c?/t?�?D/�?�? �/�?�? OO�?"O8O nO�O.?�O�O�Ov?�O _�?"__:O<_._h_ v_L_�_�_�_�_�Oo !o3o�ODoio_�o�o �_�o�o�o�o�o�o >P�_w��Fo� �|o��
��8� F��Z�p�����fߏ ����9��Z�T� r�t�f�������؟ � �ΏG�Y�k��|� ��L�¯��ڟܯί� ��*�@�v���6��� ��ӿ~��	ϴ�*�$� B�D�6�p�~�TϒϨ� ���Ϟ��)�;��L� q�ϒߌߪϬߞ��� �߼����F�X��� ���Nߴ�������� ���@�N�$�b�x� ����n������� A��b\z�|n� ����(��O as��T�� ���//�2/H/ ~/�/>�/�/�/��/ ?�2?,?J/L?>?x? �?\?�?�?�?�?�/O 1OCO�/TOyO$?�O�O �?�O�O�O�O�O__ N_`_O�_�_�_VO�_ �_�Oo�__ooHo Vo,ojo�o�o�ov_�o �_$I�_jd �o�v����� �0��oW�i�{�&�� ��\ҏ̏��ޏ� &���:�P�����F��� џ㟎����ď:�4� R�T�F�����d����� � ���'�9�K���\� ��,������������ ��̿
� �V�h���� �ϳ�^����ϔ�
�� "�$��P�^�4�r߈� ����~���	����,� Q���r�l�ߌ�~�� �������&�8���_� q���.����d����� ������ .BX ��N������� !��B<Z\N� �l���/�// A/S/�d/�/4�/�/ ��/�/�/�/�/?(? ^?p?/�?�?�?f/�? �?�/OO*?,OOXO fO<OzO�O�O�O�?�O _#_�?4_Y_Oz_t_ �O�_�_�_�_�_�_�_ .o@o�Ogoyo�o6_�o �ol_�o�o�_�o�o( 6J`��Vo� ���o�)��oJ�D� bd�V�����t���ȏ ����7�I�[��l� ��<�����ʏ̟���� �ܟ�0�f�x�&��� ��ïn�ԯ������ 2�4�&�`�n�D����� ο࿎���+�֯<� a����|Ϛ��ώ��� �Ϭ��� �6�H���o� �ߓ�>Ϥ���t����� ����0�>��R�h� ���^��������� 1���R�L�j�l�^��� ��|�������? Qc�t�D��� ���� �"8 n�.���v� /�"//:</./h/ v/L/�/�/�/�/�? !?3?�D?i?/�?�? �/�?�?�?�?�?�?O >OPO�/wO�O�OF?�O �O|?�O�O
O_�O8_ F__Z_p_�_�_fO�_ �_o�Oo9o�OZoTo r_tofo�o�o�o�o�o  �_GYko| �Lo���o������*�@�v�\��$�CR_FDR_C�FG 9Z���q
UD�1:�w�tJƄ  �Ҁ�|��HIST� 3:Z�  ���  ?�r�@�A�B�C��p�D�E�I��g�p�o�w��h���INDT_�EN��t������T1_DO  �u��z��T2����VAR �2;���� h�'� j�f��j��r��k��k΍C��rZ��S�TOP����TRL?_DELET6�Ɣ� n�_SCRE�EN Z���_kcscy�U_��MMENU 1<~��  <�|%����tۯ�:��s �=�v�M�_������� ⿹�˿�*���`� 7�Iϖ�m�ϥ��ϵ� �������J�!�3�Y� ��i�{��ߟ߱����� ���F��/�|�S�e� ������������0� ��f�=�O�u����� ����������) b9K�o��� ����L#5 �Yk���� /��y��_MANUA�Lc���ZCD���=㙵�/%  "���rԆ
*n'
*?�|(��pd<'GR�P 2>��cB� h ���"~h �$DBCO���RIG�����"G_�ERRLOG 	?ʫ�q�/1?C?U?� �!NUMLI�Mē�!��
�!P�XWORK 1@ʫ ?�?�?�?�?�?�m�DBTB_y� CA=���!;B�l ��DB_AWA�Y�#�qGCP Γ�=�ׇ2UB_AQLs0..�"_�"Yb��������S@ 0 1B>�+ , 
�?�O0
$�O_H_M����_L@�%UONTImM������GV�I
}P�GMOT�NEN.�.&}[RECORD 2Hʫ� �_�sG�O��Q�_
+`B	oo-o ?o�XGono�_�oo�o �o�oqo�oo4�o Xj|�)�!� E���0��T�� x��������ҏA��� e����>�P�b�t�� �����+������ ��:���3�͟������ ��'�ܯǯկ���� �J�\�˯��k�y��� %�7����m�"�ϣ� X�ǿٿ�Ϡ�7ϯ��� E���i�{�0�B����� x��Ϝ������������QBTOLERE�NC^DBȧBl@L���� CSS_CCSCB 2I�,	DP
$�O
.c�� ���?�������(�@:�L��p���
+�`� ����������!3 EWi{���� ���/AS ew������ �//+/=/O/a/s/�/�/ ���/�/��Y�+:�LLE�JI��UQ4<C:A 7C��C�{0.0\��F? A�+�p+�ɴ�C�P�q1�- 	� A�k0�0B<�ߍ9?�  �6�0�?�?�(DP��qP��B���HC[�3OEO(WO��{O�(kO�O�[O�OO��K���L�d������?8;V�Oȥ[�O���OPH_#21��@��7_ �_�_�_��vPA.��_c8.�A �_o�WqQ m1�1m1!m�QB�QBo Lb)e�Yo�o�o�oQZ�P��`�`0�Dz20Ca� @��
�!X�&R[��	 5_��>7�����Y@k}�"w�a$1W2 �!"{$5�ךO��O���8�J�\���MaC�H+�>1�?3B�Dz��D~���%O��ď��ݏ��K	���2x%���"DYWA���1_�/�t��= R�t�r�R���ʟ���� Пޟ�9��#�q`H� ��������a����*3 Ʃ������!��E� W�6�{�Z�l���ÿ�o��b�"��q2��Az&�4���B7YB�#�@�m@$Y*���ʿ B�T�f�x����"H �ܪ������ϑȴ�!� �E�W�i��0ߝߐ� ����r��߮��-�?� Q��u������� �������)�;���_� >�P���t��s����x� h���0' 9f]o���� ����,��O Y�}����� ��(//1/K/U/�/8���/�/  z/�� �/�/??5?(?Y?L? ^?�?�?�?�?�?�?�? �? O1O8UOt/^O�O �O�O�O�O�O�O�O_ _$_Q_H_Z_�_FO�_ �_�_�_�_�_oo o 2oDoqohozo�o�o�o|�oԷ	  �a+��`�����p#Z�`�/- R�=va�C� �<�q
S�����"h�:�2���#���K�����i�A   x����m�@�  Տ��͂С���BѠ=�賖 �����+Ă�C�  �M�3�t��Ӄ>�/{�����S���@@�������BȲS�>����C�����͂��<�o�?�PH�)S�B����������CBܿ�ͅ1�+��9�� m�b�i�!�3���w��]A�����@q�B]���т��¡`  �?��ͥͿ�u�{?����e�ܱ�Ծ�$�DCSS_CLL�B2 2K�����p�~'�NS�TCY 2L����   h�믊�������ҿ� ����,�B�P�b�tπ�ϘϪϼ��Ϸs)�D�EVICE 2Mm���(��>� P�}�t߆߳ߪ߼��� ������C�:�g�y���������)�HN?DGD Nm�p�Cz�k)�LS 2Om�G�9�K�]�o������������PARAM P8�����H��RBT 2R�m� 8�p<�	������Q�T�������R��1��@� �CW  �B\`6�B	D�� ������@R����b���$�����.�� �	>,�YkJk����c��; M�T� ���0///f/��A�S�D �C���ׂ!т1@�#��@I&�@�R�\@g�;?���j��B�&f�B�DC�C3$C2�o�C3Ф����A���B8�y�BB�A��.��m�B���C�R�C3�C4
/C3��a�(�35	P<8�@"E/W/�? ?/m??�?�?�?O�? �?8OO!O3OEOWOiO �O�O�O�O�O�O�O�O __j_A_S_�_�_l� �_�_�_�_o	oBoTo ?oxo�[?�_�_q_�o �o�o�o�o4/ ASe����� �����f�=�O� ��s������_o�� ,��)�b�M���q��� �o��ŏ򟭏۟�:� �#�p�G�Y���}��� ���ůׯ$����Z� 1�C�U���y���ؿ�� ��� ϛ�D�/�h�S� ��wω��ϭ������ �.���)�;�M�_� �߃ߕ��߹������� ��`�7�I��m�� �����������J� \��π�k��������� ������"��+�=�j AS�w���� ��T+=O as����/� �//'/9/�/�/ �/�/�/�/?�/(?? L?^?9g/y/�?}?�? �?�?�?O�?�?OZO 1OCO�OgOyO�O�O�O �O_�O�OD__-_z_ Q_c_u_�_=?�_�_
o oo@o+odoOo�oc? u?�_�o�_�o�o�o N%7I[m �������� !�3���W�i������� ����yo"��F�1�j��|�g�����ğ�h�$�DCSS_SLA�VE S��}���ښ?_4D  ���AR_MENU T� ��R�d�v��������bA�֯��֞'�SHOW 2}U� � �� Ձ/�9�@�^�p�����@������ܿ� � (� "�L�I�[�m�ϑϣ� ʿ��������6�3� E�W�i�{ߍߴϱ��� ������ ��/�A�S� e�w�ߛ������� 
���+�=�O�a��� �������������� '9Kr�[�� ��������# 5\�k}��� ����//1/X U/g/���w/�/�/ �/�/	??B/??Q?x/ �/�/2?�?�?�?�?�? O,?)O;OMOt?nO�? �O�O�O�O�O�OO_ %_7_^OX_�O_�_�_ �_�_�_ _�_o!oH_ Bol_io{o�o�o�o�o �_�o�o2o,VoS ew����o�� ��@=�O�a�s� �������͏ߏ� � *�'�9�K�]�o������"���ɟ��CFG �V������FRA:�\	�L�%04d�.CSV�	��}�֟ ���A O�CHW�z��g�񏋯��
��u�����į֯��u���JP�(����������RC_OUT -W����+�۟�_C_FSI ?�Q�  �u�������޿ٿ� ��&�!�3�E�n�i�{� �϶ϱ���������� �F�A�S�eߎ߉ߛ� ������������+� =�f�a�s����� ��������>�9�K� ]��������������� ��#5^Yk }������� 61CU~y� �����/	// -/V/Q/c/u/�/�/�/ �/�/�/�/?.?)?;? M?v?q?�?�?�?�?�? �?OOO%ONOIO[O mO�O�O�O�O�O�O�O �O&_!_3_E_n_i_{_ �_�_�_�_�_�_�_o oFoAoSoeo�o�o�o �o�o�o�o�o+ =fas���� �����>�9�K� ]���������Ώɏۏ ���#�5�^�Y�k� }�������ş���� �6�1�C�U�~�y��� ��Ư��ӯ��	�� -�V�Q�c�u������� ������.�)�;� M�v�qσϕϾϹ��� �����%�N�I�[� mߖߑߣߵ������� ��&�!�3�E�n�i�{� ������������� �F�A�S�e������� ����������+ =fas���� ���>9K ]������� �//#/5/^/Y/k/ }/�/�/�/�/�/�/�/ ?6?1?C?U?~?y?�? �?�?�?�?�?O	OO -OVOQOcOuO�O�O�O�O�O�O�C�$DC�S_C_FSO �?���Q� P  �O�O<_e_`_r_�_�_ �_�_�_�_�_oo=o 8oJo\o�o�o�o�o�o �o�o�o"4] Xj|����� ���5�0�B�T�}� x�����ŏ��ҏ�� ��,�U�P�b�t��� �����������-� (�:�L�u�p������� ��ʯܯ� ��$�M� H�Z�l���������ݿ ؿ���%� �2�D�m��h�z�_C_RPI^._������Ϩπ_���W߀�{�^SL��@Lߎ��� ��� ��H�C�U�g��� ����������� �� -�?�h�c�u������� ��������@; M_������ ��%7`[ m������ �/8/3/E/W/�/{/ �/�/�/�/�/�/?? ?/?X?S?e?w?�?�? ��9��߬?�?OO+O =OfOaOsO�O�O�O�O �O�O�O__>_9_K_ ]_�_�_�_�_�_�_�_ �_oo#o5o^oYoko }o�o�o�o�o�o�o�o 61CU~y� ������	�� -�V�Q�c�u������� ������.�)�;� M�v�q���������&��NOCODE }X=��'��PRE_CHK �Z=�АA А�< �Ր�=�E�W�=� 	 < 9������3y�ïկ�� ������A�S�-�w� ��c������������ �+�=��a�s�i�[� �ϻ�U���������'� ��]�o�Iߓߥ�� ���ߵ����#���G� Y�3�e��ϗ����� q��������C�U�/� y���e����������� 	��-?KuO a�������� );_qK�� �����/%/� I/[/5/G/�/�/}/�/ �/�/�/?�/E?W? �/{?�?g?�?�?�?�? �?O�?/OAOOMOwO QOcO�O�O�O�O�O�O _+_!?3?a_s___ �_�_�_�_�_�_o'o o3o]o7oIo�o�oo �o�o�o�o�o�oG Y3}�I_w�� ����1�C��/� y���e���������� я�-�?��c�u�O� ��������󟍟� )��5�_�9�K����� ��˯ݯ������� I�[�5����k���ǿ ��ϟ��ϩ��E�� 1�{ύ�gϱ��ϝ��� ������/�A��e�w� Q߃߭߇ߙ������� �+���a�s�M�� �����������'� �K�]�7�����m�� ����������5G =�/}�)��� ����1Cg yS������ �/-//9/c/Yk �/�/E/�/�/�/�/? )??M?_?9?k?�?o? �?�?�?�?OO�?O IO#O5OO�OkO�O�O �/�O�O_�O3_E__ i_{_U_g_�_�_�_�_ �_�_o/o	ooeowo Qo�o�o�o�o�o�O�o +�oOa;m� q������� !�K�%�7�����m��� ɏ��Տ���o5�G� �S�}�W�i���ş�� ���՟�1���g� y�S���������寿� ѯ�-��Q�c��K� ������ϿΏ��� ��M�_�9σϕ�o� ���ϥϷ�����7� I�#�m��u�gߵ��� a�������	�3��� i�{�U������� �����/�	�S�e�?� q����ߣ�����}��� ��Oa;�� q����� 9K%W�[m� �������5/G/ !/k/}/W/�/�/�/�/ �/�/�/?1??U?g? A?S?�?�?�?�?�?�? 	OO/OQOcO�?�O �OsO�O�O�O�O__ �O;_M_'_Y_�_]_o_ �_�_�_�_o�_o7o -O?Omooo�o�o�o �o�o�o�o!3? iCU����� ����	�S�e�?� ����Uo��я㏽�� ��=�O�)�;����� q���͟����ݟ� 9�K�%�o���[����� ���������#�5�� A�k�E�W�������׿ �ÿ������U�g� Aϋϝ�wϩ���ɯۯ 	�ߵ�'�Q�+�=߇� ��s߽��ߩ������ ��;�M�'�q��]�������������$DCS_SGN� [��-��^��>	29-�NOV-25 1�5:52 ��6�0�- 7-31   12:49 `��`� [}S=�n�P�f4n�j��`��k�2�ե�U��Þ�;"0>�~�  �HOW �\��� `��VERS�ION %�V4.5.2���EFLOGIC �1]���  	������+	��:�PROG_ENB  ��"c�[ULSE  @�s_ACCL{IM��u�d�WRSTJN�T�-���EM�Odb�w� IN�IT ^
����OPT_SL �?	���
 	�R575��E7�4J6K7K50o1o +	�(TO  4����V� DEX�d�-�`�#PATHw A%�A\��S/e/��HCP_CLNTID ?��" ,���/���IAG_GRP� 2c������b�	 @��  �"ff?a�G��%��� B�  ?��1� 0C?1>�@c��j2!�7�@�z�@^��@
�!��m�p2m15 89�01234567��0����  �?��?�=q�?��
?޸R�?�Q�?���?ʼ0��0�(��?�z���0`�@o�  AG�Ap�0,�10A� 0 0G�;B4�� ��4�`�
�1@�@���\@~�R@�xQ�@q�@�j�H@c�
@�\��@U�@Mp����?�?D���#@��7IH��@C�\@>L@9��@4�x0/\)@)�@#�\@{@��jO|O�O�O�O8G?�/��?��0�� G@�?}p�?u�?n{?[@?\�0Q��O__,_|>_PX�
=?��0�tP_U� 0z�H�?p�0h��?^�R�_�_�_�_�_PX��5�\P�� � 0�, `�0?�tP�� #` o o2oDoVo8G� ���oAS�o'q� y��[m��+� 	�O�a��m���qbRB��@jRcQ�`
=?�Śʆ�\Pׄ
=5!{��4V����@
=�b��a&���?� �@C��``3=q��=b��=��E1>�J�>��n�>��H
=<w�o ~��s������ �`�C�`<w(�Ub� 4�"i��@ß���A@`�?5������8�J� �Ȼ�V����������xگ쯖�>J����bN�
=��GI�6���@{`^��pPy��0k�@ffZ>9!T@��33푒��(��
=C�� ���I�CH�)�C.dBت 
= B׿ݱɼ'�  � 
��a'�B3Ğ���N�B��`�X��wω� ����Ϸ���`�s��ψo��˻6�<҂��D&t�����D/�´ �²X³��AD
ߋ�߯�����߾��������n���*Iҥ	�W��!C�T_CONFIG� d�'�d��egA�!ST�BF_TTS�
@s	�����e����MAU� h��MS�W_CFv�e�+ � @��OCVIE�W��f	�1�� ��[�m���������� I�����&8�� \n����E� ��"4F�j |����S�� //0/B/�f/x/�/ �/�/�/�/a/�/?? ,?>?P?�/t?�?�?�?X�?�?^�RC�gΥ��!j?��O;O*O_O�NO�OrO�O��SBL�_FAULT �h�:��AGPMS�K���Gj�TDIAOG iz�������UD1�: 67890123451R��%Q���EPD�m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�oLV!V�i��
\_�od�TREC	P
_Z
*TCW{ [_Xj|���� �����0�B�T��f�x��o�o�o���U�MP_OPTIO2%��NځTR��:�I��PME����Y_TEMP  �È�3B+�rO��*�9�UNI�����O���YN_BR�K j4��EDITOR���(����_�`ENT 1k��9  ,&�IP�ANUC_S�MPLGRP_C�LOSEȏ&�FS_MOV_5�DEG �OPED%��������EAS_WRK2�FpG��ANIM=A�_DROq�W���30�K�� ��-BCKEDT-� _PICɯ���HOME �*��&PROG_1� �������J��M�AIN q���&�DE�C���GE�TDATA˿ݿf��1 ���&&��1 �B���AAA �R��&�y϶ϖ�TE�� ?���&@�1 ���&�O4��1䜐MGDI_S�TAb�>�O���NC�_INFO 1l<	������@��ఔߢ�n�V�1m	� C�~�������
��d��=�O�a�s��� �����������'� 9�K�]�o��������� �������	*� 8J\n���� ����"4F Xj|��
��� ��/!+/=/O/a/ s/�/�/�/�/�/�/�/ ??'?9?K?]?o?�? �?�?��?�?�?�?/ #O5OGOYOkO}O�O�O �O�O�O�O�O__1_ C_U_g_y_�_�_�?�_ �_�_�_Oo-o?oQo couo�o�o�o�o�o�o �o);M_q ���_�_���� o%�7�I�[�m���� ����Ǐُ����!� 3�E�W�i�{����� ß՟�����/�A� S�e�w���������ѯ �����+�=�O�a� s���������Ϳ߿� ��'�9�K�]�oρ� �ϥϷ���������� #�5�G�Y�k�}ߏߩ� ������������1� C�U�g�y������ ������	��-�?�Q� c�u����ߓ������� ���);M_q ������� %7I[m�� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?A? S?e?w?���?�?�? �?�OO+O=OOOaO sO�O�O�O�O�O�O�O __'_9_K_]_o_�_ �?�_�_�_�_�?�_o #o5oGoYoko}o�o�o �o�o�o�o�o1 CUgy�_��� ��_�	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ������˟���� �%�7�I�[�m���� ����ǯٯ����!� 3�E�W�i��������� ÿտ�����/�A� S�e�wωϛϭϿ��� ������+�=�O�a� sߍ��ߩ߻������ ��'�9�K�]�o�� ������������� #�5�G�Y�k��ߏ��� ����������1 CUgy���� ���	-?Q c}�o������� �//)/;/M/_/q/ �/�/�/�/�/�/�/? ?%?7?I?[?u��? �?�?�?��?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_�??�_�_�_�_�? �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9K]w_� ����_���� #�5�G�Y�k�}����� ��ŏ׏�����1� C�U�o]�������� �����	��-�?�Q� c�u���������ϯ� ���)�;�M�g�y� ������]�ӟݿ�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�_�q�{ߍߟ߱� ˿��������/�A� S�e�w������� ������+�=�O�i� s��������������� '9K]o� ������� #5Ga�k}�� ������//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Y K?u?�?�?���?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_Q?c?m__�_ �_�?�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/�_ [_ew���_�� ����+�=�O�a� s���������͏ߏ� ��'�9�S]�o��� �����ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� K�9�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����������)�C� �$�ENETMODE� 1n��_�  S�S��N�p߂�R�OAT�CFG o��������C����DATA 1�p_��М��*��*���!�3�E�"T�dT�u몱M�y� �������������� ��E�W�i�{������ ��=�����/A ����w����� �]o+=Oa s������ //��K/]/o/�/�/�/�-R�RPOS/T_LO��r��C%�
���/??/?Q�R�ROR_PR� �%_�%4/q?@8TA�BLE  _�ి�?�?�?�+RSE�V_NUM n�?  �i�@��!_AUTO_ENB  ��g�@4w_NOA s_����B  *�*`@�`@�`@�`@@�+_@yO�O�O9DFLsTR%O7FHISC�E!g�2K_ALM �1t_� �C$`LM�+�O9_K_]_�o_�_�_�O_�2?@  _�^A���ZR��TCP_VER �!_�!`?�_$E{XT� _REQ�Fs�0I*cSIZ3o�%dSTKPiNE��'bTOL  �E!Dz�B�A %d_BWD�P�`�Fعa�ҢcDI�a �u���'��E!�kST�EP�o�oR��`OP�_DOroP�FDR_GRP 1v_��Ad 	�_p��ap�s�Y�q'��M"���l���T� ����vas��}��� ��2��V�A�S����w�����?԰W@�/Ơ@9�?���ܷ�
 F@E"ԁ�����S"� ��F�1�j�U�A����O@S33��P�@�� ��O�؟�ap� �Ŝ�apG�  (�Fg?�fC�8R4�ȝ�?�΀Q�Ǟ6�X��x��875t���5���5`+��ȟH ���?����%V�Ar�EATURE �w���`���LR Handl�ingTool ��E"Engl�ish Dict�ionary��M�ulti Lan�guage (C�HIN)�&�KA�NA/�4D St��ard���An�alog I/O�^�g�gle Sh�iftz�uto �Software Update���matic Ba�ckup�ͱgr�ound Edi�t���Camer�au�Fy�Comm�on calib' UI��n��Monitor(��tr�Reliayb����DHCP���Data Ac�quis7�`�ia�gnosɱr�z�i�splay�Li�cens^�d�oc�ument Vi�eweC�b�ual� Check S�afety#���hanced#�����s��Fr����xt�. DIO 3�f�i��D�end�E�rrB�L��`�8�s�_�rp�O� �`�F�CTN Menu��v^ò�TP I�n��fac����G�igE�����p �Mask Exc��'���HT��Pr?oxy Sv��#�igh-SpeЇSkiҳ#��S�m�municȰonsZ�ur�С�u�v����connect� 2��ncr��sGtru	����e�����J����KARE?L Cmd. ���Run-Ti@�E�nv���el +:̰sʰS/W���������v�Book(System)�MACROs,Q�?/Offse��0�aHSв�s�5�MR<�D8®�M����R�l���MechStop"/�t����0�iqґ�� x�r�ʰ��od>��witch.����.��TOptm�f��0�fi����g���0�-T���P?CM fun���	�a��tiz��o^��Regii�ru��ri��F�4s�Num Sel��|O>� Adjue��Jw���tatu�0�����RDM �Robot�scgove��ea��@�Freq An;lyu�Rem��S��nU���Serv�oS�A ��SNPX� b1�SN��C�li��_.��Libr�/� � K&�oN�t��ssag����P ����a��P�/I���%MILI�B?�"P Fir�m���.P��Acc<��TPTXo��$eln��?�!���-orqu��imGulaA���6uH �Pa*��.�\�b&�/�ev.�%��ri���t?USR E�VNTO-@nexOcept� n��X(E9�{�VC�rp�g���V���B<?�E�+��KSr SCn5�OS�GE�O�EUIa�Web Pl�^=!���ET7������ZD?T Appln��QEOAT�!Ѵ���iPj�ax)�_ G�rid����]�_iR�B.U�f���O���RX-10iA��_m�ll Smo�othU���c�sc�ii/�vLoad���tjUpl�`��t�oS��0rity�AvoidM,�sbW�t�0g`	�yc��`�;@�c�CS/��. c�� xJo =tL�r x��u��� xc��abo���RL�0>�2Y�Ճor��O�0�S�F�it��{tl�n�t���wHMI Dev�� (S!m�����in�#?�
����sswo\���R?OS Eth(��a@�!��$�[L%�g �b�L%dhUpvE!�%f[�t �НiRs���{�64MB D�RAM��FROp#����l<f FlH�����6m �aZ�op�q���e``v��sh�����Ɨc�Õ��p,�6؜ty��saȂ)�r'��j"~ .z�pq/sJs�dŰ �vx��� 2�ap�pornv��<"�V�q�T1*�FC�/��E�Fs=��H�el�U!��Typ��FCE h��vR@aSt�{����luA x$ꃨPG j����Rj��No md �c߷ dOL;��Sup���0OP'C-UJk"�T遼�05��j��cr.p��lu� �����quir��� Om��%p�T0.
���estL%?IMPLE ��V�J'S;�eq�tex��dhz�I(p��[B�?CPP���E����bTeaH �9�ߚDrtu���v�Y����4���UIFg�po�nsRfstdpn�Ke SWIMEoST f� F01���� bC�:�L�y�p� ���������	� � �?�6�H�u�l�~��� ����������; 2Dqhz��� ���
7.@ mdv����� ��/3/*/</i/`/ r/�/�/�/�/�/�/�/ ?/?&?8?e?\?n?�? �?�?�?�?�?�?�?+O "O4OaOXOjO�O�O�O �O�O�O�O�O'__0_ ]_T_f_�_�_�_�_�_ �_�_�_#oo,oYoPo bo�o�o�o�o�o�o�o �o(UL^� �������� �$�Q�H�Z���~��� �����؏��� � M�D�V���z������� ݟԟ��
��I�@� R��v�������ٯЯ ����E�<�N�{� r�������տ̿޿� ��A�8�J�w�nπ� �Ϥ����������� =�4�F�s�j�|ߎߠ� ����������9�0� B�o�f�x������� �������5�,�>�k� b�t������������� ��1(:g^p �������  -$6cZl~� ������)/ / 2/_/V/h/z/�/�/�/ �/�/�/�/%??.?[? R?d?v?�?�?�?�?�? �?�?!OO*OWONO`O rO�O�O�O�O�O�O�O __&_S_J_\_n_�_ �_�_�_�_�_�_oo "oOoFoXojo|o�o�o �o�o�o�oK BTfx���� �����G�>�P� b�t�������׏Ώ�� ���C�:�L�^�p� ������ӟʟܟ	� � �?�6�H�Z�l����� ��ϯƯد����;� 2�D�V�h�������˿ ¿Կ���
�7�.�@� R�dϑψϚ��Ͼ��� �����3�*�<�N�`� �߄ߖ��ߺ������� �/�&�8�J�\��� ������������+� "�4�F�X���|����� ����������'0 BT�x���� ���#,>P }t������ �//(/:/L/y/p/��/�/�/�*  ?H551�#�!�2�(39�(0�%R�782�'56J6{14�%ATUP'6�545'86�%VC{AM�%CUIF'7�28c6NRE65�2V6R63�&RS�CH�%LIC�6DwOCV�6CSU6�866J6026E�IOC�746R6=9V6ESET?7U7�J7U7R68�&M�ASK�%PRXY�o87�&OCOH3�?86@&83^FJ6�%8 :�GLCHFFO�PLG?70vFMH�CRGFS�GMAT��6MCS>80"G5=526MDSW+WiG;OPiGMPRjF�0��H06PCMn75`qW@26�@�G51J7�51�X0J6PRSvG69^FFRDb6�FREQ6MCNz�&97SNBA�7^�GSHLBfM1gt�0X26HTC>6�TMIL86TP�A�6TPTXcfELf�@�7870�&wJ95z6TUTjFwUEVFUECFFwUFRb6VCC�h�O�FVIPnfCS�C�fCSG�6�0I��%WEB>6HTT�>6R6�8�h;0FvC�G]wIGEwIPGmS�vRCnfDGiGkH7�X6�'R7	G]R�XR51�86vH%2vH5V6�0JX�X�6z7L=i�'J87�"G87�G83J6R�55vF@26R64��g5��R6�GR8�4��79�H4z6S�5]GJ76^FD0u626F �RTSfwCRDFCRXjF�CLIZXI7CMS��6S�>6STYng6�)WCTO>6�0�778�7�0z6ORS�F7@�6FCB�6FCFv�WCH>6FCRF�FCI�vFC�GJԋpOWG*�M�XNO�M�6OLWKP�6O�P��SENDGFL]U�FCPR�WL	wuS��C�8ETS^��T��0zgCP�6TE�%�S60�&FVR��6IN�WIHagI{PNnfGene�$ �(1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������ /ASew��� ����+= Oas����� ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e�w������� ��џ�����+�=� O�a�s���������ͩ�  H5�51ϧ�2�39z��0�R782﫽5�J614�AwTUP?�545?��6�VCAM�C�UIF?�28��N�RE�52~�R6�3�RSCH�L{IC��DOCV���CSU�86�J{60N�EIOC���4.�R69~�ES�ET_�}�J7}�R{68�MASK﩯PRXY��7�OCO�3_�.���>��3��J6=���L{CH��OPLG_��0��MHCR��S�}�MAT��MCS�^�0��55N�MD�SW����OP��M�PR��۰.�0�PCM��5M��N��ж.�51n�51��0nn�PRS~�69���FRD��FREQ��MCN�9�S�NBAϻ�SHLEB�MM�۰��2��HTC^�TMIL���TPAN�TPTX��EL���.�q8-�+��J95��wTUT��UEV~�wUEC��UFR���VCC^O��VI�P��CSC��CS�G���I�WEBn^�HTT^�R6ͼ���[��
CG�IG޽IPGSRC���DG��H7m�6��R7m�R��R5U1^�6��2��5~�R�J�ܞ�6��L]�n�J87��87.�;83n�R55��k��N�R645�+R�6��R84n+79��4��S5��J7]6��D06N�F<wRTS.�CRD~�wCRX��CLI.�m�CMSN�{0^�S�TY��6��CTO�^��N�7-�˰��O�RS�ګ��FCBnN�FCF��CH^�wFCR~�FCI>KFC��J�G��M��NOMN�OL�����OP]KSE�ND��LU~�CPUR��LmS�<C̇ETS�K|<;���C�P��TE=;S60n�FVRN�IN��IH��IPN��Gene�Ψ�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y��k�}�������ů  }נSTDҤ?LANG�� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z�x������RBT�OPTN������	 -?Qcu�������DPN �);M_q �������/ /%/7/I/[/m//�/��/�/�/�/�/�/?ted �ʨ9? K?]?o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�_�_�_�_�_	o o-o?oQocouo�o�o �o�o�o�o�o) ;M_q���� �����%�7�I� [�m��������Ǐُ ����!�3�E�W�i� {�������ß՟��� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9� K�]�oρϓϥϷ��� �������#�5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u����� ����������) ;M_q���� ���%7I [m��������/!/3/E/  �N/l/~/�/�/�/�-�99�%�$FE�AT_ADD ?_	����!0?  	�(? ?/?A?S?e?w?�?�? �?�?�?�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy� ������	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q���������˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a�s߅ߗߩ߻� ��������'�9�K� ]�o�������������$DEMO �w�)    �(4�*�<�i�`�r��� ������������/ &8e\n��� �����+"4 aXj����� ���'//0/]/T/ f/�/�/�/�/�/�/�/ �/#??,?Y?P?b?�? �?�?�?�?�?�?�?O O(OUOLO^O�O�O�O �O�O�O�O�O__$_ Q_H_Z_�_~_�_�_�_ �_�_�_oo oMoDo Vo�ozo�o�o�o�o�o �o
I@R v������� ��E�<�N�{�r��� ������ԏޏ��� A�8�J�w�n������� ��Пڟ����=�4� F�s�j�|�������̯ ֯����9�0�B�o� f�x�������ȿҿ�� ���5�,�>�k�b�t� �ϘϪ���������� 1�(�:�g�^�pߝߔ� ���������� �-�$� 6�c�Z�l����� ��������)� �2�_� V�h������������� ����%.[Rd �������� !*WN`�� ������// &/S/J/\/�/�/�/�/ �/�/�/�/??"?O? F?X?�?|?�?�?�?�? �?�?OOOKOBOTO �OxO�O�O�O�O�O�O ___G_>_P_}_t_ �_�_�_�_�_�_oo oCo:oLoyopo�o�o �o�o�o�o	 ? 6Hul~��� �����;�2�D� q�h�z�����ˏԏ ���
�7�.�@�m�d� v�����ǟ��П���� �3�*�<�i�`�r��� ��ï��̯����/� &�8�e�\�n������� ��ȿ�����+�"�4� a�X�jτώϻϲ��� ������'��0�]�T� f߀ߊ߷߮������� ��#��,�Y�P�b�|� ������������ �(�U�L�^�x����� ����������$ QHZt~��� ��� MD Vpz����� �/
//I/@/R/l/ v/�/�/�/�/�/�/? ??E?<?N?h?r?�? �?�?�?�?�?OOO AO8OJOdOnO�O�O�O �O�O�O_�O_=_4_ F_`_j_�_�_�_�_�_ �_o�_o9o0oBo\o fo�o�o�o�o�o�o�o �o5,>Xb� �������� 1�(�:�T�^������� ����ʏ��� �-�$� 6�P�Z���~������� Ɵ����)� �2�L� V���z�������¯� ���%��.�H�R�� v������������� !��*�D�N�{�rτ� �ϨϺ��������� &�@�J�w�n߀߭ߤ� ����������"�<� F�s�j�|������ �������8�B�o� f�x������������� 4>kbt ������ 0:g^p�� ����	/ //,/ 6/c/Z/l/�/�/�/�/ �/�/?�/?(?2?_? V?h?�?�?�?�?�?�? O�?
O$O.O[OROdO �O�O�O�O�O�O�O�O _ _*_W_N_`_�_�_ �_�_�_�_�_�_oo &oSoJo\o�o�o�o�o�o�o�o�o}  x.@Rdv �������� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ����"�4�F� X�j�|�������į֯ �����0�B�T�f� x���������ҿ��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
.@Rdv ������� *<N`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6 HZl~���� ���� �2�D�V� h�z�������ԏ� ��
��.�@�R�d�v� ��������П���� �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������  ��2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ��(�:�L�^�p��� ������������  $6HZl~�� ����� 2 DVhz���� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|����@���������� ��6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p ������� � �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ� ������������0� B�T�f�x������ ��������,�>�P� b�t������������� ��(:L^p �������  $6HZl~� ������/ / 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFoXojo|o�o�o��o�o�o�o�oy��$FEAT_DEMOIN  #t��Np�$p6tI�NDEXC{Rq��6pILECOMP x����q�Qr1uzpSETUP2 y�u��r�  N� �qws_AP2B�CK 1z�y � �)x��{%� �$p�p�K�!u �w����*���я`� �����+���O�ޏs� �����8�͟ߟn�� ��'���4�]�쟁�� ����F�ۯj������ 5�įY�k�������� B����x�Ϝ�1�C� ҿg����ϝ�,���P� ���φ�ߪ�?���L� u�ߙ�(߽���^��� ���)��M���q�� ��6���Z������ %���I�[������� ��D���h�����3 ��W��d��@ ��v�/A� e���*�N��r�/�y�pP�� 2�p*.VR /j/�*m/�/�0�/�/�T PC�/�/>�FR6:�/>�/>?�+Tbpb?t?�5_?�<Ep/?�?�G*.FW/�?�	3��?"L�?FO�;ST�MQO{O20gO�M5O�O�;H�O�O�G�Op�O�OO_�:GIFY_��_�Eo_,_>_�_�:JPG�_o�E�_�_�_�Wo�*JSao�o��cxo5o%
JavaScript�o�_CS�o�F�o�o� %Casca�ding Sty�le Sheet�s:�
ARGN?AME.DTi��@\};�a�t��j�pDISP*���t���q4��B��CLLB.cZI_��@:\���\��Ɖ�aCol�laboƏr�
PANEL1�O ��s�	�C��qiPend�ant Pane�lJ��	9�:�"�@5���R�d����2?��(�3��ԟ�{���2 ß������X�j����3G�0�3��ܯ���3˯������`�r���4O�8�3�&�����φ�4ӿ�Ϸ����h�z��vtTPEI?NS.XML�=��:\)��ϥqCus�tom Tool�barj��yPAS�SWORD����FRS7���n�P�assword ?Config�ߥ 7���0�m���� �� ��V���z��!���E� ��i���
���.���R� ��������AS�� w��<�`� ��+�O�H� �8��n/� '/9/�]/��//"/ �/F/�/j/�/?�/5? �/Y?k?�/�??�?�? T?�?x?O�?�?CO�? gO�?`O�O,O�OPO�O �O�O_�O?_Q_�Ou_ _�_(_:_�_^_�_�_ �_)o�_Mo�_qo�oo �o6o�o�olo�o% �o�o[�ox� D�h���3�� W�i�������@�R� �v�����A�Џe� 􏉟��*���N���� �����=�̟ޟs�� ��&���ͯ\�񯀯� '���K�گo�������4�ɿX�j�����$�FILE_DGB�CK 1z������� < �)
SU�MMARY.DG�	���MD:=�}����Diag S?ummary~��CONSLOGsϠV�h���ߐ��s?ole lo	TPACCN���\�%D߁ߌ�TP� Account�in#ߋ�FR6�:IPKDMP.'ZIP�߹�
�����ŝ�Except�ion
��i�ME?MCHECKw����lύ��Memory Data���Jn )x�RIPE��f�x�����%�� Pac�ket L"��L��$�K���STA�T��� ��� �%)�Statuys��F�	FTP�����|������mment TBD�F� >I)ETHERNE_���L��]���Ethe�rn2��figu�ra)DCSVRF������  verif�y all"�(�14�DIFF���#�9di�ff�ZL�� CHG01���)/��X�Q/\2��2/�//�/�N/`/�3p�/�/�/1? �/�X?�&VTRND?IAG.LS]??� ?�?��u1 Op�e�4� ��nos�tic�׉�)�VDEVy2DA�T�?�?�?�?��V�is�1Devic9e�?�;IMGy2���O&O�O"�QDImsag]O�;UP@�ESO�OFRS�:\_B]��Up�dates Li�stB_���@FL?EXEVEN��O�O�_���Q UI�F Ev55��-�vZ)
PSRBWLD.CM�_µ�-R	oD_�PS�_ROBOWEL<;�:GIG��o��_�o��GigE��H�_�N�@�)}�aHADOW�o�o�oO��Sha�dow Chansge����Cdtr?RCMERRG,�>����pCFG� ErrorW@t�ailv MA��S�CMSGLIB���Y��b����bPic ���)E�ZD�o��B�׏n��ZD�`ady��� rNOTI����ȏ]���Notific����,�AG)CR?SENSPK�O�����\���� CR�_ؑOR_PEAK柍�.�@��d�� �������M��q�� ���<�˯`����� %���̿����ϣ� %�J�ٿn����Ϥ�3� ��W���{ύ�"߱�F� X��|�ߠ�/߱��� e��߉��0��T��� x����=������ ���,���=�b���� �����K���o��� ��:��^p+�# �G��}�6 H�l��1� U��� /�D/� U/z/	/�/-/�/�/c/ �/�/?�/�/R?�/v? �?C?�?;?�?_?�?O �?*O�?NO`O�?�OO �O7OIO�OmO__�O 8_�O\_�Om_�_!_�_ E_�_�_{_o�_4o�_ �_jo�_�o�o[o�oSo �owo�o�oB�of x�+�Oa� ��,��P��t�� ����9�Ώ]����� (���L�ۏ폂���� ��s�ܟk� ����6� şZ��~������C��دg�y����$F�ILE_FRSP�RT  ���������'�MDONLY �1z;��� 
 ���~�˯��ﯯ� ؿ������ �2���V� �zό�ϰ�?����� u�
ߙ�.߽�;�d��� ��߬߾�M���q�� ��<���`�r��� %��I��������� 8�J���n������3� ��W�������"��F���S|%�VISB�CKY�C�h�*.�VD��; FR�:\� ION\DOATA\�^; �Vision VD file� ASiwa�* ��`��/+/� O/�s///�/8/�/ �/�/?�/'?�/8?]? �/�??�?�?F?�?j? �?�?�?5O�?YOkO&O �OO�OBO�O�OxO_ �O1_C_�Og_�O�__�,_�_!�LUI_C�ONFIG {�;���[ $ �S^��V#o5oGo`Yoko}o�i`|x�_ �o�o�o�o�o|�o0 BTfx��� �����,�>�P� b�t��������Ώ�� 򏉏�(�:�L�^�p� �������ʟܟ� �$�6�H�Z�l���� ����Ưدꯁ�� � 2�D�V�h��������� ¿Կk��
��.�@� R��vψϚϬϾ��� g�����*�<�N��� r߄ߖߨߺ���c��� ��&�8�J���n�� ������_������ "�4�F���j�|����� ����[�����0 ��Afx���E ���,�P bt���A�� �//(/�L/^/p/ �/�/�/=/�/�/�/ ? ?$?�/H?Z?l?~?�? �?9?�?�?�?�?O O �?DOVOhOzO�O#O�O �O�O�O�O
_�O._@_ R_d_v_�__�_�_�_ �_�_o�_*o<oNo`o ro�oo�o�o�o�o�o �o&8J\n� �������t�Robot S�peed 100%�:�L�^�p����r�  x������$FLUI_DA�TA |��}�Ł�q���RESULT �3}Ņ� ��T�/wiz�ard/guid�ed/steps/Expert�� %�7�I�[�m�������ǟٟ��Co�ntinue w�ith G�ance�"�4�F�X�j��|�������į֯� ���-��Ņ�0 ��p�ǃƁ6'����ps�r� ��������̿޿�� �&�8����_�qσ� �ϧϹ��������� %�7ߏuт�q'��+�z=�+M�cllb�ToolSet���g/Dist�Work@�������%�7�I�[�m���.0����������� ��%�7�I�[�m�����w{ݐqo߁�?��&M�rip���N�um/NewFram�+=Oas���������0x��
.@R dv��������p��c�/��E��M���imeUS/DST�y/�/�/�/ �/�/�/�/	??-?�?Enabla? s?�?�?�?�?�?�?�?POO'O9O���`/sO5/G/Y&24d/ �O�O�O�O_#_5_G_ Y_k_}_<?N?�_�_�_ �_�_oo1oCoUogo yo�oJO\OnO�OB���>
�ditor�o /ASew������� Touc�h Panel �s (recommen�)�$�6� H�Z�l�~�������Ə؏� ��o�o��o|�oracces`� p���������ʟܟ�� ��$�?�Con�nect to Netw��g�y��� ������ӯ���	��-�싘O���#����!E�pIntroduction6� ˿ݿ���%�7�I� [�m���u��ϰ��� ������
��.�@�R� d�v߈����]��߁���Us�_#�5� G�Y�k�}���������q1����%� 7�I�[�m�������������a
������ߤ����)����A��ve���{����������
0xFE/^p�� ����� //$/2*�c.L/ 2~D/Macro�s/New�"_��/ �/�/??(?:?L?^?|p?�?�0x0�? �?�?�?�?�?OO)O ;OMO_OqO�OB&��]/��O�/�,�/�+�"Open�#_5_G_Y_ k_}_�_�_�_�_�?�� �_oo1oCoUogoyo �o�o�o�o�o�����O��O��-�O�OoClos�w�����������_2 +�Q�c�u��������� Ϗ����)��o�i�R���=��S�etMethod .���ӟ���	��-��?�Q�c�u�8�c��[�����W��n�𒼐��������̯ޯ ���&�8�J�\�n��� ="iqr�Oa��s���$����tra�ightOffset���,�>�P�bπtφϘϪϼ���=��X�g����g ������,�>�P�b߀t߆ߘߪ߼��ߍ�l0�����ѿ�%�S�M�X��o���� �����������#�>.0<�'�Q�c�u� ��������������$)A��h ��+�=�O�Y*��� �/ASew 6�������/ /+/=/O/a/s/2D`V�/z��tZ~/ ?)?;?M?_?q?�?�?�?�?�?�117.762��?OO 1OCOUOgOyO�O�O�O��O�/�/�$B�%ȯ/�/׺)�/��Ro�tationIWW �Oo_�_�_�_�_�_�_��_�_o�?180 �Ko]ooo�o�o�o�o �o�o�o�o#�OX�C3�_%_7_I_onP&����� �/�A�S�e�$o��� ����я�����+� =�O�a�s�2�/�/hz��nRz��)� ;�M�_�q���������x�-99o��� (�:�L�^�p�������0��ʿ����´������,"ݟ�tp3Z�dir/Tp3z οd�vψϚϬϾ��� �������?<�N�`� r߄ߖߨߺ������� ��ӿ��O��� �+1��Measu�rement/S?traigh?�� ��������+�=�O� a� �2ߗ��������� ��'9K]o�.�@�R�d�v��/W�e��Nums/New�sv'9 K]o����v�0x��� //$/ 6/H/Z/l/~/�/�/�/�/-`��)��#�y.��Tool�Use�/l?~?�?�?��?�?�?�?�?O)j1OAOSOeOwO�O�O �O�O�O�O�O__-a	
�/���/Y_?-?�PartR?�_�_ �_�_�_o#o5oGoYoko*B2oo�o�o�o�o �o�o%7I[�m,_��K_��(�_�s/G���r � �2�D�V�h�z������������ ��0�B�T�f�x��� ��������{}���#�)��yPayl?oad1Cm�b� t���������ί�������p�[��c�Ȃ��c-���L�^�p����� ����ʿܿ� ��}�ٟ�/5���3��Y ϶����������"��4�F�X�j��10 ׏�ߤ߶��������� �"�4�F�X�j�՟WɃA ��[���=�2 O���,�>�P�b�t����������'��ێ�5��� $6H Zl~���υ�C����}P&����Advanced� \n������p��/{�0x�� :/L/^/p/�/�/�/�/@�/�/�/ ??u����1?u�%%��M�ass/Center�1?�?�?�?�? �?	OO-O?OQOcOҏ �O�O�O�O�O�O�O_ _)_;_M___v�0?�0�_f?��?ss��j_ oo+o=oOoaoso�o �o�ohOzO�o�o '9K]o���@�v_�_�_�_�[,�_J��G.c�2�XX� ^�p���������ʏ܏ � ��o�o6�H�Z�l� ~�������Ɵ؟��� ������'�9�sY���į֯��� ��0�B�T��%��� ������ҿ����� ,�>�P�b�!�3�E�W�i�{���sZf��� *�<�N�`�r߄ߖߨ� g�y�������&�8� J�\�n�����uϐ�ϙϫ�.����p �P�\L�[�m������ ��������������3 EWi{���� ��������� ��$�6�rt���� ���	//-/?/Q/ "�/�/�/�/�/�/ �/??)?;?M?_?�0BTfx�rt ��OO'O9OKO]OoO �O�O�Od/v/�O�O�O _#_5_G_Y_k_}_�_ �_�_r?�?�?�?���<�TCPVerif�y/2cMethod�_Vohozo�o�o�o��o�o�o�o�LDi�rect Entry8J\n� ��������HA�_'��_�_j'o+ofyJ�����ȏڏ ����"�4�F�X��O |�������ğ֟��� ��0�B�T��_A��_0��[�m��fy��� 
��.�@�R�d�v��� ����k�п����� *�<�N�`�rτϖϨπg������ϯ���ӯfy�?L�^�p߂ߔߦ���������� ￰1?17.762ǿ/� A�S�e�w�����������������B냆%������/mW �������������`1CU�80ÿ ��������!3EW�D�CA39�G�Y�k�}�PZ �//+/=/O/a/s/ �/�/�/���/�/�/? ?'?9?K?]?o?�?�? �?d���Ϛ���yR�?IO[OmOO�O��O�O�O�O�O�O�-9m&_8_J_\_n_�_ �_�_�_�_�_�_�_�?F�9´�?�?L*O~#OfyMeano �o�o�o�o�o�o0B_*gtS�� �������"� 4�F�oou�3oEoJ1)eowo�`axV�� ��)�;�M�_�q��� ��Tf˟ݟ��� %�7�I�[�m������ b�������K"��ˁ�Introductio�o?�Q�c�u� ��������Ͽ��% �2�$�6�H�Z�l�~� �Ϣϴ��������ϵ A��ѯ���B� ˀ ߇ߙ߽߫����� ����)�;�M��q� ������������ �%�7�I��6�,�>�� M#a�file2�/cyclepo=wƆmodeT��� ��1CUgy����#�z�b��g�X�^�[�g���� 0BTfx���&-e�!� �������La�uide�dȄSafety �5/G/Y/k/}/�/�/ �/�/�/�/T�??1? C?U?g?y?�?�?�?�?�?�?�?g�g��Ox�����/don�� �O�O�O�O�O�O�O_  _2_D_?h_z_�_�_ �_�_�_�_�_
oo.o @o�?O#OmoGO/ȄReg,��o�o�o "4FXj|���?EuropO� ����#�5�G�Y�Pk�}�����abzc�o}o�oML�o Toimez}@EU�� 5�G�Y�k�}��������şן韨wEETw Ea rn �sa�o+�=�O�a�s����������ͯ߯񯰇�c`�ߏя㏡o��24����������Ϳ ߿���'�9�P_]� oρϓϥϷ������� ���#�5�G�^o�*��<�RO`�24/currentL����� ��)�;�M�_�q�����s29-NO�V-25 17:29 ��������� �*�<�N�`�r������_����yߋߝ� <�߿�Year��2 DVhz��������v2025 �*<N`r�������� 
<����  ���-/��!��Month��/�/�/�/�/�/��/??)?;?�u11C?j?|?�?�?�?�? �?�?�?OO0OBO/' /�O�U/��DayFO�O�O�O_ !_3_E_W_i_{_�_L829�_�_�_�_�_o o*o<oNo`oro�o�oUOgHsO�o���O��Hou -?Qc u������L97��$�6�H�Z�l� ~�������Ə؏ꏩo"gH�o)���"�og(inute��� ����̟ޟ���&� 8��_\�n��������� ȯگ����"�4�� ��o-�;�Q Q���?NetDonr�ѿ �����+�=�O�a� sυ��nA�ϻ����� ����'�9�K�]�o��ߓ�W�W����ߍ� O"��	��-�?�Q�c� u���������� ��)�;�M�_�q���@����������I��� �߽�����Xj| ������� 0��Tfx�� �����//,/ ����!3E�/�/ �/�/�/??(?:?L? ^?p?�?A�?�?�?�? �? OO$O6OHOZOlO ~O�OO/a/s/�/�/�O _ _2_D_V_h_z_�_ �_�_�_�_�?�_
oo .o@oRodovo�o�o�o �o�o�o�O�O�O�O���W�Summary �ov������ ���*��_N�`�r� ��������̏ޏ��� �&�8���	-?���RobotOp <�ʟܟ� ��$�6� H�Z�l�~�=�����Ư د���� �2�D�V�h�z���O�O�a���􅟗�&��cllb�WtToolSet�ting�Off ��(�:�L�^�pςϔ�`�ϸ����ϛ�1�� ��)�;�M�_�q߃�@�ߧ߹����ߣ�
�i ͷK���%��n��{��������@������/���23� Y�k�}����������������1�����q��.E�/�S�peedLimit/Max�6� �� 2DVh�z��	1000.�0������ /!/3/E/W/i/{/�+yIsDz  g�y����Val �/,?>?P?b?t?�?�? �?�?�?��OO(O :OLO^OpO�O�O�O�O��O�O�/�/�/�/����//Introductioi�p_�_ �_�_�_�_�_�_ oo $o��HoZolo~o�o�o �o�o�o�o�o 2 M���M'_��A_� �lectWork 4������/��A�S�e�w�6iLi_ghtwe�� �qpiece����Ϗ ����)�;�M�_�\q���  Er��Sew�4�/L�oad�NotH'W_l��W�W���� .�@�R�d�v�������8��Я;d.3�?�� �"�4�F�X�j�|��������Ŀֿ�OÙ>�#����ɟ7�8�����CenterMassڿ�ϘϪϼ� ��������(���? Q�c�u߇ߙ߽߫��� ������)���C���3Z5=�O�a�omml�.����������1�C�U�g�y�<c�EOAT w/o par������� ����
.@Rdv;xA﫟�w��/ ����+=Oa s�����8�� //'/9/K/]/o/�/ �/�/�/�/4�X����2��g�n? �?�?�?�?�?�?�?�? O"O�FOXOjO|O�O �O�O�O�O�O�O__`�/�/?c_%?�/9? K?���_�_�_�_
oo .o@oRodovo���_�o �o�o�o�o*< N`r�C_��y_�+�_���"�4� F�X�j�|�������ď�h10;O���� ,�>�P�b�t�������0��Ο9_�yA Y_� }_��~a?k�}����� ��ůׯ�����6O C�U�g�y��������� ӿ���	��ڟ�V_`�"�,5�G��_���� ������*�<�N�`�tr߉b�cith�o �߷����������#� 5�G�Y�k�<Ϧ���r��6��/� Co�ntactSto�pInvalid�Area/�PlusZz�$�6�H�Z� l�~���������ݏ�� �� 2DVhz ����-ϓ�������7�����Min�v����� ��//��</N/`/ r/�/�/�/�/�/�/�/ ??������51C�XY	�XY"?�?�?�?OO%O 7OIO[OmO,/�O�O�O �O�O�O�O_!_3_E_�W_i_(?:?L?^?p?���)�?��NotHW_l�o!o3oEo Woio{o�o�o�o�o�A R��o�o&8J \n������PA�_����_���_ U����\�n������� ��ȏڏ�����o4� F�X�j�|�������ğ ֟�������9����� -��1Spe?edLimio�� ïկ�����/�A� S�e�$���������ѿ �����+�=�O�a�@s�2�D���h��S����Modet��� )�;�M�_�q߃ߕߧ����|GDo no�t Use (R�ecommended)�� ��$�6� H�Z�l�~��������"���ϡϳ� �\��9�K�]�o����� ������������|� 5GYk}���@����yH�� ���7�#���� ����//*/</ N/`/�/�/�/�/�/ �/�/??&?8?J?\? -?Qcu�?�? �?O"O4OFOXOjO|O �O�O�Oq/�O�O�O_ _0_B_T_f_x_�_�_ �_�_?�?�?�?�?,o >oPoboto�o�o�o�o �o�o�o�O(:L ^p������ � ���_�_�_oo ~�������Ə؏��� � �2�D�V�g��� ����ԟ���
�� .�@�R�d�#���G�Y� k�Я�����*�<� N�`�r���������˯ ޿���&�8�J�\� nπϒϤ϶�u��ϙ� ����"�4�F�X�j�|� �ߠ߲���������� ˿0�B�T�f�x��� �������������)� ��M����������� ������(:L ^������ � $6HZ� {=��a�u��� / /2/D/V/h/z/�/ �/�/o�/�/�/
?? .?@?R?d?v?�?�?�?�k���?��/�wizard/c�llb/step�s/Summary�?HOZOlO~O�O�O �O�O�O�O�O�/ _2_ D_V_h_z_�_�_�_�_ �_�_�_
o�2�7�?��?�?�(O/Co�nfigurat�ionCompleteo�o�o�o�o �o(:L^_ ������� �@�$�6�H�Z��6#o�5o�Yo�3qo/S�ignalNum�berAssـment/SPIރ d�	��-�?�Q�c�u�0������ju1��ٟ ����!�3�E�W�i� {��������1
�9��a���2ŏ׏�D�U�g�y������� ��ӿ������-�?� Q�c�uχϙϫϽ��� �����į֯�����
ߐߢߴ����� ����� �2�D�V�m z������������@
��.�@�R��:� ��{�U�������� &8J\n�� �c�����" 4FXj|���?�?�������/./ @/R/d/v/�/�/�/�/ �/�/�/�?*?<?N? `?r?�?�?�?�?�?�? �?O���GO	/nO �O�O�O�O�O�O�O�O _"_4_F_?W_|_�_ �_�_�_�_�_�_oo 0oBoToOuo7O�o[O �o�o�o�o,> Pbt����o� ����(�:�L�^� p�������eoǏ�o� �o�$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ������ۏ =����v��������� п�����*�<�N� �rτϖϨϺ����� ����&�8�J�	�k� -��ߡ�e��������� �"�4�F�X�j�|�� ��_����������� 0�B�T�f�x�����[� ���������,> Pbt����� ����(:L^ p������� ������/E/l/~/ �/�/�/�/�/�/�/?  ?2?D?h?z?�?�? �?�?�?�?�?
OO.O @O�/#/5/�OY/�O �O�O�O__*_<_N_ `_r_�_�_U?�_�_�_ �_oo&o8oJo\ono �o�o�ocOuO�O�o�O "4FXj|� ������_�� 0�B�T�f�x������� ��ҏ����o�o�o;� �ob�t���������Ο �����(�:��K� p���������ʯܯ�  ��$�6�H��i�+� ��O���ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ�Y��� }��ߡ���*�<�N� `�r��������� ����&�8�J�\�n� ���������������� ��1����j|� ������ 0B�fx��� ����//,/>/ ��_/!�/�/Y�/�/ �/�/??(?:?L?^? p?�?�?S�?�?�?�?  OO$O6OHOZOlO~O �OO/�/s/�O�O�/_  _2_D_V_h_z_�_�_ �_�_�_�_�?
oo.o @oRodovo�o�o�o�o �o�o�O�O�O9�O `r������ ���&�8��_\�n� ��������ȏڏ��� �"�4��o)�� M��ğ֟����� 0�B�T�f�x���I��� ��ү�����,�>� P�b�t�����W�i�{� ݿ����(�:�L�^� pςϔϦϸ����ϛ�  ��$�6�H�Z�l�~� �ߢߴ������ߩ��� Ϳ/��V�h�z��� ����������
��.� ��?�d�v��������� ������*<�� ]�C���� �&8J\n �������� /"/4/F/X/j/|/�/�M�/q�/�+�$F�MR2_GRP �1~�%�� �C4  �B�� 	 � x!?3<0F@ I?y@�+0G�  q1�Fg�fC�8R<}5a=?�  �?�,�06�X��2�8�75t��5��ߛ5`+�a=A�3  �?�;BH�4_0�E@S33!E�,4COTM0@AjO`> TO�O�O�O�O�O�O_ �O2__/_h_S_�_�#��"_CFG ;T32�_�_�_�_�Y�NO :
�F0.a 3`�\RM�_CHKTYP  �!� 00� �!�ROMI`_MIN\O`�#��{`�:@]X� SSB�S��% 6��o�%�c�o�o�UTP�_DEF_OW � �$3�gIR�COMN` �$G�ENOVRD_DeOpf�-}TH�0�rd dJud3t_E�NB 3pRA�VC�#��g�` �A5�o�y_�a<q��1J �q�OU 0�<6a818r15<x`�?���/�}���͏�#C���3�!���o"��!>W����Br0�p49p��o�pSMT�#ሡy0�`��$HoOSTC�R1�9Ν`���0 M5C�$
�ȟ�&  27.0�=1�  e��E� W�i�{��*3�����Я�������	ano?nymous	�7�I�[�m�� ǟ0���������,�	�� -�?�QϘ�uχϙϫ� οh������)�;� ���Ϧ�������� ������Z�7�I�[� m������������� ���V�h�zߌߎ�{� �ߟ���������.� /ASv���m� ����*�<�N�+ bO��s����� ���//8�� ]/o/�/�/�/�� "$/?X5?G?Y?k? }?��?�?�?�?�?? B/T/1OCOUOgOyO�/ �/�/�O�?�O,?	__ -_?_O�Ou_�_�_�_ �O�_O�_oo)o;o �O�O�O�O�_�o�O�o �o�oZ_7I[ m�o�_�_������|���ENT {1�P� P!�.V�  'pD��� p���h�ɏ��폰��� ԏ"�G�
�k�.���R� ��v�ן�����П1� ��U��y�<�N���r� ӯ�������ޯ�Q� @�u�8���\�����ɿ ����ڿ;���_�"� ��Fϧ�j�|��Ϡ�����%���QUIC�C02��!19�2.168.1.10K�@�1��^� ߄��D�2�߮���!�!ROUTER"����!r�I���P�CJOGr�M�!�* t�0{�=�C�AMPRT���!1r�����RT;������`� !Sof�tware Op�erator Panel=�oغ��NAME !3�?!ROBO����S_CFG 1��3� ��Auto-sta�rtedidFTPtoI�o�t�o �����- (:]K���� ��Kn"4F#/Z |:/k/}/�/�/h�/ �/�/�/?0/�/C?U? g?y?�?�?Rodovo�o ?	OP/-O?OQOcOuO <?�O�O�O�O�OO�O _)_;_M___q_�?�? �?�_�O�_$Ooo%o 7o�O[omoo�o�o�_ Ho�o�o�o!3z_ �_�_�_�o��_�� ����o/�A�S�e� w�������я��� �N`rO���s�� ������͟������ '�9�\�]�🁯���� ��ɯ�"�4�F�H�� |�Y�k�}�����h�ſ ׿����0���C�U� g�yϋϝ������� �	�P�-�?�Q�c�u� <ϙ߽߫������߆߀�)�;�M�_�����_?ERR ���o���PDUSIZ � �^�����>��WRD ?����  ?guest�������%�7�I���SC�D_GROUP [3� 
�wIFT��$PA��wOMP�� ���_SH��ED�� �$C��COM��T�TP_AUTH �1��� <!iPendanU��`'!KAR�EL:*`i{�KC���� V�ISION SETy���'?:�^p���������/CTR/L ���I(��
�'FFF�9E3/��FR�S:DEFAUL�Tn,FANU�C Web Server��\!L"/ ����,�/�/??,?�>?}�WR_CON�FIG �~����cn/�ID�L_CPU_PC�� �B����0 ;BH�5MIN�<��~�5GNR_IO�������0HMI_EDIT �~��
 ($IPL�_�"_SMPLG�R3 LOSEIc�on 2B��OO�PEN2Bt7H5s1 FOXO22mO�O$ bktle�ad-inst_�basicpic?k_star^I/ �O�O__;_&___J_��_�_Z!($*uninit�t[�_ �_�_o�_/oo,or_ wo�oto�o�o�o�o�o��o�?$INPT_SIM_DO�6��:NSTAL_oSCRN�6 �Uz�TPMODNTOqLkwT{�!RTYJxp�1Yv3 ENBkw���3OLNK 1���������1�C�U�g��rMAS�TE�0�yH"�qSLAVE ����H D�uSRAMCACHE����5O_CFGǏ�s߃�UO�ۂCMT�@� �2���YCL�Ə��� _ASG s1�s7��
 i� ������ԟ���
� �.�@�R�d�v�q�_�WNUM����
ۂ�IPďևRTRY�_CN(���gq_UQP�����q��� ۂ����</  0�I$3��0@gr?���� ��Dm�plGrp/Sa�r�e_Config.stm��������ѿ�ր���#� 5�G�Y��}Ϗϡϳ� ����f�����1�C� U����ϋߝ߯����� ��t�	��-�?�Q�c� �߇��������p� ���)�;�M�_�q� � ������������~� %7I[m��� ������!3 EWi{
��� �����//A/S/ e/w/�//�/�/�/�/ �/?�/+?=?O?a?s? �??&?�?�?�?�?O O�?9OKO]OoO�O�O "O�O�O�O�O�O_�O �OG_Y_k_}_�_�_0_ �_�_�_�_oo�_Co Uogoyo�o�o,o>o�o �o�o	-�oQc u���:��� ��)���_�q��� ������H�ݏ��� %�7�Ə[�m������ ��D�V�����!�3� E�ԟi�{�������ï�R�K�_MEMBE�RS 2�"�]2� $"����^������RCA_ACC �2���   [}~�� �T�` 6��ps��T�*T��T�g�6z�� �w�i��T���I�BUF001 2�V��= {�u0 _ u0{����U�������곫|���'��2�=�K�U��d�rāĎ�ĜīĹ�Ȫ�������}V!�}����-�ĕ:��J��V��a�}�o��{�ĉ�~{�N�  N�~���0u ~�
Ա�
��
��O  WOz�z	�z��z��!�{)�{��9�{3�A�M��X�f�q�}"괊����ǹ2Կ��������� ���	��������  �%�)�%�1�%�9�%� A�%�I�%�Q�%�Y�%� a�%�i�%�q�%�y�%� ��%��%��%��%� ��%��%��걸��� ���������������� ��������j������u  �����.�FP ��)�� 1��9�:�@��H�M� �X���*�h���q��� B���҉��ґ��ҙ� �ҡ��ҩ��ұ��ҹ�@��������ǹ3�� ����������	�� ���'�.)�7�.9� G�.I�W�.Y�g�. i�w�.y�.�� .�§�.�·�T��� ������������� ���������	�� ���!�/�1�?� T�@�O�N#X�g��� ;p����ҏ���� ����ү���ҿ����+����CFG 2�V� 4T���*�T�T�<�!!��HISѲ�V�� �g� 2025-11-29T�� M;  AGs#�/�/�/R�XT�� `�$h�$pr$x�r$i�#�/??T�[|�pY(8e)?^? p?�?�?�?�?�?�?�?�T���! R�x��Y"1-07-06@A?.O@OROdOR�^%�v �":�$ �$x��/�O�O�MR�X�H5O
__._@_o  T�#X�{/�p_�_�_�_�J▁H2�O�_�_
oo.o@oRoP����O�oR��QgAY"0-08-31�_�o�o�o�o
gAso0BT\f�boP�g2��o���E^��;� �"v fa#oP�&�8�Ӯ7&��C/U/g*bQdy ��G���ɏ�*!d� �� ��� ��� ��i��@ cԏ'�9�'?9?��� ������ɟ۟���� �6�Oh�U�g�y����yH6  [� 8��`� ����@� ��߯��O�OL�9�K�|]�KZ8  ^]P }�h�������ѿ�_�_ ��+�=�O�a�s�ao ���ϗo�o�����|'�x9  _0� [�m��m������8����	 U@ c�p��ɯ:�L�^�L�9$��h�z�g*� qy ��������*�� �� �ⶠ��� �� � ��G�Y�G�Y��ߡ� ����������1 ���2���z���yH��)��@6�� ���lYk}k�� ]P������� ��,/>/P/b/t/�/�/ �ϩ�/����)/?(? :?L?x�/{?�?�?�? �߱��?�?OO�sra �6B�p6B�j?_OqO��Oq�A_I_CF�G 2��� H�
Cycle �TimeqB�usywIdyl�B�Dmin{=QUp�F�A�Read�G�Dow�H�O��Q��CCount�A	ONum �B�C�{�s]pKQY�PROmG�B�������)/softp�art/genl�ink?curr�ent=menu�page,113[3,� s^�Uo�W�631,�P le�_Config.stm�Oo�MJUy��SDT_ISOL�C  ���~���OJ23_DSP_ENB  ^j���`INC ��^kul`A   ?��  =���<�#�
ka�i:�o �a�o�o��o$VxgOB�PC�c�E��f>qG_GROUoP 1�^k��< �tP�a�	�,?��_��! ���(��L�^�p�䂏�6yG_I?N_AUTOKt�i}`POSREF�XvKANJI_M�ASK膯h��RELMON ���|_�yG�`�r�����P���N��S��WՃ��ʕ�քKCL;_L��NUM�`���$KEYLOGG'ING�����*�e��PLANGUAG�E ��f���ENGLIS�H t�|�LG�A١�ZR�'���  ��H  ��� '�7  � +
���� /o=f� ;��
�(�UT1:\��� ��'�9�P�]�o����������ɿ��(�O���HQ�N_DISP ��o X���z�LOCTOLu��Dz�Pga�a���GBOOK ����-��Q��-� �Ԫ������/�A�`Qݑ�Sc�?�	��@ԩ�q9j�߼�Q���_BUFF 2��^k ��%�����>b��G C�ollaborativ �%�7��v� ������������ �E�<�N�{�r�����?DCS ��Y�b �a`ܟ���E'|9��IO 2���� �@n�@�P� r������� $6JZl~ �������/�"/MER_ITM[nd��{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�?���P"SEV��F�.L&TYP[nj/KOp]OoO�=�RST����SCRN_FLW 2�[�P��� �O�O__+_=_O_�O�TP3�[o:B�NGNAM�d��f�6�UPS_ACR�@�ꏾTDIGI�X~IU_LOADCp�G %|Z%ANIMATIO=��ROP\_yeMAXUALRM��Q���e
Bb�Q_PD�U�P ��a�B`CA���͜o������d�dpP 2��� �=�	:O�o+ OaD�p��� ����'�9��]� H���d�v�����ۏƏ ����5� �Y�<�N� ��z�����ן�̟� ��1��&�g�R���v� �������Я	���� ?�*�c�N�����|��� ���Ŀֿ��;�&� _�q�TϕπϹϜϮ� �������7�I�,�m��Xߑ�:hDBGDEF ��e��o���_LDXDISA��P{[KMEMO_{AP�PE ?|[
 ��z��-�?�Q�c�u���B`F�RQ_CFG ���g��A z�@i���|�<��d%��������b��k���*Q�/S� **:\�|�O� a���|և��������� ����2~ߍe[2 `L�p��,(0 �C��(9 ^E�i������ //�6/8jIS�C 1�|YB� � ��~/���ߔ/��/�/��/B/T"_MSTR� �M5SCD 1�
��/c?�/ �?r?�?�?�?�?�?O �?)OOMO8OqO\O�O �O�O�O�O�O�O_�O 7_"_4_m_X_�_|_�_ �_�_�_�_o�_3oo WoBo{ofo�o�o�o�o �o�o�oA,Q wb������ ���=�(�a�L��� p�������ߏʏ���'��K�6�o�?MK����#=�ၟ$M�LTARM���:���� �������METPU���b���+9ND�SP_ADCOLx����CMNT.� !�FNJ�N��FSTLIo�`�0 �#>®���گ|�!�POSCF��=Y�PRPMM����ST,�1�#; 4��#�
^�j�^� n�|�Z�|�~���ҿ�� ƿ����>� �2�t� V�hϪόϞ�����!��SING_CHK�  r�$MODA���\+����տDEV 	��	�MC:N�HSI�ZE��b���TA�SK %��%$�12345678�9 �����TRI�G 1�#; l �����		�J��֣YP�ѣ0��E�M_INF 1��6�`)AT?&FV0E0O����)��E0V1&�A3&B1&D2�&S0&C1S0}=��)ATZ����H�F���:�n���Av���Y��������� ��������� w*��������� �+O� 8J\���/: '/��]//�/h/�/ �/j�/����5? �Y?�/j?�?B/�?n? �?�?�?O�/�/CO�/ ??�O�OP?�O�?�O �O�?_�O?_&_c_u_ (O�_LO^OpO�O�_�O o)o`_Mo _qo,o�o�o�o�oG�NITO�R��G ?b�  � 	EXEC�1f�r2x3x4�x5x��v7x8
x9f�r�Rytr ytryt+ryt7rytCr ytOryt[rytgrytsr�ys2�x2�x2�x2��x2�x2�x2�x2��x2�x2�x3�x3�x3r�R_GRP_SV 1���� (j������~�l�w���oХ�_Djb��ԃ�ION_DB$й|(�b�  �Q�=��+"��b��=��`N ˠ"� }"=�-ud1t�������� �PG_J�OG ���ƫ
�ˠ2��:�o~��=���?�ˠ ����*�ܞD�V�ˡm���n�0�'�ˠ+��@�����ѯ�  ��ѧ�L_N�AME !��� ��!Defa�ult Pers�onality �(from FD�)Y��RMK_E�NONLY�G�R�2�� 1�L��XL� �O�l dm�������ѿ �����+�=�O�a� sυϗϩϻ������� ߥ��$�6�H�Z�l��~ߐߢߴ����� "����#�5�G�Y� k�}���������� ����1�C�U�g�y� ��������������	 -?Qcu�� �����) ;M_q����@���//��<�� ;/M/_/q/�/�/�/�/��/�/�/?��E�a��*/ݟ*?_?��PN?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�Oh?z?�O�O�O __)_;_M___q_�_ �_�_�_�_�_�O�Oo %o7oIo[omoo�o�o �o�o�o�o�o!o�ots���`r}x�d����~���w ��G{���N�A��p .�Y�O�a�s� ������׏-�Ӑ��
���	`C�=�O�a� �3�AD�������[� A�̙(��q*�q��"���tS|���  թtp�pE�C{  &�G�"� k�V�{�����ů�x�qHH�j�p����p+�� � ���� @D�  &)�?�/��?Ā1�ā@I�)���˯�  ;�	lA�	� �X � ����y� ��, � 񈙰����K�o������]K���K]�K	�.���_�Z�����@
��J��Կ���T;f�I���Y�,A�{S��ٽ�>  �3����Ck�j�#3��?2}H���bāO��|S-��π��B����X�畨� kD	�����g  �  ��!ֵ�?��	'�� � ]�I� �  �ٕ��:�È��È�=��͙�-�@�߯�ھ���G���-���N}�+� � 'A��B�I���@�p�Q�V�Czj�Cn�C�� y�~�J1�|�η�{ Nſ A 0ݹB}���|��弝���āDz��$���H�3��X�~�i���������А #4P���ąz��؄�  �p��?��ff������� !�&8j�8ĀN�\
>L����=�ݺ(Ā�P������������q�� xi�;e��m��KZ;��=g;�4�<�<����/����yɐ?fff?���?&;�@==0M?��YH� |�6B�ݹ1��/�� u���	/�-/ /Q/</u/�/r/�/J�zF}��/�/�/? �,?��/_?�/�?n? �?�?�?�?�?O�?%O OIO4OmOXO�˜O�� X�?�OB?_�O_A_ S_e_z_�_&_�_�_@�_�_�_o����3dՙG�Cojoo�o���ؘo�o�o�oH���{�k�}��dD
p,�L�d��`�aUq�I��!n,ȴA2�=q@��T@|�j@$�?��V�^�z�Ð���=#�
>�\)?��
=��G�}�{=�r �,��C+�?�Bp���p}�B6��C7n����?6`���(��5}G��p�Gj��F��}�G�>.E�VD�K�����I2`�F��W�E��'E���D��;�����I+aE��G��cE�vmD��� ��9��ď���ӏ� ��0��@�f�Q���u� ����ҟ������,� �P�;�t�_������� ί���ݯ��:�%� ^�I�[��������ܿ ǿ ���6�!�Z�E� ~�iϢύ��ϱ����� �� ��D�/�h�S�x� �߉��߭�����
��� .��+�d�O��s��@���������p(�q�34�]�����9���!�7��U3~�qmU�g�I�5Q����I�������Q��������=+aO�EP�P��A�O����x����� #\Gl�}�� ����"//��O0�OL/�/p(��/�/ �/�/�/�/�/??C?@1?g?U?w?�?�P2/�?  B�;`p�1KCHpz;`�P@Bo OO+O=OOOaOrM�C�?�O�O�O�O�O�S�?��C�  @�SJ$�P�P�aS�4�U
 �ON_`_ r_�_�_�_�_�_�_�_�oo&o8o�z(Q ���}��'x#�$�MR_CABLE� 2�} ȽtT� �f���o �	�owI�`q�c�ow }�7]1g� �y������ 3�Y��-�c�����u� ����珽�Ϗ��/�U� ��k�1{B��o�� ��˟����������w*A�** qc�OM �~i���[� *[� ���%% 23�45678901�~��� {�����{@��{@�1{@{A
����mnot �sent J�ӣ�W�TEST�FECSALGRO  eg{J�1dC�dQڡ
S�� � {DXbp�n�������� 9UD1:\�maintena�nces.xmlܬ��  +Z��DEFAULT�vLqbGRP 2�^b�  �{@}6�*[V{F  �%�!1st cle�aning of� cont. v��ilationW 56��ڏ�	P����}5+*�}J���ϰ����X�%i�m�echp�cal �check�  �S��@]�d�}5�ϑߣߵ����(�~y�roller;�M�_߭���U�g�y������(�Basi�c quarte�rly���$��,�D��#�5�G�Y� �1M2ߋ�{@"8��N�N���}5�����b�t�C��O��s��������&�(�Overha�u��|�' x{@18}5�ew���{@$V��� �wIT)/;/M/_/q/ ��/��/�/�/? ?%?7?�/[?�/�/�/ �?�?�?�?�?:?�?!O p?O�?iO{O�O�O�O  O�O�O6O_ZO/_A_ S_e_w_�O�_�O�O�_  _�_oo+o=o�_ao �_�_�o�_�o�o�o�o Ro'vo�o]�o� �����<N #�rG�Y�k�}���� �����8���1� C�U���y�ȏڏ쏢� ӟ���	��j�?��� ������������ϯ� ���T���x�M�_�q� ����䯹�˿��>� �%�7�I�[Ϫ��ο ࿵���������!� p�EߔϦ�{��ϟ߱� ������6��Z�l�A� ��e�w��������  �2��V�+�=�O�a� s������������� '9��]���� ��������N #r��k}�� �j�8�\1/ C/U/g/y/��/�/� �/"/�/	??-???�/ c?�/�/�?�/�?�?�? �?OT?)Ox?�?_O�?��O�O�O�O�O@JnB	� X�O__(_lIB IOW_UOWE__�_�_ e_w_�_�_o�_�_7o Io[oo+o�o�o�oso �o�o�o�o�oEW i'9�������| �wA?� ; @nA 5_0� B�T�nF�������lH�*ŏ** F�@ �q�vp������!��E�W�i�{���zOFFߏ��ϟ� 󟵟�)�;�M����� ������������� �Y�k�}��m���� S���ǿٿ�1�C��� 3�E�W�i�+ύϟϱ������WDnA�$M�R_HIST 2���u�� 
 �\B$ 2345?678901�#��Ͽ��9Ozߌ� C�u�O�����߯��� .�@�R�	��i��� c���������*��� N�`����;�����q� ������8��\�n%�nD��SKCFMAP  �u��q����n@��ONREL  nD������EXCFENB��
��FNC�JOGOVL�IM�d�^�K�EY�aj_�PAN�|x�R�UNQa	�SFSPDTYP5< �SIGN��T1MOTS��_CE_GRP7 1��u�� �@r�_/nCL/�/�s/ �/k/�/�/�/?�/? D?�/h??a?�?U?�? �?�?�?�?O.OORO 	O\O�OoO�OcO�O�O�O_�K�QZ_E�DIT���TC�OM_CFG 1�͹e_w_�_ }
FQSI �6+B����_�_��_�o���O@oXT__ARC_��@T_MN_MO�DE��=Z_S�PLco#UAP_�CPL�o$NOCHECK ?�/ � �o /ASew����������N�O_WAIT_L��;W& NTNQ���E�Y�_ERMR0!2й	���� '���Ə؏��_��/�~`O��ю�| ��/aBw?������Z������­+�/A�׈�	<���?��v��� ����_PARAM��ҹ���0o������(� = V�E�W� _�9�����o���ɯۯ`��������C��U��y��cUM_RSPACE�i��Q������$ODRD�SP�c� OFFSET_CAR1P��o�DIS���S;_A~`ARK�<Y�OPEN_FIL�E���Q<VαPT?ION_IOr��s�M_PRG %��%$*�Ͼ�O��WO;��6'���r����:!5�����	�j�	�	 ���	���$d�ϰR�G_DSBL  ��� r�v��R�IENTTO� f�C�� �A �U�`IM_D{�����ϰVӰLCT �c�8RҼ��yd����_PEX�`���RAT�g d� ���UP )���b�; �{���s����$PAL�]��c���_POS�_CH<�&���Ő2�/#�L�XL;���l�j� D�V�h�z��������� ������
.@R@dv����22� ���#5GYk}����� ��//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ k���_�_oo+o=o�Ooaoso�o�o�o��E�a:Ҭ��o�����o	:�P�o3E Wi{����� ����/�A�" w���������я��� ��+�=�O�a�s��� T�f���͟ߟ��� '�9�K�]�o�������ȷ�ɯۮ��;��(��j�dg�8�J� /�m�{���e�������进�
�׷��� 	��9�?�]�����h�ϲ�:�ֵ	`������	���:�o���'�9�K�]�f�A��  t�и_�_���"�x���~���  �����#���C{  ο��ʿ��� #�I�4�m_��Z���OU��D�_�D�H'���� � ����� @D� M ��?�����?���៑C4����s�  ;�	l��	� �X � /�4�%� ��, � �E�J��Hʪ��U򏓤H����Hw�zH��P���������B�  ������������>  �3���C�����c���������B��=������R��f�ek������ծT D�������g  � � ��]����	�'� � 	�I� �  y��Ռ�=���-?��@U[�����[������yN%��  '���C C C��� �*�/�a�`��$�z�� Nq� A 0��B%Ѕ%$�`�%d�l�%��DzV��//�/�/?*?����A2��I2?А 4PI"Z5"��z��^�|���l ??�ff���?�?/? ���?�;��18���?J>LO~ $���(��6EP?HZ9�<�3�7�C1 xޜ�;e�m�B�K�Z;�=g;�4�<<�m��O�?������%Bq�?f7ff?l?&�@���@=0�E?��U�Y$��A����� =_��\_�G!��?�_|_ �_�_�_�_�_�_!o3o oWoio@o�oxo�o(_ J_L_�o�o/S >wbt���� �����H��� �o���o��z������ ��O&�8�ҏk�V��� z���ş��"�ߔ}ق�C�����:�%�?��D�K���o������ %�~�D��د�^��^�]���@I�͞,ȴ�A2=q@��T�@|j@$��?�VT��z��Ð��=#�
�>\)?��
�=�GH����{=@�,��C�+��Bp���[�B6��C7n���?����(��5�G�p�Gj���F�}�G�>�.E�VD�K������I2`��F�W�E���'E���D���;�����I+a�E�G���cE�vmD�����:��7�p�[ϔ� ϸϣ���������� 6�!�Z�E�~�iߢߍ� ���������� ��D� /�T�z�e������ ����
����@�+�d� O���s����������� ��*N9r] o������ �$J5nY�} �����/�4/ /X/C/|/g/�/�/m�=(m�34�]�/mA����%�%�/�/U3�~�m??�"�5qQ-???�"��Y?<k?Q����=�9��?�?�?�?O�<n�P�BP?N^�[�hO�/�tO�O�O�O�I�����O�O_�O_>_)_ b_M_�_q_�_�_�_�_��FP�R��_.oh� 1o;oqo_o�o�o�o�o �o�o�o#Is0y2�_t  B��,���qCH��z�s0@������t�cH�Z�l�~�̐�s3?���=@ @*s35ts0s08�q��[ts5
 �� ����0�B�T�f�x� ��������ҟ�c�ԁ� ��);�'x#��$PARAM_MENU ?�5��  �DEFPU�LSE�	WAITTMOUTH��RCV[� �SHELL_WR�K.$CUR_S�TYLF���OsPT�q��PTB�����C��R_DECSNS�0E�\���!� J�E�W�i����������ڿտ���"��SS�REL_ID  ��5YA�1�USE�_PROG %�,�%σ�2�CCR�_�C�YA4���_HO�ST !,�!���ϐ�TP@���û������0ߏ�_TI�ME]�Cƫ��GDEBUGA�,�2��GINP_FLM3SKY߈�TR�߈�WPGA�� x�7����CH�߇�TYPE)�5���M� v�q��������� ���%�N�I�[�m� ���������������� &!3Eni{���������WO�RD ?	,�
 �	RS���C�PNS�E��:J9Oɡ�BTE�DCOL�E���׭L_� �0�s0����dm�TRACE�CTL 1ׅ5�6� =@ *=@7@��_DT Q؅5 ��D � ]i� ' 	+$
+$+$+$�0-"E+$+$C�-"+$U+$+$+$+!/C�/WA-"��-" Ѐ-"��-"Ȁ-"Ā-"+$*/</N/`/r/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n���#!�%k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w���g������� �����!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O���O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�w��� ������џ����� +�=�O�a�s����������ͯ߯������$PGTRACE�LEN  � � �����3�_UP _����b�j��N�c�3�_CFoG �b�L�*�
c�����������E���  ����w�DEFSPD� ۂ��E���3�H_CONF�IG �b�J�� ��d)��&B� �,�PôƱlH���3�INz�?TRL ނ����8õ]�PE����b���(����3�LID{����	~��LLB 1��_ �I�B8�sB4Ӵ� I��!��LŶ� <<7 �?�K�j� K�b߄߲ߘߺ�����  ����8�f�L�n����4���������M���<�/�A�r���G�RP 1������@A!���4�I��A �C�u�C�OCWjVFx����-�`Ʊ����(�(����0q�C���´B$BE lL6H��l��&�B3�4����`�j4MJ�n ��,����%//  DzJ#S/�� :/{/*/�/�/�/�/�/ �/�/??A?,?>?w?�b?�?�?�?�:)�1�
V7.10be�ta1��+�@��*�@�) @ߺ+A )�?���
?fff>�����1B33�Aж�0
CB(���A���AK���9AD	AVOhOzO(�O�O��p���8�@@>K��@A���??�ff?�@�������Mb��������?� �?�,_>_(_b_L_�_$�1)�l��u)A�Z b��_��_o���1EEl�A�S BڰB�:o�,eBHbc�T���MdI���T��Q��Tx�dxo�o o�o�o�o l���2�� -?s)WM_	t�����KNOW_M � ������SV ��?�Y�i/ �� ��_D�/�A�z�������M����� �B	��6� �I�^��Z����O
�b�T�@ ڱ�1ڰ$� �2����+MR��鯍T�_^+�����~�OADB�ANFWD���S�T��1 1�b���p4EOAT� w/o par!t��B�����=L Q�0�B���f�x����� ���ү�)���,� >�P�b���������ܿ�R��2򜻁4ڿ � �</���3 �+�=�O��4l�~��Ϣ��5�������ς�6�$�6�H��7 e�w߉ߛ��8����X�����MAҐ�����OVLD � �ޏz��P�ARNUM  �����#���SCH]� k�
�������UPD���|^��_CMP_���`����p'ޕv�E�R_CHK�����ޑǂ������RS8q�՟�q_MOҟ���_��
�_RES_G���
ROʽ_ d������� 7*[N`3�@P�5k�� ��7����/7 �/</A/7d�\/{/ �/7�Л/�/�/7
���/�/�/7V 1���fې��@`h����THR_INR�q�bፂޕdm6MA�SSz? Z�7MN�y?�3MON_QU?EUE ���ޖ� �@ 
�N{�U��N�6�8�3END8AIEXE*OE�@�BE)@O�3OP�TIOG(�0PR�OGRAM %��:%�08?���2T�ASK_I_�qNO?CFG ��?���OPDATA���&[`a��2ƅu_ �_�_�_�_h_�_�_o o)o�_Mo_oqo�o6_�INFO���S]� �4?o�o�o $6 HZl~���� ���� �2�D��g�d�S\ nQ��?DIT �_��|��TWERFLKH�`3�CRGADJ ��A���?� ��1��1
P��a��?���z���cQ<@����f%� �r�وn!�MQ2��/��b	H�0lA7�_2<�>����ɻt$�*�/� **:�� ������6�1����;���a�C2[�)� ��9�K�y�o������� ���ۯ�g��#�Q� G�Y�ӿ}�������ſ ?����)��1ϫ�U� gϕϋϝ������� ��	߃�-�?�m�c�u� �ߙ߫�������[�� �E�;�M���q��� ���3�������%� ��I�[�������� ��������w!3a Wi������ O�9/A�e w���X6	"_F/ ۀ4/m/X$㙏/�[/�/W/�/�/���*�SYSTEM�V�9.40107 �27/23/2021 A%݀�
7��#�PREF�_TLA( $G�RID@ES ? $BARcB]2�STYLE]1��~?0OTOENTJ0�  $Po_NAMs0!�0�{2]1z1XY(�J1� � $LIS?T_PORT]2�3wENB�8SRV�0�)�4�6DIREC�T_1�2�42�93��94�95�96�97��98�1  �PF�_HRK0  Q0V�ALUEv�S0O�UPv�$AXI�SzAWC�4� �!$ENABr0� �1G�3%�$CUR��wERA�N�C�Bn0AR�0Y�PoA$TOTA�L_TI�Ar@�CP�WRpBIC1�DRE�GEN�JRpBEXE\A�A$]C�A^1�REe0�EMONT�R_R)Q�2�A_S�x@WWP:SV_LI�M�0tV@�1EGR�E�CG0?PHzBOVsERU0�TV_Hd0�DAYSV�QS_�Y�A$MAXS�IZ9SSUMMA�R�P2 $C�ONFIG_SE�T�CUP�2{ALAf�0RUQ=QC_o6_$CMPR�4 cGDEV�@�P/bI�@�Z c�S]1XBEN�HANCE�A | 
�E*a�@TT�Q'INT�0QM(�^1���_MASKj3P�D_OVRD�3GfE2IX�0JPAXyP�Z5OVCyQ�TBU�qR�YAF5 4� S?e71[o6�P�SLG�P�A \? $PS_�V=p#MO�P^1�AS�0ra3aU<q�fTv��SbtAUx1-p80P>�A (0Q�A�rJvOPCrF�IL_McS�qVE�L:S�0TQLP�3Nt�0.PCPSUL�P�  	$V�{CF�P_�po@�M'�[V1&�V14�2C�U24�3C�34�4C�144��A�0 ��@����0��MINщVGIB1+0��2�*1����3��3��4"��4���@�L��@�@��@̇Ʌ݅ɅP�LUS_TORQ�nA؅����+pSAV�ba	d $�MC_FOLDE>R`	$SLđÑ�se�@M�pIsc��L�OA�`  $��2cΐKEEP__HNADDّ!��R#�CCOMi0�;�{1ڒ=p<�OP  �b�ؑ_0<�xg<�REMS�;��A�2�x�����U�4e;�HPWD  ��SBM�a�0COL�LABLt�@>p�AE:�a�@ITSa��r�$NO�FCA9L(c�CDONrb�q�Ò�a�0
 ,Q0F�LANGoA$SSYNҐI�M�0Cb���@UP_DLYz�1C�DELA{���Ak2YPAD�Q�$TABTP_R��� �QSKIP�:� Ĵ0�POR0k������P_�Pʰ ι�@J��b�}Q���Q ��@��@��+@��8@���E@��R@��9�a�{RA�3 X�P��B�gMBa�NFL�IC�3��REQUx�0�cqwNO_H���r�,`�_SWIT�CH�2RA_PA�RAMG�q ��_0mhUSE_W�J[r
��SscNGR�LT{�O�q$W�ARNWpYp(c�S�T�@J1���rAP�#`WEIGH�3Jg4CH�01�OR�1�1��bOO�@;RAT+IO/�J�@D�0�b�SA��&e�ӓ�OBiO�D^0x0J2����1�bEXD_R{TQTD_IT�C���@0����a�x0R�DC�A=� � ��`�`��R݀��T�H?Q����RGEAFPRIO��8�W�G �`Y�?PER���SsPC���UM_��>�s2TH2N�a����� 1  ����{1�2  �D liX�LVLW2_P���Sgq��QP�L10_CA�q����a  h:q�0��j�0(S���qJ�H��М�Ձ �b񩓁�@�Bb��zA'���`�� }P��DESIG"����1
�1�����;10��_DS�q�|��G0POS11�1 l�B�ZrH��C���ATq����pU��EIND�`�1=� ��=0���HOM]Eg 	2/ASew0�
3����(��4)�;M_q5 ��������6/#/5/G/Y/�k/ 0�7��/�/�/�/�/�/}'8??/?A?S?e?���Sߠ1���QP���`����B T��D�F&CIO�q=II�0bO�_OPIEaC�B؋�� WEӁ# @H��/��D� C��B$DSB?pGNA���v��C��P��S232N#E  �9��5H��3`ICE��SPE����Q��IT�Q qO�PB��RFLOWF�PTR1ТQ��U�S�CUPi�a�UXT��a�Q�`ERFAC�T��U%PS;CHca! t�Ր�_	P`^�$FR?EEFROM�Pvs�Aq�(�A`ۑUPD��)��PT�0&eE�Xذ�X�S!��FA��p2b��@PdPca"�� 塏5�A�L�q�9P�EX`PIHQb�P1PY8e�B_�r0��4aQSfWR�a�?��9DP�wfP��6FR�IEND:�p$�UF��t�`TOO�L�fMYHՐ�bL�ENGTH_VT�E�dI�q�c��$� �`�hUFINV�_ y�ARGI��q6�ITI��gXؕ��g=vG2=gG1�Ga^P��WrhwPRE_�b���D���a�� ���S�cEQӀC��b��q�v
���lS~Q# @.@P�Q꒬zWhpjU�jU���B�|�P�T$X �-M�PCTQcH��YhPP�/U)d�SG��WI`�m�҂�D��a@K�q���ʰ������=$�v 2#�qa� wi1�hr`2uk2
�3uk3�j։-��i��I��60`�0`!�$)V�
rV>uV!�
qQ��q�rP%7�kV ��ߡO��vCR�����b�Z���Ee��	s����5$AG���PR����p�S!�PR�q�"�R&A& �����+�ˀ$�В�ˀ% π�P�p^Pβ
���R�S�A' ؠ�Rp��7A\�/@UNN�@SAX%Q�pA�`L�a�r´�THIC���G���@�^PFERE�NZ���IF_CH�kc��Iug���6��G�1���0$��
pn<�_JFE�PRL�	 �RVW�A~Q(�  $X�;Q ] ^�VALE� ���j�:�)�Bn�  2�( �S,�0*_
  �$�_�� �a��@γT�Ь��γDSP嶫�LILSpE
��A��šȳ���AX��UVK�P_GMIR�!āpMD�&B�AP2� �E/`b�AԶ�SYS8�lB��;PGw�BRK�r�V�NC��I�1  `��vc��в��AD;A<γ;�BSOCٶ3@�N��DUMMY1�66�bSV\�DE�fASFSPD_O�VR��^���LDL��ORצ0N��b�F�֫�OV�CSFTڥ�W��Fp��mA%Ås���alCCH�DLY�RECOQV��pT�W��M��@���������
�_���\� @��,pVE\z@�1OFS,pC���cWD8���4����2,[���TR��	A���E_FDO[�MB�_CMKAF�B BAL��@�hⰑ+�VlQ �R�PY�ƳP�Gi�|�AMz�\��P������_M��NRMŰ9B���T$(���Q�3T$�HBK�Qg��IO�ue�YA��PPA �?�$�O�7���YB��?DVC_DB/s��@h��B����2ј�1������3����ATIEO�@]Q,��Uzc�8FCAB
�tb�s@=����0���QT�_RP~g�SUBCPU���Si��@R��P��Sp���B�$HW_C<P������Akq���$UNI�T��� � ATT�RIj���CYC=L�NECA��L��FLTR_2_F�I��H��F�QLPx�����_SCT�sF_�F_�8�
�FS�A��CHA��a y��CRxRS�D�зB��գ��Y@_T��PRO��@�9PKEM�0_�Ц�Tf�w� f���D�I`i�RAILAiC��4M��LO���c��7�b������V��PR��S�qπ�W!Ct��@	��FUsNC���RIN�p`s�o` w$8QRA� �b �#
@	��#gWAR5���BL�q��'�$A�+��(�(D�A���!8�#�%LD@�PЅ�33汪!ᑆ33TI�S5ɱ���$�PRIA�QRAFD P0�~3�Є5p󀘂��MOI� C�DF_�`�ӸQ;P�LM��FA��HR�DYPdORG80H���ao`0�5MULCSE�`j�S����J�J6�K�F�FAN_ALMLV5S�RAWRNYEHAR�D���V`�p�P� 2�QAQƱ��_��g�A�UmPRkORTO_SBRv�E��J� �v�!�CMPINF���D)1�CRE�GvfNV�P!c��D�A�`R�FL���$M0��RG�ࠠ�`HgUCM�N��Y�#NONI�NE�PpYBjRs&� �I��๱+ ���a]$Aa$Z$q��|����,$ �o��EG�γ��QAR�����23#e� |�wAXE�ROB店RED�W�a��_]m��SY��8a��fS�gWRI��f� �STR䵼@��*�E���d8�AB�`���f9'#��O�TOQ����AR�Y�r!!�����F�I��,�$LINQK�1��'qc�_�c�����3O��`OqX�YZwBYz�jsOFIF��&rNrBxp	B�l"�t���p �sFI� �ww����l"��_J���(Ҡ3s���@�d�j3p�F��TB�qB5�C� &k�DU���32�7"TURT@XZ3n�qb�BX�`���FLm�@��`��pu�i39��
� 1+��K
�Mg�\�54%S�S%�ORQ��# #���␂�1��0�<�pj��#QQ�OVEX���M,0��Sr��Sr� �Rq��@o�p�� o� B�q ,�0��Y�9��� ��0�j�Y�v����S��L���ER��!	8"!E��|�D#9�A瑠��u�%�w11AX�ӆ�1� �(r �����A��ƀ��� ������3 ���`���`��1fp���0���0�� �0���0˩�0۩�0� �0���0��0�8�,�x� �2~�DEBU}$x!�C���JrCAB'�8�R�V�| 
©��/� m;�e�;�Ɓ;��;� ��;�3!;��a;��a�4p:��2ϒ�sLAB�rq�y ��GRO� 4�}L��B_� � �d��p�@������A �ANDڀ8 .� ��Su1��A]� ��Q��`q�1��� RpNT8d@�ӣ�VEL�͔���!���r�0/B�sNA��phbC�T�`s�3#,��b
 �SE�RVE���P- $��p� ��!)�P�OJ�� _�T9P�!�P��1�P. � $M�TRQ"��
L�hbV�/Z�2�2.k�b0 _ �0 lT�AER	R�ra�I���͔��'TOQ͔ʐL<`��(�b���G+�%<q|�� �V`0 1 �,'�o��/ёRA~� 20 d0�rf��b� 2�P�$f���0����L�OC1x�3 � ��COUNT��a n�FZN�_CFGU�4 4� %V�T|�z��ೈ����Z����S5 �,�M�+B�`�pɓo��FAq0ؕ6XX`-	��H�Ga,�� XaPzB��HELAP��6� 5�pB_B;AS|�RSR$V` ERcS<L1� 1�窙 2�
3�
4�
5*�
6�
7�
8���RO�� �-pQpNL��Q@�AB8�
 � A�CK�IN^�T_�UUU�@	@�AL_P�UX�~Be2OU:�P�� %Xy��@�`y�T�PFWD_KAR���-Q��RE7��0P8#p1� QUE$Yf� Y�I���~@�AIU@��yOp���VOqSE�M�q?&E��0AS�TY[SO* P�D�Ig�@��!x��1_�TM9SMANRQܘ&OpENDN�$�KEYSWITCaH��z!$HEI��BEATM�PE�(`LE��� ��(UҾF.$�S$DO/_HOM�0OzAOEF9�PR�q��ja�`UUC
0O�1���OOV_M��pE�pGOCM;�'E��RvzHK�Q7 DLq$&W��U��"M`��K�<�FORC*SW{ARձ��x�OM` 8 @����s�@U�cP`1(FgPD3F4�D���Sc�O�L�29<�%XUNLO���mZDED�A  �P+0��: <NP�1y�}�MSUPGN���ACALC_PLkAN�C1�pAY��a�yC��; � �@9�PA�$�MQ{Aϵ �·`���%Md0��`�r�F�Td��RSC��M�P�ѱ� �<Q����p�OTYWZZWZEU AR㐡PTaՈR�P��Vj�NPX_AS��< 0� ADD|����$SIZeA�$VA���MU/LTIP<�S@�A�1= � A$��P>2�p6bS���aC��"fFRIF�a�^�S�IB4`N=F�$ODBU�`��0#efcai7�CM�!$�ձ������Ƃ�|� !�> � �P���TE��
��$SKGL�aT5r��&����c���`�`STMT<��sPSEG8" q�BWY��dSHOW�ub�BAN�@TP��p���,��7���V+�_G��? �$PC��_�+���kFB�1P�xSP 1Af�un�VD�p��@� ���A00���q@�w@�wP)@�w3@�w5�y6�yU7�y8�y9�yA�y �@�w @�w���v�@�w!F�x+����y1�y�`T���1$�11�1>�U1K�1X�1e�1r�U1�1��1��1���:�x��y2�y2
�2��2$�21�2>�2�K�2X�2e�2r�2��2��2��2��3��y3�y3�y3
�3
�3$�31��H�K�U3X�3e�3r�3�U3��3��3��4�yU4�y4�y4
�4�U4$�41�4>�4K�U4X�4e�4r�4�U4��4��4��5�yU5�y5�y5
�5�U5$�51�5>�5K�U5X�5e�5r�5�U5��5��5��6�yU6�y6�y6
�6�U64�6A�6>�6K�U6h�6e�6r�6�U6��6��6��7�yU7�y7�y7
�7�U74�7A�7>�7K�U7h�7e�7r�7�U7��7��7����VP_UPD�qAs Z��C 
�0�V\b�qB x �$TOR��`  �7SO�� l ��Q_w�RE�r��'��`��S��C1����_�U;`�� ��PYS�LO�C �  �Udb��Qd�W$05�0<�RVALU��q����R�F
�ID_YL�#z�HIu�I�2?$FILE_���Ƶ$?3�p�SA�V�qD h����E_BLCK���q>��D_CPU���P ���Pu������� ��R E � �PW�`.I`XLAqSR��]ngRUN�@G�\��g� ��\�gHВs� g��0T2��_LI�2F � 'G_O:">�P_EDI2�@�T2SPD�G��PIDq`I`
��DCSy Gi�H� � 
$JPC�w�s� SPCOC�^$MDLQ�$u0~TCP�U�F� SCO�B� � ;�r�pI��0M\��O�z�aTABUI�_<�pJ�B< sHD"RI$2#�A�S�`LLB_AVAI2.�P2#��qK $� SEL�� NEs� RG_ N�`�Aq2#SC��0L �o!Bb@TB�q� _M�@��pM \��PFo1LI_���&M�b-@G�p�Uy2]t6:rPS_JXbP�` �P,5Ew"��TBC2�EN a��`�@�@�B$��FT@qag4"PZ�TDC�e� �0�P;c�5&{7THX`�1�4��ڴ7R�$�PERVEn3�4{3�4�aF2�_AC�0 OX -$A�@n3D�{3@� PI`aPL�OW�'F1A��2�HG*P��`3C\`ERTIA5T��pI��@�KDE�EXaLAC�EM��CCcC��V�2�P�F�E�G�ATCqV�L�A�GTRQ�L UZ�r�C�q:U�C�q!JQ��QZ�Ja��pR�E�Q�EA2�`9p*!@�C�0JK�VVK|q�Q�1�Q�a�P�Jpq�Q�SJJ�SJJ�SAAL�S�P�S��P�V�a�R5�3)PN�1\)`�K�@uD�!_�qq`]�H0CF�"P{ `��GROU`�(�aZB�qN^0CpS�`?REQUIR�2>�GEBU3�1�� 2O�a�0�fG1�SGL5Q�  A�PPRPCw ��
u$� N�hCLO-�yS�5y�E~ BC�� AR �d0M��0�@P�2Wt_MG��apC�p��kx�0�lwBRKjyNOL�DjvSHORTM!O��z�}[uJ�!3CP�T�@�S�@�S�@c��@c�@#1�r7�u8�1{��1M4S� �b(Bn1G��1U�PATHQ�j�`�j��-Hf�Gp�`R��NT¼ A%�w�b`qINF BUCt@[A��C?PKUMɈYJ@��iP Ё~��1늣0��P뀿PAYLOA�wJ;2Lf�R_A� *��LY 6�2�&�B�kuR_F2LSHR�4o�LO7���p�̓~�̓ACR����������2HS�uB$H�krޒFLEX�cuXG0JK6T P�b�\?n?�?�?��� EU :OF�@p����"O�1�@+O=OOLF1��ե�^OpO�O�O�O�O�E�O�O�O�O 
__._@_R_��TW ��T���s_�_�_���ZTa��X�����U \�D��U�ŗ��_�_�_ �P�Ue�Ueo1oCotUibbJhdV �W0`uo�o�oZ�g�AT��a^PELp��"�ҳh�J�`U�`JE�pCTRw"��N���֤gHAND_VB�Q��_�M4W� Q@4kv�4M�SW��D3�EvX� $$M T�Xy���q��q�쳰��r��A��#�[v��D��d}Au|C��zA�{AA�{��v{ �zD�{�D�{P��Go m�S�T�wu�yu�N�xDY� �`kv����4�@ f���f���%��WDį����uP�u�u�
����%�.��[�M4Yc w�\�O� *�xs)qASYM��P`�`��XR`������_SH\b��؄�}��H�����*�J�1��pC�cYb��_�VI+��)s�V_UNI�3���n�J�U������� �&��^P���pß՟Df%����D2E�p�CHh Z ���dO�TO��P�PD�V�3�$�5��R��P�q��Xq� �$�!� _u����0�%�!�����PROG_NA��$Tj$LAS9T�qR�CAN���3~� XYZ_SP��@�$X7�� �l6S� �05q1EN�p14CU�R�(�0�`HR_TF�b[A�1y3N���pS�O�4 ����1�\ ����I�A�$�� A��C�����0s��0 ]o � Y�MEX����)Bc"�T�0P�TFe�q�QAU`Yd �(VHqAeITGZa� $DUMM�Y1��$PS_6 �RF   q��F��FLAj`YP�R��BYC$GLB_T���5�EQ@���wLIFh^�E���f�@OW+@O�UV�OLY�� 0Q_2Ɂ�D2.��@�pP�6R��00S�@TC�$�BAUD��SST�6�B��@ARIT�YpSD_WA�TAeIUYC��r�OUv���Q�YTLANS��@�[��SZ\C'�BUF_�RL����X�0޹YCHK_0CE�Sɡ��JOG@E��AQ!4hRUBYT:�KiH�Kd�rn�nf@`�Q��!��fH��>���1_ X
���a�STY���SBR�U M21_� ��T?$SV_ERR�e��cCL�@�bAq�Ol�"�0GL�EWh�` 4 $[A�$�Q$�Q$W 3sy��!U�#0Rɂ�@:sUua b�"4�$GI�}$�q  psLphb� L$pnv}$FzEvvNEARR�N?2$F�yO�TG1�Z/�J0R�� �cw�$JOIN�T���uMSET.hd  kwE�ur��S��t��he��  ��UX�?����LOCK_FOx��`��0BGLV��GLg�TE:0XM��&�EMP�p��8���BR�$UP�rF{ 2a��Ls��b|�h\�W���`�aCEo�|sҀ $KAR��}M�3TPDRAp��qVEC�� ��pkIU��c��HEY�OTOOLɣ%�VȤ;RE�IS3H�E��6/��!CH�� d&�1ONWE�D3Wc;��I�"6P@$RAI�L_BOXE{!���ROB0��?�~�aHOWWARp!x���@m�ROLM�B Ǖd�j�ؒ��6P�;�O_F��!��HTML5x1K3��P� ��� r_�hf�~^ � W�hg�r���q��qv�Phh t�Ђ��`NA�Ҵ�R���P�O[�1IS0��N P�;���_����2��!ORDEDW�� Q�&�pXT��%1)�3���O@ i D �@OB���W� ��C�@���SYS�ADR�Ѱ0Q@|� �� j ,b�NV$A^�!5\�|=5%APVWVA,A?k � 0r��5PR�"$E�DI1��VSHWeR������IS�p�Q`ND;@wcس�cHEAD+` �;���KE�Q�@CP\i0�JMP�L�5� PRACE�4l���Q�I��S��C�%�NE.����TISCK/��M�1�1�2�HN�am @(��O��7C7�P�6����@STY�"k�LO��Ad�2�ns�
L0 6%$��"4=��SW�!$�{ @A��Ea�EP� �6SQ�U�RLO�B�T�ERCU@ZC�T=S�o up�`@�׭ s����N�OV@�ICU IZ�D"1�E@�A%a�B���A�PP�RN��_DO?2[�X�P9S�1�3AXI�Q�!���3E� T����P�REQ_�,�E�T-�*P33���Fd���A���D�9BX�0 VrSRdplmз���@�s��
����VJ1��h���A���q��@��A8���I���� ���D+��P?���C��,�C=�%7I��pTSSC�@ 7q h�DS����f�@SP� AT*��J2�ь�[BAD�DR)c$�P� IyF3��_2CH+��/`O���m �TU��`I�� r�rC�U�PN��XpV<�I��2sM�t�.�C�
�
C�� ���0t 	\�`��������@0�C^��Q��
���b���TXSCRE�E�u�0_P��IN!As|pL"4� F�sQ_.Pv TA� �`�B,��a�����+��ҕ��RRB`�q+����D�1UE7�w# ���!a�@Sq,�'RSM����U۠W��6!�0S_Fs#&�� !&)A'��.�CL��ހ 2vGUE���x�2�bf&1M_TN_FLj��1��`���q��BBL_ro�W�@�0y ���j�"O@q�"LE^��#����$RIGH�TRD�dTCKG�R�@5Tܠ
71WIDTHBSͰB����A+b �UI��E9Y���z d$p
��Ɛ��6P��BAC�K���B~5q4@F�Oɡ�7LAB��?�(4@I-�P�$UAR���0pW0:@H�� { 8 $��0T_�l�2;@R��PR�GSu��A^��1O�e�`|��w�PU�� /CR`�ґLUM8/C�N ERV���3�P�p^4} � b�GE�2�qY��ﰓLP�EW�ET���)��G��H��HY��I5
�K6�K7�KMP�@R� �Ӹ��pDU1Y�=`�A |V1US=Rt~ <�`�01Urr�rrFO� rrPRIj�my��рP�TRIP��m�oUNDO6�ip�ЙP�չ����8��+�` ��2KP.$aG ��T���Lm�ROSr��VR1���S+��!�"4s;~$b��U0��U�A�!��o.o<#�B���SOSFF��� � Dc�O�`�����d�d��GU&�P�a\��c����gk1SUB�� }��E_EXE6��V���SWO�� e�c`�W�WA���KPq��J V_CDB-sEpC�KPT`䅖��q��;#OR�o�uuRAUD vtTȋyD�[q_��7��s |��D�OWN��>s$SRC��0��D���u��MPFqI����-�ESP�� ��d=�^CޱZGK�Ra8�r���� `e`rrs��2�COP�$���P_�px�o�k�v�7rCT3q)��qK���DCSŐP�L��4 COM\P�Q�{�xҏ���}�HcCq�a��o��VT�Qg`�bY�Zޱr`K�F�� ���SB$�>�r����_�M*�e��DI�C_�AY���P�EE0T�1��VR�q������ �0C�� <�����W��� ~ Gg5�vs�!������ ��SHAD�OW�Q
�_UNgSCA���OW����DGDE_LE�GACi�� �V�C��C\c�� A��%������R��w�0�w�@Cr@w�D�RIV��8��C��!��h�� ܂ MY_UBY+T���c ��1�d)��0�̱�_ ���&�L��BMv�!$Z�DEYI�cEX� ��o�MU&�1X=�l� US*��{P_RbC�pPc���D�G_�PACINj��RG�q����zc`��9c��K#o�RE�2�ba\�\���� �S � a�G��P/H����]�R`� �f0�(@�L1�b	n���RmE=�SW��_A����`k���OAQ-1A(o�s¨�E��U��ϒg ��]�HK���%@��EП�o����EAN��prprż�P]�MRCV�!�; �z@ORG�Б�	Ҍc���REF�'$����a�k@[� I�PP�Z��Z�)�|�ֱ�_�p�ʲ�����SP��ˣڅeA]��$� ��?�Q\Q�Х�OU�؛� g����2�� 0Mq�jP�-���F� N UL_ �f.�CO�i��\�Y�NT)��䩂��A��8Q��e�L)���0����A��8Q�VI�Av� �pHD<w v0$JOP�"��$Z_UP|���Z_LOW5���d��1�"���$EPY��S�Y%��@�G\FG �q���o 5-PA81{ -CACHf�LONѷ���]���C1T���C��I_F�����T������$HO�rps��Á���O � 3�L2���q}A���VP����_SIZf��Zd��5�؇7q3MP�
FA�I��GV���AD�	o�MRE����GP R��py�AS�YNBUF�RT�D-9�3OLEO_2D_tcUW9c$����UK���Q���ECCU�VEM�հ�����VIRC �M5�9_~�jX�P�P�AGIR_�GXYZE -#_�W/� (L�$k1�Tb�L��IM�L�C0��G�RABBa<�{�L�ER��CN�{�F_1D(���.V50�()���%B���Y���2LAS902ћ�_;GE��� ����q�O�%T���b�/��9R�I4����B�G_LEV�1��PaK����Q�GI� N�0t�p�"����Hk��P��S� ��N�4O��VL
q�����σcAO�*SbD�QDEY��q�8��8B�W�C�����p�b�WPA�:ڄ0T8S��Q�MDtQ� ��rPTĂ�Ufq� $&qIT��RyP�1���bVsSFd���  �P�o���_�URf���S�M�U��R�xAD�J]@���ZD�F�3 DHV�AL?�� �t U�PERI�"�$MSG_QM�$���`7r��gp���RzG�Q^�cG �X�VR�T��"�PT_����2 �ZABCBbu�RڃC�
����AACTVSg� � � $�U<3 
SCTIV�1G�IO���SB��ITlU���DV�
���Y0�p��q `P	Sݑ�r ��rGސaGLST��G���M�\f_S�� ��R��CH�r� Lmq�c�U���j�8D��А GNAET`x��G��_FUN?��G ��ZIP�t�LTRQ�$LˢA��!_ZMPCFbu��B�p�R�qڡLNK�0�
Cq ct�� $@��tCWMCM��Cx�Cb��Zq0�P�Q $JxsrtDv~r�r �w���u��rw�ԍr��wUX!uUXE q��v!�u�u�u�q�qp�y�q�wpFTF��~s8�2���Z�eG� �K�dY�	Q��Y^�Dg  � �8��R� U�$�HEIGH��zH?(a�gVB�%�R��� � �D/ѱP�$Be�����SH�IF�HRV��FPC����PC�srhq x�@���3p�#9�kYDI�b`CE�PV��}�Q�SPHER�� � ,a�����6���y@GNp�)�ޏP�����W�X@X@
X@� ��IORITYy Y���ʒ���$`SP�@�P品���֓��;��r
@ ʒגODU��&x�����W�5�G�GL�H�1��HIBHQO���T�OE�1D� � (!AF��E� �ӯާ!tc�pޯ�!ud���.�!icm��V�5�XY�� ��� �ԑ)�� *������X@���Ϳ�������� ��S�:�w�^ϛϭ� ���ϸ����*4�p�	���%+�=�O�a�� >�M#c�z	�/�� **:���9߮�����ض��A��,  �ΐ����*��`���Z��m�������ENHAN�CE (���A�>�d�����  ��1�����ѓ�P���QkR�X@����RTREPx�w�g�SKST�`�㖡�SLGu ������ԑUnothing� ���� ��CUg�Y���TEMP �D�xz�4 _a_seiban�	Š����2 VAzew�� ����//@/R/ =/v/a/�/�/�/�/�/ �/�/??<?'?`?K? �?o?�?�?�?�?�?O �?&OOJO5OGO�OkO �O�O�O�O�O�O_"_ _F_1_j_U_�_y_�_�_�_�_��VERS�׀A�` d?isable��]SAVE 	D��	2670H7K00�X�_po!��0ro�o/��o 	�h*�H|��o�e�o�e ;M_qz*|�op�9�/gƁ 1
��]`�p'��5����'���URGh�Bu���h�WFA���䔄��/�W̠b�K�f�W�RUP_DELA�Y ����_?HOT %3�,�����s�R_NORMALňL�Տ*���SEMI	�/�n�֑_QSKIP�s3��sx�_���_ן��� ��3�"�0��P�b�t� :�������ί�򯸯 ��:�L�^�$�n��� ����ʿܿ�� ��� 6�H�Z� �~�lϢϴ� �ό������� �2�D��3��$RACFG� ����|��~b�_PARAM���3�� @��s@`��|�2C��5�|���Cg�G�=Bb�BTIF����~b�CVTMOU������b�DCR��s�� ��ʑ=t�B8�*B(^P@����@-�S;���������}վ-��T3�
�x̟���;e�m����KZ;�=g;�4�<<���pJ���� � :�L�^�p���������������� }�RDI�O_TYPE  �7��u��
EDPR�OT_f���,C�|�BHg�E��Xv��2h ���B��Я�
����� �+�\[�� ��ߴ���� "//F/T'rw/��>/ �/�/�/�/�/�/�/�/ ?B?d/i?�/�?$?�? �?�?�?�?O�?,ON? SOr?$O�O O�O�O�O �O�O_�O(_JOO_nO 0_
_p_�_�_�_�_�_ �_o4_9oKo
oloo �o~o�o�o�o�o�o 0o5TohV�z �����@1����XINT 2�ȉ��q�G;� �o�����祐j�f�0 Ǐً����	� ��S�A�w�]����� ��џ����۟�+�� O�=�s���k�����ͯ �����'��K�9� o���g�����ɿ��ٿ����#��G�T�EFPOS1 1'	?  x��� t���ϩ����ȈϚ� ��5� �Y���}�ߡ� <ߞ���r��ߖ��� C�U����<����� \����	����?��� c����"�����X�j� ����)��M��q n�B�f�� %��mX� ,�P�t�/� 3/�W/�{/�/(/:/ t/�/�/�/�/?�/A? �/>?w??�?6?�?Z? �?�?�?�?�?=O(OaO �?�O O�ODO�O�OzO _�O'_�OK_]_�O
_ D_�_�_�_d_�_�_o �_oGo�_koo�o*o �o�o`oro�o�o1 �oU�oyv�J �n���-��� �u�`���4���X�� |�ޏ���;�֏_��� ����0�B�|�ݟȟ� ��%���I��F���k�2 1w�!�3� m��֯��3�ίW� �T���(���L�տp� ���������S�>�w� ϛ�6Ͽ�Zϼ��ϐ� ߴ�=���a���� � Z߻ߦ���z���'� ��$�]��߁���@� ��d�v����#��G� ��k����*�����`� ������1������ *�v�J�n� ��-�Q�u �4FX���/ �;/�_/�\/�/0/ �/T/�/x/?�/�/�/ �/[?F???�?>?�? b?�?�?�?!O�?EO�? iOOO(ObO�O�O�O �O_�O/_�O,_e_ _ �_$_�_H_�_l_~_�_ �_+ooOo�_soo�o 2o�o�oho�o�o�o 9�o�o�o2�~� R�v���5���Y��}��������3 1��N�`���� �<�B�`�������� ��U�ޟy����&��� ӟ����k���?�ȯ c�쯇��"���F�� j����)�;�M���� ӿϧ�0�˿T��Q� ��%Ϯ�I���m��ϑ� �ϵ���P�;�t�ߘ� 3߼�W߹��ߍ��� :���^�����W�� ����w� ���$���!� Z���~����=���a� s����� D��h �'��]�� 
�.���'� s�G�k��� */�N/�r//�/1/ C/U/�/�/�/?�/8? �/\?�/Y?�?-?�?Q? �?u?�?�?�?�?�?XO CO|OO�O;O�O_O�O �O�O_�OB_�Of__ _%___�_�_�__o �_,o�_)obo�_�o!o�oEo�o��Ƅ4 1я{o�o�oE0i oo�(�L��� ��/��S�� �� L�����яl������ ���O��s����2� ��V�h�z���� �9� ԟ]������~���R� ۯv�����#���Я� �}�h���<�ſ`�� ���Ϻ�C�޿g�� ��&�8�Jτ�����	� ��-���Q���N߇�"� ��F���j��ߎߠ߲� ��M�8�q���0�� T��������7��� [�����T������� t�����!��W�� {�:�^p� �A�e � $��Z�~/� +/���$/�/p/�/ D/�/h/�/�/�/'?�/ K?�/o?
?�?.?@?R? �?�?�?O�?5O�?YO �?VO�O*O�ONO�OrOx�O�o�d5 1�o �O�O�Or_]_�_�O�_ U_�_y_�_o�_8o�_ \o�_�oo-o?oyo�o �o�o�o"�oF�oC |�;�_�� ���B�-�f���� %���I�������� ,�ǏP�����I��� ��Οi�򟍟���� L��p����/���S� e�w������6�ѯZ� ��~��{���O�ؿs� ���� ϻ�Ϳ߿�z� eϞ�9���]��ρ��� ߷�@���d��ψ�#� 5�G߁�������*� ��N���K����C� ��g��������J� 5�n�	���-���Q��� ������4��X�� Q���q� ��T�x �7�[m�/ />/�b/��/!/�/ �/W/�/{/?�/(?_ T6 1+_�/�/ !?�?�?�?�/�?�?O �?OAO�?eO O�O$O �OHOZOlO�O_�O+_ �OO_�Os__p_�_D_ �_h_�_�_o�_�_�_ oooZo�o.o�oRo�o vo�o�o5�oY�o }*<v��� ���C��@�y�� ��8���\�叀����� ޏ?�*�c�����"��� F����|����)�ğ M�����F�����˯ f�﯊�����I�� m����,���P�b�t� �����3�οW��{� �xϱ�L���p��ϔ� ߸������w�bߛ� 6߿�Z���~����� =���a��߅� �2�D� ~��������'���K� ��H������@���d� ����������G2k �*�N�����1�U;?M47 1X?N� ���/�8/�5/ n/	/�/-/�/Q/�/u/ �/�/�/4??X?�/|? ?�?;?�?�?q?�?�? O�?BO�?�?O;O�O �O�O[O�OO_�O_ >_�Ob_�O�_!_�_E_ W_i_�_o�_(o�_Lo �_poomo�oAo�oeo �o�o�o�o�ol W�+�O�s� ��2��V��z�� '�9�s�ԏ������� ��@�ۏ=�v����5� ��Y��}�����۟<� '�`��������C��� ޯy����&���J�� ��	�C�����ȿc�� ��ϫ��F��j�� ��)ϲ�M�_�qϫ�� ��0���T���x��u� ��I���m��ߑ��� �����t�_��3�� W���{������:����^����hz8 1�/�A�{����� #�A��e b�6 �Z�~���  aL� �D� h�/�'/�K/� o/
//./h/�/�/�/ �/?�/5?�/2?k?? �?*?�?N?�?r?�?�? �?1OOUO�?yOO�O 8O�O�OnO�O�O_�O ?_�O�O�O8_�_�_�_ X_�_|_o�_o;o�_ _o�_�oo�oBoTofo �o�o%�oI�om j�>�b�� �����i�T��� (���L�Տp�ҏ��� /�ʏS��w��$�6� p�џ���������=� ؟:�s����2���V� ߯z�����د9�$�]� �������@���ۿv� ����#Ͼ�G����� @ϡό���`��τ�� ��
�C���g�ߋ�&���ߕ���MASK +1�������~��XNO  ��� ��MOTE  �"��X�_CFG _��Tԓ��PL_RANG[��WѶ����OWER� �����S�M_DRYPRG7 %���%\�����TART ����UME_PR�O����v���_EX�EC_ENB  y���GSPDO������TDB̴���RM����IN�GVERSION� #�e���I_AIRPUR��� W�0�l��MTE_��T��]�����OBOT_ISO�LC ��h ���^�NAME�-���OB_CATEG ���1�$�8@�ORD_NUM� ?��e�H700  �T�{����PC_TIMEOUT��{ x��S232x��1 #��� L�TEACH PENDAN�tד�$[�Y����� ����� ce Cons�T�/-&"'/U�?мֳ e-W/�/K�No Us��/�/�/�NPO�)��������CH_LR�!̙��	F1?!OUD1:l??R�ЏVAIL\�T �����PACE1� 2"#�
@?���,zӑ��U |i)L< ��0?��;PO�?0O�O�O ~O�O�G�?�?OO�O >O`OV_w_6_�_�_�] #�#��]�O�O__�_ B_d_Zo{o:o�o�o�o �o�O�_oo,o�oPo roh�o�����o �o(�Lnd� ��D�������Џ� � �$�6�H�Z�|�r�@� ����ɟ������ � 2��V�x�n���N��� ů��گ��
��.�� R�d�j���J������� ������*�<��`� ��xϙ�HϺ��϶��� ��&�8���\ώ�t� ��Tߪ��ߢ���;�12�<� �?�*� <���`ߒߕ���u���������3�'�9� K�]��������� ����"#�46�H� Z�l�~�0�����@�.CD5W i{��Q����>�./O/&/d/e6 x����r/�/ ?_/�/O?p?G?�?�/7�/�/�/�/�/�?? 7?:O�?OpO�OhO�O�?8�?�?�?�?O�O &OXO[_�O;_�_�_�_��_�OG &�K� �_�
(` o  �EHoZolo ~o�o�o�o�CX�m_ �_�o�_2�dHp-o ?om����� �o�o�n�z!�3�P�C U�������ˏݏ� ��	��=�O�p�c� u�����ǟٟ�������)�;�]�o� `�_ @Ш� ����������� ������*�l�~��� R���ƿؿ������� 2�����JόϞϼ� rϤ�����������߈R��"�
֯���_MODE  �I�R��S '�K��L�J�/_ү��M��r�	m��+�CWO�RK_AD�������-�R  ��K�@������_I�NTVAL��T���C��OPTION�� �N V_�DATA_GRPg 2)(��AD��P��o���~����� ��������,< >P�t���� ��(L:p ^������� / /6/$/Z/H/j/�/ ~/�/�/�/�/�/�/? ? ?V?D?z?h?�?�? �?�?�?�?�?O
O@O .OdOROtOvO�O�O�O �O�O_�O*__:_`_�N_�_���$SAF�_DO_PULS�����o�c�Q�PCAN_TIM�ў�0���QR *D��E�^��&`&b,��A�cK��Q�� ��6oHoZolo~o�o o�o�o�o�o�o�+o��b27t�Q"�QdCx:qJq���Sy���������fyz \��t��w_ ��  T�����#�5�B�T D��B�k�}����� ��ŏ׏�����1� C�U�g�y����&�xz��ڟ쟱��  @�;��o��
�K�p���
�t��Dik�|a7�  � ��b ��e�Q��F������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ�������@��� �2�D�N��� r߄ߖߨߺ������� �Q�%u.�@�R�d�v� �����������0�r\�S�h���!� 3�E�W�i�{������� ��������/A Sew����� ��+=Oa s������� \�/'/9/K/]/o/�/ �/�/�/"��/�/�/? #?5?G?Y?k?���� �b�?�?�?�?�?OO )O;OMO_OqOI�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTofoxoM�衟Q��o�o �o�o�o,>P bt��������z�o�$�.�����2��	12345678s��h!B!ܯ� 
F��` ��������ʏ܏� � �$�*��oM�_�q��� ������˟ݟ��� %�7�I�[�m�~�<��� ��ůׯ�����1� C�U�g�y��������� ������	��-�?�Q� c�uχϙϫϽ����� ����ֿ;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m�,ߑ� ������������!� 3�E�W�i�{������� ��������/A Sew����� ����=Oa s������� //'/9/K/]/o/. �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�?�?�?����?�?�5��/O1OCO_�Cz�  A��j   ���h2�}� >OF
�G_�  	��2�? �O�O�O�O\�oL��OR_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o7_�o �o�o&8J\ n������� ��"�4�B�A�A:�B<_� U��A?  �o����sCu@l��A�At C v@��ŏ�@(ۃ `Rl����iMu@�0\�$SCR_G�RP 1,E+�E4� �{ ��B |E�	 `��h�y�r��^�~E����������ڟRM3��@גD�#\���כ0\CR�X-10iA 0�12345678+90�@N� \��@�N�0 k��A
�X���	���K ��h��W���W�0SD^�בv�����	�����*�<�N�^����H����l� W�������ſ׿���o�A��Ϯ�?�XG0��w�\Ch_@,[}x�x  �䄑B�  BƊψ¡Ą�9Av@��  @�@��愑@����� ?���Ǆ�H��߳ʄ�F?@ F�`+�3� *�W�B�{�fߋ߱ߜ� �����ߤ�������$�0�!�3�E�B�S��� ������������ �;�&�_�J�����/^ �ß����|G�@��D@I���e@nM B�bX� �����?�TA����H���� 0Q��A ���/��DPb1 	(�@�(���� {��� /)L�����='£�7�ECL�VL  Q   ���Ǣ� Q@P!L�_DEFAULT|X$L!��@�l#HOTSTR�x-��"MIPOW�ERFW ZE�%ޮ$WFDOy& ��%6�ERVENT� 1-_!_!�# �L!DUM_E�IP/8�j!?AF_INEx =?�T!FT?l>�3?�?!���? ��?�?!RPC_OMAIN�?�8��?�(O�3VIS�?�9��OtO!OPCU�AuO�JcO�O!7TP�@PU�O&9�d�O_!
PMON_PROXY_�)6e�OX_�B&_"=f�G_�_!RDM_'SRV�_&9g�_�_G!R��o'8h�_�<o!
�0Mo_#<i�+o�o!RLSY3NC�o�i8wo�o�!ROS?�l�y4�o !
CE�@�MTCOM!)6k�l!	5rCON�Sm(7l[�!>5rWASRC�_)6�m��!5rUS�B�'8n�P�!GSTM� j�%:o?�����?���S����#I�CE_KL ?%��+ (%SVCPRG1�1��21�6� �3Y�^� �4���� �5���� �6џ֟ �7���� �Hy�A�<�9I�N�� ov� �#��� �K�Ư  �s�� ���� �ß >� ��f� ���� � ;��� �c�޿H���� H���.�H�ܯV�H�� ~�H�,���H�T���H� |���H����H�̿F� H���n�p��� � � ������@��&�� J�5�n�Y��}���� ���������4��X� C�j���y��������� ����0T?x c������� >)bM�� �����/�(/�/:/^/I/�/�_D�EV �)��UT1:�'4����$GRP 2�1�%� �bx 	� 
 ,� �/?�"�/.??R? 9?K?�?o?�?�?�?�? �?O�?*O<O#O`OGO �O�O�/�OqO�O�O�O _�O8_J_1_n_U_�_ y_�_�_�_�_�_o"o 	oFo�O;o|o3o�o�o �o�o�o�o�o0 T;x�q��� ���_o,�>�%�b� I���m��������Ǐ ����:�!�^�p�W� ��{���ʟ!��� $��H�/�l�~�e��� ��Ư������� �� D�V�=�z�џo���g� Կ����
��.��R� d�Kψ�oϬϾϥ��� �������<ߓ�`�r� Yߖ�}ߺߡ߳����� ���8�J�1�n�U�� ����������U�"� ��F�X�?�|�c����� ������������0 T;x�q��� ���,>%b I������ �/�:/!/3/p/�#d Խ&	^/�/�/��/�/�/�/?";%�x"?G?�#���`1 1`5p?~7h?�?�?�? �?�?�94?O\9�?FO 4OjOXOzO|O�O�OO �O*O�O__B_0_f_ T_v_�O�O�__�_�_ �_oo>o,obo�_�o �_Ro�oNo�o�o�o :|oa�o*�� ������T9� x�l�Z���~����� ď�,��P�ڏD�2� h�V���z����ן� ����
�@�.�d�R� ��ʟ���x��Я� ���<�*�`�����Ư P�����޿̿��� 8�z�_Ϟ�(ϒπ϶� ��������@�f�7�v� �j�Xߎ�|߲ߠ��� ���<���0���@�f� T��x�������� ���,��<�b�P��� �����v������� (8^�����N ���� �$f K]6~�� ���>#/b�V/ D/f/h/z/�/�/�// �/:/�/.??R?@?b? d?v?�?�/�??�?O �?*OONO<O^O�?�? �O�?�O�O�O_�O&_ _J_�Oq_�O:_�_6_ �_�_�_�_�_"od_Io �_o|ojo�o�o�o�o �o�o<o!`o�oTB xf����� 8�,��P�>�t�b� �����я������� (��L�:�p�����֏ `�ʟ��ڟܟ�$�� H���o���8�����Ư ��֯د� �b�G��� �z�h�����¿��ҿ (�N��^���R�@�v� dϚψϾ� ���$Ϯ� ߪ�(�N�<�r�`ߖ� �Ͻ��φ������� $�J�8�n�ߕ���^� ���������� �F� ��m���6��������� ����N�3E�� ��f�����& J�>,NPb �����"�/ /:/(/J/L/^/�/� �/��/�/�/? ?6? $?F?�/�/�?�/l?�? �?�?�?O�?2Ot?YO �?"O�OO�O�O�O�O �O
_LO1_pO�Od_R_ �_v_�_�_�_�_$_	o H_�_<o*o`oNo�oro �o�o�_�o o�o 8&\J��o�� p�l���4�"� X����H����� ď֏���0�r�W���  ���x���������ҟ �J�/�n���b�P��� t��������6��F� �:�(�^�L���p��� �Ϳ��� ϒ��6� $�Z�H�~������n� ���������2� �V� ��}߼�F߰ߞ����� �����.�p�U��� ��v��������6� �-������N���r� ���������2���& 68J�n��� �
���"2 4F|���l� ���//./�� {/�T/�/�/�/�/�/ �/?\/A?�/
?t?? �?�?�?�?�?�?4?O X?�?LO:OpO^O�O�O �O�OO�O0O�O$__ H_6_l_Z_|_�_�O�_ _�_�_�_ ooDo2o ho�_�o�oXozoTo�o �o�o
@�og�o 0������� �Z?�~�r�`��� ����������2��V� ��J�8�n�\������� ����.�ȟ"��F� 4�j�X���П����~� �z�����B�0�f� ����̯V������ҿ ����>π�eϤ�.� �φϼϪ�������� X�=�|��p�^ߔ߂� �ߦ���������� ��6�l�Z��~���� �������� �2� h�V��������|��� ��
��.d�� ���T���� �l�c�<� �����/D)/ h�\/�l/�/�/�/ �/�//?@/�/4?"? X?F?h?�?|?�?�/�? ?�?O�?0OOTOBO dO�O�?�O�?zO�O�O _�O,__P_�Ow_�_ @_b_<_�_�_�_o�_ (oj_Oo�_o�opo�o �o�o�o�o Bo'fo �oZH~l��� ��>�2� �V� D�z�h�����׏� ��
���.��R�@�v� ����܏f�Пb���� ��*��N���u���>� ����̯��ܯ��&� h�M������n����� ȿ��ؿ��@�%�d�� X�F�|�jϠώ���� ���ϴ��ϰ��T�B� x�fߜ�����ߌ��� �����P�>�t�� ����d��������� ��L���s���<��� ������������T�z� K��$~l��� ��,P�D� Tzh���� (�/
/@/./P/v/ d/�/��/ /�/�/�/ ??<?*?L?r?�/�? �/b?�?�?�?�?OO 8Oz?_OqO(OJO$O�O �O�O�O�O_RO7_vO��A�$SERV_MAIL  �E�vP�\XOUTP�UTkX��@@`TRV 22v V  yP (QxF_�_`TSAVE�\�zYTOP10 2}3�Y d |O 2oDoVohozo�o�o�o �o�o�o�o
.@ Rdv����� ����*�<�N�`� r���������̏ޏ��`��&� UeYP�_�]SFZN_CFGw 4 UyS�{D�Q�Uf�GRP �25p��Q ,B�   A���AD;� B���  �B4&cRB2�1�VHELLi�!6 U�V�P�_���>(�%RSR(�)� ;�t�_���������� ˯ݯ��:�%�^�I�􂿓����  �Q%��Կ濡������@���S�zG��2�@d��|�ۖHK 17� ϚϕϧϹ� �������*�%�7�I� r�m�ߑߺߵ�����~՜OMM 8��)�ڒFTOV_E�NBkT�Q�YHOW_REG_UII��^RIMIOFWD�L�9~�WAITF�Ɉ���Prj��T��TIMj�7����VAjP��>~�_UNITE��v�YLCc�TRYj��U`PMEi�:@���Q	���f�;r�� ������<����X�@Đ `	P?�  �����_'P@6�V�VMON_�ALIAS ?e��Phe1_�� ���
�%7 �[m��N� ���/�3/E/W/ i/{/&/�/�/�/�/�/ �/??/?A?�/e?w? �?�?�?X?�?�?�?O O�?=OOOaOsO�O0O �O�O�O�O�O__'_ 9_K_�Oo_�_�_�_�_ b_�_�_�_o#o�_Go Yoko}o(o�o�o�o�o �o�o1CU  y����l�� 	��-��Q�c�u��� 2�����Ϗ�󏞏� )�;�M�_�
������� ��˟v����%�П 6�[�m����<���ǯ ٯ�����!�3�E�W� i��������ÿտ�� ����/�ڿS�e�w� �ϛ�FϿ�������� ��+�=�O�a�s�ߗ� �߻���x�����'� 9���]�o����P� �����������5�G� Y�k�}�(��������� ����1C��g�y���Z�$S�MON_DEFP�ROG &����� �&*SYSTE�M*���REC�ALL ?}�	� ( �}4xc�opy fra:�\*.* vir�t:\tmpba�ck?=>192�.168.56.�1:11320 `fm��}76�mdb:home�.tpCemp\��Uk�// }�86s:orde�rfil.dat�C��|/�/�/}/ �@Y/ge/�/??�35>Pb�/z? �?�?�4E?W?j?�?�OO }\�:i�pl_fanuc�_smplgrp�_close.ls�=OOE�?�?�O3/ E/�/�2nO�O_�/�/ �O�/�OQ__"_4?�? X?j_|_�_o�?�_�_��3�_Xo�o�tp?disc 0}o�0�Rodovo�o�t�pconn 0  �o�o�o�o�*z�c =Oas���O�O D_�O����'_9_T� ]_o�����_�_Jo�_ �V�!�#o5oF��k� ՟�� ��o�?�������1�7r1}�O�a� s����)�;�ď_�� �������T�ݏo��� �%�7�ʟ[��V�!� ����F�ٯk��Ϗ� � 3�E�οi���ߞ߱� L�տg�yߋ��/��� ��e���	���>�P���u����95Ea�nimation_pick����0������%�7�dropK���o���%�7�I��� ��\��߶� Q��l���4��� X������C~��4o�/%L
xy�zrate 11 ѡ����/�//B95'},202ϡ}/ g/y/�/?��A����' �/?�?%?����[?m? ?�?#5G�?�/�? O�O�NO�+eOwO�O�_�3�$SNPX�_ASG 2<����@Q�� P 0 '�%R[1]@g1.1!_kY?��3%k_�_z_�_�_�_�_ �_�_'o
oKo.o@o�o do�o�o�o�o�o�o �oG*kN`� �������1� �;�g�J���n����� ��ˏ��ڏ����Q� 4�[���j�������� ğ����;��0�q� T�{�����˯����� ��7��[�>�P��� t���ǿ���ο�!� �+�W�:�{�^�pϱ� �ϻ�������� �A� $�K�w�Zߛ�~ߐ��� �������+�� �a� D�k��z������ ����'�
�K�.�@��� d������������� ��G*kN`� �������1 ;gJ�n�� ����/�/Q/ 4/[/�/j/�/�/�/�/ �/�/?�/;??0?q? T?{?�?�?�?�?�?O��?O7OD3TPAR�AM =@U�JQ �	�;JP��D�@�H�D�� ��3POFT�_KB_CFG � zCFU0SOPI�N_SIM  @[�F�O�O_�@Q@�RVNORDY_�DO  �E�E�%RQSTP_DS�B�N�Bi_uHQ@S�R >�I �� & IPL_�FANUC_SM�PLGRP_OPENu]yD�@Q@�TO�PN_ERR�2_OB�QPTN ��E
`�D��RRING_PR�M�_DRVCNT_�GP 2?�E�A�@x 	e_do|@Ro��ovo�o�WVD9`ROP 1@`I�@�a �I�g�o�o 2Y Vhz����� ����.�@�R�d� v������������ ��*�<�N�`�r��� ������̟ޟ��� &�8�J�q�n������� ��ȯگ����7�4� F�X�j�|�������Ŀ ֿ������0�B�T� f�xϊϜ��������� ����,�>�P�b߉� �ߘߪ߼�������� �(�O�L�^�p��� �����������$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@gd�v�����bPRG_COUNT�Fs�
b�ENBo��M#�D/_UP�D 1A�[T  
�{Bf/x/�/�/ �/�/�/�/�/??C? >?P?b?�?�?�?�?�? �?�?�?OO(O:OcO ^OpO�O�O�O�O�O�O �O __;_6_H_Z_�_ ~_�_�_�_�_�_�_o o o2o[oVohozo�o �o�o�o�o�o�o
3 .@R{v��� ������*�S� N�`�r���������� ޏ���+�&�8�J�s� n���������ȟڟ������_INFO� 1BT%: \�	 3�w�b������?*&�?����>Y�L=��n-�����h>F��d9��]/�𡯈��'� D�&t����D�)�´ ��E�³��*��<��YSDEBU)G�U �*�d=)e�SP_PASS��B?w�LOG �CQ�^!  r*�#�0�  �9!�*�UD1:\x��7���_MPC���T%%�7�T!�U� �T!�SAV D���!�̱�$���SV��TEM_TIME 1E���_  0  P(��#����ù��MEMBK  T%9!̰̿9�K�[��X|: � @[�(��}ߢ߲�v�d������r� �@���,�>�P��h��z�������� � ������0�B�T�f�x����e�������� ��*<N`r ���������SK���$߰Tfxl��*�|��2�߷#� ��� )����������</�N/`/7.e�� ��/�'�7/�/�/�/���2�?;?M?_?q?�?*�U�?�?���?'�n�?�?OO1O COUOgOyO�O�O�O�O��O�O�O	__-_=�T�1SVGUNSP]D�� 'w��HP�2MODE_LI�M F��{�DT2�QPqQG��CUAB�UI_DCS 	J7w�F�'�_�$��$G�6_�\o�WG�*7���9a 
?`�$9o'�Sh��Scɼ��UEDIT �K�_�XSCRN �L���R�G �M�[�U�:�eS�K_OPTIONpl��{��b_DI��?ENB  �%w���aBC2_GRP 2N�Y���o���0C��s<\BCCeF�`P]{�� ����v`����� !�G�2�k�V���z��� ��׏ԏ���1�� U�@�y�d�������ӟ �������?�Q�g ^�p�������0�ٯį ����3�a�N��#� V�|�j�����Ŀ��� ֿ�����B�0�f�T� ��xϮϜϾ������ ��,��P�>�`�b�t� �ߐ؆`������ �� ��6�$�F�l�Z��� ����������� �� 0�2�D�z�h������� ��������
@. dR�v���� ���0N`r �������/ /�8/&/\/J/�/n/ �/�/�/�/�/�/�/"? ?F?4?V?|?j?�?�? �?�?�?�?�?�?OBO 0OfO~O�O�O�O�O PO�O�O_,__P_b_ t_B_�_�_�_�_�_�_ �_�_o:o(o^oLo�o po�o�o�o�o�o �o $H6XZl� ��|O��� �2� �V�D�f���z��� ԏ������
�@�.� P�R�d���������� П����<�*�`�N� ��r���������̯� �&��>�P�n����� �����ƿ�ڿ�"� 4��X�F�|�jϠώ� �ϲ���������B� 0�f�T�vߜߊ��߮� ���������,�b� P��<���������� p���&�L�:�p��� ��b��������� �� $ZH~l� ������  D2hVxz�� �����/./@/R/ �v/d/�/�/�/�/�&�� �$TBCSG_GRP 2Q�%��  ���! 
 ?�  ?+??O?9?s? ]?o?�?�?�?�;�"�#�S <d�H�A?�!	 HA�����5>���>�=q?�\�5?AT��A 2HO�THJ�ff?aG'�?L G>BpTOVN	�t@#E� @wA� 6Jy��O�M@��RjI�>�33*A�5�ABCO�O�H�BPOQY9�,_.^��HBY�ArBU�PB�t_.^�H �6�H�U�_�_�_ o=o@ooho�o�kjh��a	V3.002�	crx�c�`*��`�d�"8T�O ?�dS� Hqji p��m  �3C��oY`s�!J2�#T� =`lxCFG [V�%
1 0V�z��r,r��x�����  �E�0�i�T���x��� ��Տ��ҏ���/�� S�>�w�b�������џ ��������=�(�:� s�^�������ͯ2+  د�����/��?�e� P���t�����ѿ��� �¿+��O�:�_υ� �!�/�϶/�ϼ���� ��(��L�:�p�^߀� �ߔ��߸������ � "�$�6�l�Z��~�� �����������2� � V�h�(/����<����� ������
@.P v��X���� �*<Nr` �������/ /8/&/\/J/l/�/�/ �/�/�/�/�/�/?? "?X?F?|?j?�?�?�? �?�?�?��O$O6O�? fOTOvOxO�O�O�O�O �O__,_>_�Ob_P_ �_t_�_�_�_�_�_�_ oo:o(o^oLo�opo �o�o�o�o�o �o$ H6X~l�� �������D� 2�h�V�����HO��ȏ ����
���.��R�@� b�d�v�����П���� ���*��N�`�r��� >�����̯��ܯ�� &��J�8�n�\�~��� ��ȿ���ڿ���4� "�D�j�Xώ�|ϲϠ� ����������0ߪ�H� Z�l�ߜߊ߬����� ������>�P�b�t� 2���������� �����L�:�p�^��� ������������  6$ZHjl~� ����� 0 VDzh���� ~����ߺ@/./d/ R/�/v/�/�/�/�/�/ ?�/�/<?*?`?N?�? �?�?�?t?�?�?�?�? O8O&O\OJO�OnO�O �O�O�O�O�O�O"__ F_4_V_X_j_�_�_�_ �_�_�_o�_oBo0o fo�/�o�oLozo�o �o�o,P>t ���h���� �(�:�L�^����p� ����ʏ��ڏ܏�$� �H�6�l�Z���~��� Ɵ���؟���2� � B�D�V���z�����ԯ ¯��
��o"�4�F�� v�d������������� ��*�<�N��r�`�p�τϺϤ�  ����� ��������$TBJOP_G�RP 2W����  ?_���C��	���Y�����X  ���Y� �,? � �x��ï @��?}�	� �A��͔�C�  D�ǌь��>0�>\?��е�aG�:��o��;ߴAT3�ͰՌ�A��Ӭ����ߦ�>�я\�)?��D�8Q��Ѵ�L��>̼����;iG�Ҍ�z�Ap�Љ� ��A�ff��0��m�������:VM��ҹ�R����)���@��RD�Cр��щ�pi�e�H�Q��ff���:�6/D�33��B   ������D�V�h�Q�Q�x���:ǲS���}�,B�x6?Q@��Hd���r����d�=m�<�#�
���0�;/˚�d���B� ����ٰ��"� �:kF �� ������/4/`/,/Z/�/��C������!��	V3.{005�crx�#� *� i�������*� C�  E�$` E�h E�ܨ F� F�3� FV4 F�x� F�� F�� F�X F��0�� F�F� F�� Gs� G G�� Gk G&��#�� Y? E@� E�� E��� E� F�� F2 FN�� Fj� F��� F�� F�� F�H F�|� Fʰ 9�IIR�1t,H�5 *��T�?�2���3?����`-�ED_TC�H Z��(�#e����h���d$�(ЄO�O��� �TE�STPARS  ���SC�HR�@A�BLE 1[�� @��fւҞG�:�G�H�H����*�G	�H
�H�HU����H�H�HN�FRDI�O(�_@_%_7_I_[U�TO�_��[�_�_oo/n�BS�_&� �Z�o& 8J\n���� �����"�4�F� ��`�o'� W��po�o �o�oR_d_v_�_�_�X��Bm�NUM  V��(�p���� �@�P�B_CFGG \V����@��IMEBF_TT��A��PE��VER�SfѮ���R 1=]�K 8zO������ ����   ���)�;�M�_�q� ��������˯ݯ�� �%�7���[�m����� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/�x� S�e߮߉ߛ߱߿��� �����:Bۑ_P�Ŗ�@ϕ<@LIF �^V��0ʑ�Њ���"��( 0
u��@��@� d���W�MI_CHANꤗ ϕ ��DBG�LVL��PF��E�THERAD ?)�E����0��x7�I���ROUT!HJ!}�����?SNMASK�ϓ>$�255.���#��������#<@OOL?OFS_DI�@R0�����ORQCTRL _�K;c�?yTh������ 	-?Qcu� ����g��/�9CPE_DETA�I��>
PGL_C�ONFIG e�V�f���/ce�ll/$CID$/grp1/�/�/�/�/�/6c�d�?? %?7?I?[?�/?�?�? �?�?�?h?�?O!O3O EOWO�?�?�O�O�O�O �O�OvO__/_A_S_ e_�O�_�_�_�_�_�_ r_�_o+o=oOoaoso��}o�o�o�o�o�o �/+
}�o` r����o�� ��&�8��\�n��� ������ȏW����� "�4�F�Տj�|����� ��ğS������0� B�T��x��������� үa�����,�>�P� ߯t���������ο� o���(�:�L�^�� �ϔϦϸ�����k� ߀�$�6�H�Z�l�g ��User V�iew |)}}1�234567890�߯�����������X2�}������2�� ��a�s������,��3D�	��-�?� Q�c����2�4��� ������v�82�5��q�����*�2�6`%7I@[m��2�7 ���/!/3/�T/2�8��/�/�/�/�/��/F/?2 l�Camera �ڄ/M?_?q?�?�?�?�bE@?�?�?�>��O�!O3OEOWOiO_	   '6C�<?�O�O�O�O_ _�?7_I_[_�O_�_ �_�_�_�_ ?�'6�� p_%o7oIo[omoo&_ �o�o�oo�o�o! 3E�_�W���o�� �����o�!�3� ~W�i�{�������X �W�KJ����#�5�G� Y� �}������şן �����Ə(5�� i�{�������ïj�� ���V�/�A�S�e�w� ��0��W� �տ��� ��/�֯S�e�w�¿ �ϭϿ������Ϝ��W {)��A�S�e�w߉ߛ� BϿ�����.���+� =�O�a���9�ߢ� ������������2� D���U�z�����������c*	)50Z�! 3EWi���� X����/�� ��.00;����� ���//*/uN/ `/r/�/�/�/O)5�K ?/�/??*?<?N?� r?�?�?�/�?�?�?�? OO�/��k�?`OrO �O�O�O�Oa?�O�O_ MO&_8_J_\_n_�_'O 9Et{_�_�_�_oo &o�OJo\ono�_�o�o �o�o�o�o�_9E���o 8J\n��9o� ��%��"�4�F� X��o9EL������ȏ ڏ����"�4�F����j�|�������ğk�  o����)� ;�M�_�q����������   ə?fffB�Pߡk����� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢϴ��� ������� �2�D�V� h�zߌߞ߰������ߠ��
��.���
k�(�  ��( 	 ;�q�_���� �����������7�%��[�I����� ��������[� 0BTfm����� ������ 2 yVhz���� ���?/./@/� d/v/�/�/�/�/// �/??_/<?N?`?r? �?�?�/�?�?�?%?O O&O8OJO\O�?�O�O �O�?�O�O�O�O_"_ iO{OX_j_|_�O�_�_ �_�_�_�_A_o0oBo �_foxo�o�o�o�oo �o�oOo,>Pb t��o�o���' ��(�:�L�^���� �����ʏ܏� �� $�k�H�Z�l������� ��Ɵ؟�1�C� �2� D���h�z�������¯ 	����
�Q�.�@�R� d�v���ϯ����п� ����*�<�Nϕ�u�@ p�}Ϗϡ�p��w�[��� fr�h:\tpgl\�robots\c�rx��10ia.xml]���� �2߀D�V�h�zߌߞ߰�  �����������  �2�D�V�h�z��� �߯�������
��.� @�R�d�v�������� ������*<N `r������� �&8J\n �������� /"/4/F/X/j/|/�/ ��/�/�/�/�/?? 0?B?T?f?x?�?�/�? �?�?�?�?OO,O>O@PObOtO�O�N���� w���<<; �� ?��K�O �O�O�O#_	_+_Y_?_ q_�_u_�_�_�_�_�_ o�_%oCo)o;o]o�o�����(�$TP�GL_OUTPU�T h������` �jfffB4  �a���o 
.@Rdv� ���������*�<�N�`�r������ ��`cell/�floor/wa�ll rite �3456789012��ʏ܏� �� ���`�/�A�S�e�w� �!�����џ������}�6�H�Z�l�~� �(���Ưد���� ���D�V�h�z���$� ��¿Կ���
Ϣ��� @�R�d�vψϚ�2Ϩ� �������߰�&�N� `�r߄ߖ�.�@����� ����&��4�\�n� ����<�������� �"�����X�j�|��� ����J������� 0��>fx����F�b $$ zb����:, ^P�t���� ��//6/(/Z/L/ ~/p/�/�/�/�/�/�/?}�A(?:?L?^?p?��?�=@�O�?�?�J? ( 	 ?�? �?"OOFO4OjOXOzO |O�O�O�O�O�O_�O 0__@_f_T_�_x_�_ �_�_�_�_�_�_,oo�Po���  <<?�o�o�`to�o �o�o�o��qo7I �oUYk��% ����3�E��i� {��c���K������ ӏ�/����e�w�� ���������A�S�� +�ş3�a�;�M����� �ͯ߯y�˯��� K�]���e���-��ɿ ۿ�����o���G�Y� �}Ϗ�iϗ���#ϭ� ��ߧ�1�C��/�y� ���ϯ���[������� ��-�?��C�u��a� ��������Q���)� ���_�q�K������ ��������%��1 [������=�� ��!EW��C�gy��gb)�WGL1.XM�L�?
-�$TPOFF_LIM l`|�0ha�&�N_SV    ��42*P_MON7 ide4$�0��02)STRT?CHK jde2&�%?"VTCOM�PATG(�!6&VW�VAR kg-\�(K$ �/ ?�0z"!_DE�FPROG %��)%IPL_�FANUC_SM�PLGRP_CL�OSE�/?0ISP�LAY' �.<2IN�ST_MSK  �< x:INU�SER�/~4LCK��<�;QUICKM�EN�?~4SCRE�@de�"tpsc~4�1.@3I2"�D@_HIST�*2)R�ACE_CFG �lg)�$0	�4
?��HHNL� 2mK:D`�A�+  !2�O�O__/_A_S_�e_wZ�EITEM �2n�K �%$�12345678�90�_�U  =<��_�_�_c  !
ok0�_Wo3�_ xo�_�o�oo�o6oHo lo,�o<b�o�o �o�o �D�� (��L����N�� ��ʏ܏@��d�v��� �Z���~���􏜟� *��N��r�2�D��� Z�̟����¯&�ү ��
�n��������0� گ������"��F�X� j��Ϡ�`�r�ֿ~� �����0���T��&� ��<߮��ω��Ϥ�� ����`�P�b�tߎߘ� ��h������(� :�L���p��B�T��� `����� �����6��� l�����k��� ���� �D� z:�Jp��� 
.�R�$/6/ �Z/���f/~// �/�/N/�/r/�/M?�/ h?�/�?�??�?&?8?�O�DS�Bo�OJψ  �RJ 8�A]OT9
 jO�O�wO�O5JUD1:�\�L��AR_G�RP 1p�[?� 	 @�@_ [_>_,_b_P_�_t^��P�_�Z�Q�O�_�_<	o�U?�  $o6k  oVoDozoho�o�o�o �o�o�o�o
@.0dRt�	�5���CSCB 2q"K o��0��B�T�f�x�����LU�TORIAL �r"K�O�GV_C�ONFIG s�"M�AZO�OF���OUTPUT t"I7���R����� ��̟ޟ���&�8� J�\�n�4��������� ̯ޯ���&�8�J� \�n��������ȿڿ ����"�4�F�X�j� {��Ϡϲ��������� ��0�B�T�f�x߉� �߮����������� ,�>�P�b�t�ߘ�� ����������(�:� L�^�p���������� ���� $6HZ l~������� � 2DVhz �������
/ /./@/R/d/v/��/ �/�/�/�/�/??*? <?N?`?r?�? �2��� �?�?�?�?
OO.O@O ROdOvO�O�O�/�O�O �O�O__*_<_N_`_ r_�_�_�O�_�_�_�_ oo&o8oJo\ono�o �o�o�_�o�o�o�o "4FXj|�� �o������0� B�T�f�x�������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@߀R�d�v߈ߚ߬ߏ8��������Ѷ� �?,�>�P�b�t�� ������������� (�:�L�^�p������� �������� #�6 HZl~���� ���2DV hz������ �
/./@/R/d/v/ �/�/�/�/�/�/�/? ?)/<?N?`?r?�?�? �?�?�?�?�?OO%? 8OJO\OnO�O�O�O�O �O�O�O�O_!O4_F_ X_j_|_�_�_�_�_�_ �_�_oo/_BoTofo xo�o�o�o�o�o�o�o +o>Pbt� ���������%��$TX_SCREEN 1u����М}�ipnl/Y�g?en.htm%�x����������/pP�anel setupČ}�ď��)�;�M�_��鏖� ����̟ޟ�g���� 8�J�\�n�����	�� ȯگ����"���ǯ ��j�|�������Ŀ;� �_���0�B�T�f� ݿￜϮ��������� mϛϑ�>�P�b�t߆� ��߼�3��������(�:��(�UALR�M_MSG ?E��R� S�(z�� ������������� ;�A�r�e�������n�SEV  |����l�ECFG �wE�O�  }(u@�  A�   B�(t
 ��/sE�Oas� ������~��GRP 2xw 0(v	 9�[n�I_BBL_NOTE y
�T��l�/rJ�/q nDE�FPROx�%|� (%���2p�� � //D///h/S/y/��/�/�/�/�/dFK�EYDATA 1yzE�Ep (vHK?]?4?�?�?�j:,(�?�?(t�0�ǲ���?�?�1��� ��Z���?��>:OLO�5�һ�� e�b�vRO>�<��C��~O�O�8@��� Ə������O,O�O�O �O#_
_G_Y_@_}_d_��_�_�_�_�_�_f>���  frh/g�ui/white�home.png�oIo[omoo�o hpoint4o�o�o�o��o�hFRH/F�CGTP/wzcancel�oN` r���c����p���%nex�o�S�e�w������ntouchupC�׏������*�/infoƏZ�l�~������ Ɵ؟���� ���D� V�h�z�������?�ԯ ���
��.���R�d� v�������;�п��� ��*�<�˿`�rτ� �ϨϺ�I������� &�8�oG�n߀ߒߤ� �����������"�4� F���j�|������ S�������0�B�T� ��x�����������a� ��,>P��b ������o (:L^��� ����k�/$/ 6/H/Z/l/��/�/�/ �/�/�/y/? ?2?D? V?h?�/z?�?�?�?�? �?�?�?O.O@OROdO�vOM��K�`����O�O�M�O�O_�F,�_5_�_Y_ @_}_�_v_�_�_�_�_ �_o�_1oCo*ogoNo �o�o�o�o�o�o�o	 ?&cuTߙ �����O�)� ;�M�_�q�������� ˏݏ����%�7�I� [�m�������ǟٟ ������3�E�W�i� {������ïկ��� ���/�A�S�e�w��� ��*���ѿ����� ��=�O�a�sυϗ�&� ����������'߶� K�]�o߁ߓߥ�4��� �������#��G�Y� k�}�������� ����1�8�U�g�y� ��������P�����	 -?��cu�� ��L��) ;M�q���� �Z�//%/7/I/ �m//�/�/�/�/�/ h/�/?!?3?E?W?�/ {?�?�?�?�?�?d?�? OO/OAOSOeO�?�O �O�O�O�O�OrO__ +_=_O_a_�O�_�_�_��_�_�_�_���[}������o@.o@mobotoNf,` �oX�o�o�o�o�o# 
GY@}d�� ������1�� U�<�y���r�����ӏ ���	��-�?�Q�c� r_��������ϟ�� ���)�;�M�_�q� � ������˯ݯ�~�� %�7�I�[�m����� ��ǿٿ�����!�3� E�W�i�{�
ϟϱ��� ������ߚ�/�A�S� e�w߉�߭߿����� ����+�=�O�a�s� ���&��������� ���9�K�]�o����� "�����������# ��GYk}���� ����1� Ugy���>� ��	//-/�Q/c/ u/�/�/�/�/L/�/�/ ??)?;?�/_?q?�? �?�?�?H?�?�?OO %O7OIO�?mOO�O�O �O�OVO�O�O_!_3_ E_�Oi_{_�_�_�_�_ �_d_�_oo/oAoSo �_wo�o�o�o�o�o`o �o+=Oa8 �c{�8 ������}����v,Џ�ȏ9� �]� o�V���z���ɏ��� ԏ�#�
�G�.�k�}� d�����ş������ ��C�U�4y����� ����ӯ�o��	��-� ?�Q�c�򯇿������ Ͽ�p���)�;�M� _�ϕϧϹ����� ��~��%�7�I�[�m� �ϑߣߵ�������z� �!�3�E�W�i�{�
� ������������� /�A�S�e�w������ ����������+= Oas���� ���'9K] o��j����� �/5/G/Y/k/}/ �/�/0/�/�/�/�/? ?�/C?U?g?y?�?�? ,?�?�?�?�?	OO-O �?QOcOuO�O�O�O:O �O�O�O__)_�OM_ __q_�_�_�_�_H_�_ �_oo%o7o�_[omo o�o�o�oDo�o�o�o !3E�oi{� ���R���� /�A��e�w�������h��я�Ӌ�������� ���B�T�.�,@���8� ����͟ߟƟ��'� 9� �]�D�����z��� ��ۯ�ԯ���5�� Y�k�R���v���ſ� �����1�C�R�g� yϋϝϯ�����b��� 	��-�?�Q���u߇� �߽߫���^����� )�;�M�_��߃��� ������l���%�7� I�[������������ ����z�!3EW i�������� v/ASew ������� /+/=/O/a/s//�/ �/�/�/�/�/?ڿ'? 9?K?]?o?�?�/�?�? �?�?�?�?O�?5OGO YOkO}O�OO�O�O�O �O�O_�O1_C_U_g_ y_�_�_,_�_�_�_�_ 	oo�_?oQocouo�o �o(o�o�o�o�o )�oM_q��� 6�����%�� I�[�m��������D� ُ����!�3�W� i�{�������@�՟�@����/�A�0C���0����l�~���h���į��, ������� �=�O�6� s�Z�������Ϳ��� ��'��K�]�Dρ� hϥό����������� #�5�?Y�k�}ߏߡ� ����������1� C���g�y������ P�����	��-�?��� c�u�����������^� ��);M��q �����Z� %7I[�� ����h�/!/ 3/E/W/�{/�/�/�/ �/�/�/v/??/?A? S?e?�/�?�?�?�?�? �?r?OO+O=OOOaO sOJߗO�O�O�O�O�O �?_'_9_K_]_o_�_ _�_�_�_�_�_�_�_ #o5oGoYoko}oo�o �o�o�o�o�o�o1 CUgy��� ���	��-�?�Q� c�u�����(���Ϗ� �����;�M�_�q� ����$���˟ݟ�� �%���I�[�m���� ��2�ǯٯ����!� ��E�W�i�{�������ڈ@����@���ܿ� �ؿ"�4��, �e�߉�p� �ϿϦ������� � =�$�a�s�Zߗ�~߻� �ߴ��������9�K� 2�o�V���O���� �����#�2�G�Y�k� }�������B������� 1��Ugy� ��>���	 -?�cu��� �L��//)/;/ �_/q/�/�/�/�/�/ Z/�/??%?7?I?�/ m??�?�?�?�?V?�? �?O!O3OEOWO�?{O �O�O�O�O�OdO�O_ _/_A_S_�Ow_�_�_ �_�_�_�_��oo+o =oOoaoh_�o�o�o�o �o�o�o�o'9K ]o�o����� �|�#�5�G�Y�k� }������ŏ׏��� ���1�C�U�g�y�� ������ӟ���	��� -�?�Q�c�u������ ��ϯ�����)�;� M�_�q�����$���˿ ݿ��Ϣ�7�I�[� m�ϑ� ϵ�����������!��P#��>�P���L�^� p�Hߒߤ�~�,���� �������/��S�:� w��p��������� ���+�=�$�a�H��� l����������� �_9K]o���� �����#� GYk}��0� ���//�C/U/ g/y/�/�/�/>/�/�/ �/	??-?�/Q?c?u? �?�?�?:?�?�?�?O O)O;O�?_OqO�O�O �O�OHO�O�O__%_ 7_�O[_m__�_�_�_ �_V_�_�_o!o3oEo �_io{o�o�o�o�oRo �o�o/AS* w������o� ��+�=�O�a���� ������͏ߏn��� '�9�K�]�쏁����� ��ɟ۟�|��#�5� G�Y�k���������ů ׯ�x���1�C�U� g�y��������ӿ� �����-�?�Q�c�u� ϙϫϽ�������� ��)�;�M�_�q߃�� �߹���������%�7�I�[�m���hp����hp��������������, E���i�P����� ������������ AS:w^��� ����+O 6s�d���� �/�'/9/K/]/o/ �/�/"/�/�/�/�/�/ ?�/5?G?Y?k?}?�? ?�?�?�?�?�?OO �?COUOgOyO�O�O,O �O�O�O�O	__�O?_ Q_c_u_�_�_�_:_�_ �_�_oo)o�_Mo_o qo�o�o�o6o�o�o�o %7�o[m ���D���� !�3��W�i�{����� ��Ï������/� A�H�e�w��������� џ`�����+�=�O� ޟs���������ͯ\� ���'�9�K�]�� ��������ɿۿj��� �#�5�G�Y��}Ϗ� �ϳ�������x��� 1�C�U�g��ϋߝ߯� ������t�	��-�?� Q�c�u������� ������)�;�M�_� q� ���������������$UI_IN�USER  ����"��  _�MENHIST �1{" � ( / ���)/SOFTP�ART/GENL�INK?curr�ent=menu�page,1133,1A����s� |�962��6HZl�36%������5�B/T/f/�//�6w/�/�/�/y/��/�/�ON_PICK�Q?c?u???��I9?�?�?�?�?,�?�?81� 2OROdOvO�M����v�A �O�O�O�O�O�O_A '_9_K_]_o_�_�_"_ �_�_�_�_�_o�_5o GoYoko}o�oo�o�o �o�o�o�oCU gy��,��� �	���?�Q�c�u� �������OϏ��� �)�,�ʏ_�q����� ����H�ݟ���%� 7�Ɵ[�m�������� D�V�����!�3�E� ԯi�{�������ÿR� �����/�A�п� wωϛϭϿ��ϼ��� ��+�=�O�a�dυ� �ߩ߻�����n��� '�9�K�]��߁��� ��������|��#�5� G�Y�k���������� ����x�1CU gy����� ���-?Qcu �������/ �)/;/M/_/q/�// �/�/�/�/�/??�/ 7?I?[?m??�? ?�? �?�?�?�?O�?3OEO WOiO{O�O�O.O�O�O��O�O__�$U�I_PANEDA�TA 1}����KQ  �	�}  fr�h/cgtp/f�lexdev.s�tm?_widt�h=0&_hei?ght=10{PlP�ice=TP&_�lines=15�&_column�s=4{Pfont�=24&_page=wholelP�'_)  rim�_�_  \P
oo.o @oRodo�_vo�o�o�o �o�o�o�o�o<N 5rY������ �  �   �� o	��-�?�Q�c�� ���_����Ϗ��� l�)�;�"�_�F����� |�����ݟ�֟��� 7�I�0�m��y��MS ������ѯ����Z� +���O�a�s������� �Ϳ߿ƿ��'�9�  �]�Dρ�hϥϷϞ� ������߄���G�Y� k�}ߏߡ�����8��� ����1�C�U��y� `������������ �-��Q�8�u���n� ���0�����) ;��_q�ߕ�� ���V�7I 0mT����� ���!//E/���� ��/�/�/�/�/�/:/ ?~/?A?S?e?w?�? �/�?�?�?�?�?OO  O=O$OaOHO�O�O~O �O�O�O�Od/v/'_9_ K_]_o_�_�O�_?�_ �_�_�_o#o5o�_Yo @o}odo�o�o�o�o�o �o�o1UgN ��O_����	� �n?�Q��_u����� ����Ϗ6��ڏ�)� �M�4�q���j����� ˟ݟğ��%���}�6�o���������ɯ)]��a�ݯ�,� >�P�b�t�ۯ����� �����ٿ���:�L� 3�p�WϔϦύ���Z���s�{�$UI_P�OSTYPE  ��u� �	 ��-���QU�ICKMEN  ���0���RE�STORE 1~��u  '���a��ߴ���a�m������1� C���g�y����R� ������	����(�:� L������������r� ��);M��q ����d���� \%7I[m� ����|�/!/ 3/E/��d/v/��/ �/�/�/�/?�//?A? S?e?w??�?�?�?�? �?�/�?OO�?OOaO sO�O�O:O�O�O�O�O __�O9_K_]_o_�_�;�SCREK�?�P�u1sc���u2�T3�T4��T5�T6�T7�T8ܼQ�STAT�� �_Ӵu��USERx�P�_�RTPSC�SSks�SWd4Wd5Wd�6Wd7Wd8Wa��N�DO_CFG ��F�E���OP_CRM5  A���f��PD�Q9i�None>��0`_INFO 2Հ�up]�0% �_Z�
K.o� d���������5�G�*�k�4��aO�FFSET ��qx�"S��*_�� Ώ�����(�U�L� ^���b��������ܟ ���$�6���`߂�p���
��ʯV�a�aWORK ��m�������z�/`U�FRAME�o�R�TOL_ABRT8i��c��ENB��{�?GRP 1���\�Cz  A�� ޱ"Q޿���&�8�!B�T�y�J�U���a~��MSK  ���q��Nf�%�i��%R��ϛ�_EVNĉ����f֑b3�
 h�aU�EV��!td:�\event_u�ser\��M�C7�Rߧ��`F׭F�SP�K�P�spotw�eld��!C6 �߈ߚ߾P��!��a� �T��ו��C�1�� ��g�y��������� ��^�	���-�?�u��� ����������6%Z �;��q�@�� ��
"�W�33�:i��8�� r����/ �'/9//]/o/J/�/ �/�/�/�/�/�/?�/�5?G?"?X?}?�?�$�VALD_CPC� 2��� 8k?�?�a O��Q�<�*�O7OIO��"S&BdpJm@j��IlD[ �OV�?�O�?�?_O /_A_S_bOtO�O�O�_ �O�_�O�O(_oo=o Oo^_p_�_�_�_�_�o �o�_ o$o9K�o lo~o�o�o]�o��o �o� �G�Y�hz ����׏b��
� �.�C�U�d�v����� ����Џ����*� +�Q�c�r��������� ̟����)�8�M� _�n���������˿گ ����%�4�I�[�m� |�����Fϴ�ֿ���� ��3�B�W�i�xϊ� �Ϯ����������� /�>�S�e�w�ߘߪ� �߾�������L�=� ,�a�s�������� �����$�9H�] o����������� � �D6k} �������� .C/Rg/y/�� ����/�	?/*/ ?N/O?u?�?�/�/�/ �/�?�/O?&?8?MO \?qO�O�?�?�?�?�? �O�?_"O4OI_XOm_ _�_�O�O�Oj_�_�O o_0_B_Wof_{o�o �_�_�_�_�_�oo ,o>oSbow���o �o�o�o��(: pa�P�������� �� ��'�6�H�]� l�����*���Ə؏� ���#�2�D���h�Z� ������ԟ����
� ���@�R�g�v����� ����Я���	��-� <�N�5�r�sϙϫϺ� ̿޿����)�8�J� \�q߀ϕߧ߶����� �����"�7�F�X�m� |ߑ��������ߎ� ���3�B�T�f�{��� ������������� ,�AP�b�w���� �������(= L^��t��� �� $&/K/Z l�/��/�/N/�� �/�/2/G?V/h/"? �/~?�?�?�/�/�/?�?.;�$VARS�_CONFIG ��i0PA�  FP53��4LCMR_GR�P 2�PK��8�1	a0\@  %�1: SC13?0EF2 *�O�@�54�.5i0��8�0��5`0`1?�  �A@�@p
@�.N &OX_.8<_�N_{_�Av_�_UA)��@�Q�52�_�_�52 B��� �Q51�U�_ og_Doo hoSo�owo�o�o�o�o =o�oRov��<DIA_WOR�K �PE�p<z0�6,		j1PE|��wG�P ��p�Y9�qRTSYNC�SET  PI��PA�WINURLg ?�b0���X�j�|��������vSIONTMOU��53<� �ʅ_�CFG �S����S۵P~Z@ FR:\̃�\DATA\�� ��� UD1��LOG�  �1�EX=�51' B@ ����P�=?��P���ş.7� � n6  ���.6|��<����A  =�����54�Q�TRAI�Nf���&� 
�7!p��v�]4#��:|B�PK (?qg� ��7y����ӯ���-� �Q�?�Y�c�u�����\��Ĉ_GE�PK7�``0�
z0x2,�c�RE���PE�.8HLEX�PLa0�1-e��VMPH?ASE  PE�3��P=CRTD_F�ILTER 2�.PK ��E�_�� ������,�>�P�b� t�.7�Ϣߴ����������� �2�D�7ISH�IFTMENU {1�PK
 <k<1%����݂����� ����������K�"� 4�Z���j�|������������	LIVE�/SNA`C%v�sflive��+̃ �U`@4menuJO������r`��5�Y�M�O�Q��@@@Z�D��.�51<Y���P�$WAITDINEND׈`1�>HOK  �Ic�Պ~S�eTIM.ׅ���GO� q+�����cRELE|�'�Hxҏ�J_ACT' �(�qc_� ���y�%�?9F�"R�DIS`@�.�$�XVR��Q���$ZABC{B1�N+ ,Y�Bu2?�2M!� VSPT ��Q͚E�
�
��?�
�?O�7�DCSCHG ���{�@�04GBph0I-P$�+A�O��O�O�:MPCF_OG 1��IA�0��X�7_�OMPn3��I��p���?o_=���  3~�� �w�?�?��vԿ�P�R����~�lD&�t����D�)��?^U���=��Q�w@t_�_ �_�_�_�_�_#`d2u�Vo<o^_�o�ei´� ²E�³#��o�h�h�`�o �o&P{�_�_o� b0&o8od4�@�����O�t_CYLINuD����K �}f ,(  *��&���O�6�s�Z� �o����͎���_� ����J���n����� Տ��Q�7��ӟ��� e�F�X��|����G�! �_�����3�o�ܯǯ �婓�0�姖�J�A��tSPHE_RE 2��}̪� ����������(�;� �(Ϥ�L��ѿ��i� �ύ�������5�G�$� ��H�/�A�~��Ϣߴ�l��h0ZZ�& ��