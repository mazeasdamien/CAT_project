��   C��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN��/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER��q�C_GRP6�P L$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� )DEX� �5O n�8BUF�7TDP�HG�_@FO�SxAV��7R?EC_TRQX��MFLG�J5�� � � N IU�
@!(UF*����4OSV3EN_CG"��0_�!�AU�SCH2�SMP]L4PEXE���2�!_�SUR}A�`jAaW�@A@bVNE|Y]QnAVA?�UY�T7D�VWWnAF�[V�A�\�WTO�0oH
e7D�f�3
e�U
e�W QT�P�0IR	 DMM��A@  @ �$la�EREG_�OFS�aME�hA1SS1�A !la�RE-   �# �0�b{F�c{ĥd� M�d�b�c$�STD�hq�gFA � �h!q�g�"�f�"�c�/ la7   �$p`TIN�@��0SUL� �R}_@  $}�@ SW@�rO:}rR%	 dp~t� �@JU� �sq�FS4D6
 �' $�0PGF`QC?!$FIL� �@�E�PmA�s&�sDIG4o@SCA��$�INTTH�RS_BI�AZ�S�MAL%�COL���qATE_TI�PROG�4U�s��!CMDA  ��FSOUTENV�6P $H_RZ_AXl�CU3VR2QLB܊�0���H������PN�T_MV_AVRʤCS!pLkp�c$�L���fO�\��STt�d�F�#STO �v�FX�LECT�EDCp�Y{���FYd��t�Z{�ړFZBc�R�e��	�/ G#P~�X $��c_IV����$!�0B"0�?0F�CC�BDDN=�CCI�c�DUMMY23<G ^�DEBU�A\!4PN�"TO�q9RP" � Q09T6�� �;!��NfBUTTSP� (~@�q֥E40N ڡFS3ՁKQ1�r�9T�I�NEW_�UI��VKP�?Up`��CCOORD8\TCH���01�P��$mP��7 �l �!�3$�WEIGH���2 Us_�aF��T���WA{Q����NTER�Q��- ޵� �c��r�AS0�$JZA7STA�� �a��P� �,�26�36āW�!Ƨ ��ä"C*��Xw�Yw�Zw�_�CM��?��D��i�RSLy�u���~� �Ǝ��ƚļ��!�@ҡ�T   E�0c"0VROUN�DCMVPERIO���$F1PUU3F2D�'TM1� ��S�_DcGAMqMc1b�TRX�U�Kt�K�K��CLt�`�&O00ADJ�GA�UPDC0R"�2��E� QRED���GFR_� _@W۲���u�DL_R���@�=�M_�5d�0 n�#��}�"��}�� k�����������}�VLj�"����A� 7���`��L�P5A8@
� 
D�A�����"�8��y"��VIBƦ�OV��DEH�֌� �`,����*�� �: RTZ�MN1SUfwMN2YUFRA q	��ShZA
`-G����OR�P�ҡAL�ҤCJ��
L��"�S8B�I$L .$M"�P30+�Q �)k�}�S"PHCmD�GVz�GV��;GVړJDO°]���S�$R�E����b�]�A�AP�)�DA��3$VF�����1LVu��@IL�A���� #��  "�@fR!��$�DC+�����B #П�5'OBOA@�vYԣW2
�G'	�$�ԍ$!#¿�E�K�`�+�eCNPRGOV6��%'PN�t_TW,��"G�3E�MNV�6c0�4WT�cW�TRL/_SKIj�J�qcMN��GW6�
eR</ENABF�|qV�!� A$SB}��xS��� {P�tyR*�tX�yRQT$���2_Q��?p����ALARMSsER�QETOTD?FRZCHK1��
��62�9NC�4N@ �5L`N@�:vJ��vE�2�2�;2�=NA9E�FFIX2��BF�䦠@qI�dD���DON�t̆95PSFW�0_D;F1"%BF2/_vJ���|��4|�Pl��33=��5|�kH|�yJ�Z(��U�23�;3�=|�9E�SDIAu �6�R�Kq�B�VvEfvC&�3GA�@�@���R <iV1<d��sP�VQ�U�Uf�S$��� ���FU�ED�S_HA�U�e�d�4GEF�k@�2�`�;�a���5!%�UzKq�#H�X���s����Y��a�_FSIW�� � *�X��RK��`H7p_�CHCK�!'�INS���w <B
U; �zH�NT���v�y�A `&| ��w�ΰP���쑜�����$���� ����2�=��=� '���SIO�e�1�  �XKC�IRTU�&@0�B�C�,SV� 2n�jp� ?X  Ф�(����͊@͉	������F@ �߀��>B�  =�[�5�a�s���������Tŕ=�d=�
ݐh�� ������6�X�$�n� W�8�P�b�|���ՒN� ����̯⯨����*� 8�f��n�X�����ҿ ����Ŀ���ڿ�� X�jτ�FϘϊ����� ߲����L�B�p�� ��b߸߮�x���6����H��7�I�X�	�MC: 567�8  Afsd�t1 78901�234q����  )y� �����c.��q�Y�'Q���`� l#�5�B�~P1�+�|�o������� ��������0'9 Rx_�����~�DMM P����A U�W�(F�Xj��POR 2]	 [�[���Z1F���B?��S4D 
!x�	/'���,/>/��v}?��B�l �e�)***@/�/#!{/�/��C�pONFIG� n����9�2[� e�$��/ّ�7  �z  D30h25Y��>�P0��e�C  C�3�h1�2D�D�/B42�3N �#� 2�,�Ӳ?o�?��:�ד�=���As!�=�O<O 3O��rO]OoO�O�O�O�O�O�O_� � :Z#S8_J_\_n_�_ �_�_�_�_�_�Y_!o oEo0oioTo�oxo�ot�o�I�� 3 [��`�g4 A�e�g ���01Bk!t�1C�`0.t���=#�
��Nn{k(EuK��Qu�LE@��eeu=D���qu��;��ʞ�u8I��u��It$ �$�m5@r�I���uFۀ3�uBQOGO�����t��+���E�.����Q���$�=�a�(4$�m�%��7�>�E���B<�~w����8E�y���;�j��ar�{�х>��݅���?s ���BHx�g!s >��� A!@��?E��qJ�b��@�sF��3{Fs�"��E~��b��vC��C��B��B ������j!AAo!k!�Bpp#B6q��f!Ju�@u�@�s @p0@�u�:p73� 	�	��l�c�u�����.pݑ Bo C��?����g ݯ��`?��33���a:�o-�?��a��c��� ����������ڿ�S?Ls�S�c�?8< ������B�����̻�p0%rk�a��8/x���
��<�>� -2��nπ�ߤ϶���e����߾�P�J�p������ �����V�A����@�� ��)qݑ��)r����� �������	��c�ѡo I��+�y����O�a� ��ڑ��)rk v�l��1��_FCCO�ORD 32 `!�?������ �r���
�= �d&�J|� ��/��*/�]/ /2/�/F/�/j/�/�/ �/�/#?�/�/J??}? 0?R?�?f?�?�?�?�? �?�?CO�?OjO,O�O POrO�O�O�O�O�O_ _�Oc__8_�_L_�_ p_�_�_�_o�_�_>o $oo�o6oXo�olo�o �o�o�o7�o^ D2�Vx��� ��$��W�
�<�~� d�R�Ïv���ꏬ�� Џ�D��w�*�\��� ��r�㟖���
�̟=� ��d�&���J�|��� �������د*��]� �2���F���j���޿ Ŀ��#�ֿ��J��}� 0�RϤ�f��ϊϼ��� ����C����j�,ߝ� P�r��߆��ߪ���� ���c��8��L�� p����������>� $����6�X���l��� ������7��^ D2�Vx��� ��$�W
<~ dR�v���/ ��D//w/*/\/�/��/r/�/�/�/
? 3��$CC_FSIW ���>1��  % 6M81Y<w? �?�4