��   C��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN��/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER��q�C_GRP6�P L$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� )DEX� �5O n�8BUF�7TDP�HG�_@FO�SxAV��7R?EC_TRQX��MFLG�J5�� � � N IU�
@!(UF*����4OSV3EN_CG"��0_�!�AU�SCH2�SMP]L4PEXE���2�!_�SUR}A�`jAaW�@A@bVNE|Y]QnAVA?�UY�T7D�VWWnAF�[V�A�\�WTO�0oH
e7D�f�3
e�U
e�W QT�P�0IR	 DMM��A@  @ �$la�EREG_�OFS�aME�hA1SS1�A !la�RE-   �# �0�b{F�c{ĥd� M�d�b�c$�STD�hq�gFA � �h!q�g�"�f�"�c�/ la7   �$p`TIN�@��0SUL� �R}_@  $}�@ SW@�rO:}rR%	 dp~t� �@JU� �s��FS4D6
 �' $�0PGF`QC?!$FIL� �@�E�PmA�s&�sDIG4o@SCA��$�INTTH�RS_BI�AZ�S�MAL%�COL���qATE_TI�PROG�4U�s��!CMDA�FSO�UTENV6�P $HRZ_kAXl�CU3VR2QALB܊�0��H�������PNT_M_V_AVR�CS!p9Lkp�c$L���f�O�\��ST�d�Fν#STO v�FX>�LECTEDCp��Y{���FY��t�ZL{�ړFZc�R�eȂ�	�/ G#P�oX $��_IVL����$!0B"�0�?0F�CCBDD�N=�CCIc�DU�MMY23G ^�DGEBU�A\!4PN�"TO�q9RP"� Q09T�6�� �;!��fBUT	TSP� ~@�q֥�E40N ڡFS3�ՁKQ1�r9T�I~�NEW_UI��VKP?Up`���CCOORD8\T�CH���01P��������7 l ��!�3$WEgIGH���2 s�_�aF��T��WAx{Q����NTER�Q���- ޵� �c���A�S0�$JZASTA�� �a��� T�,�26�36�W��!Ƨ ��ä"C��X�w�Yw�Zw�_�CM���?��D��i�RSLy�u���~��ƎŨ�ƚĆ�_Ϡ_ҡT   E0|c"0VROUNDCMVPERIO���$F1PUU3F2D�'TM1� �S��_DcGAMM�c1b�TRX�UKjt�K�K��CL�`��&O00ADJ�GA�UPDC0R"��יE� QRED���F#R_� _@W۲�x�u�DL_R��L@�=�M_�5d�0n� �#��}�"��}��k� ����������}�VLj�"����A�7���`��L�P5A8@� 
D�A�����"���y"��VIBƦ�OV��DEH�֌��` ,����*�� � R�TZ�MN1SUfM;N2YUFRAq	 ��ShZA
`-G���cOR�P�ҡAL�ҤCJ��
L���"�S8B�I$�L .$M"Pp30+�Q )�k�}�S"PHCD��GVz�GV��GVړJDO°]��]S�$R�E��h�b�]�A�AP)��DA��3$VF������1LVu��@IL�A���� #�� " �@fR!��$�DC+��Ԇ��B #П�5OBOA@�vYԣW2�G'	�$�ԍ$!#���E�K�`�+�eCNPRGOV6��%'P�t�_TW,��"G�3E�MNV�6c04�WT�cW�TRL_�SKIj�J�qcN���GW6�
eR<E�NABF��rV!� A$SB}��xS���{P�t yR*�tX�yRQT$���2_Q��?p����ALARMSERܟQETOTDFR�ZCHK1����62�9NC�4N@�5L`@N@�:vJ��vE�22�;�2�=NA9E�FFIXD2��BF�䦠@I�dD���DON�t�95P�SFW�0_DF1"%BF2/_vJ��|���4|�Pl��33=� �5|�kH|�yJ�Z��U
�23�;3�=|�9E�SDIAu �6�RKq�B��VvEfvC�3G	A�@�@���R<iV1 <d��sP�VQ�U�Uf��S$��� ��FU��ED�S_HA��U�e�d�4GE F�k@�2�`�;�a��5 !%�UzKq�#�X���s���Y��aw��@rSIW�_ � *�X��RK��`H7p_C�HCK�!'�INS����w <B
U; �zH�NT���v�y�A`& | ��w�ΰP���쑎Φ� �$���� O���2�=�=�s '���SIOe��1�  {XKC�IRTU&@�0�B�C�,SV �2n�� X  �P������͊@͉	��<����F@ �߀|��B�  =�[�5�a�s����������ŕ=�d=�
ݐh ��������6�X�$� n�W�8�P�b�|���Ւ N�����̯⯨���� *�8�f��n�X����� ҿ����Ŀ���ڿ� �X�jτ�FϘϊ��� ��߲����L�B�p� ߔ�b߸߮�x���6����H��7�I�X��	MC: 56�78  Afs�dt1 78901234q����/  )y� ������.��q�Y�'Q���`� l#�5�B�~P1�+�|�o����� ����������0' 9Rx_�������DMM P����A U�W�(�FXj��POR �2	 [��[��Z1F���B?��S4D7 
!x�	/�'��,/>/��v}?��B�l �e�)***@/�/#!{/��/�C�pONFIoG n���_9�2[�� �$��/ّ��7  �z  D�3025Y��>��P0�e�C  C�3�h1�2DD�/B4�23N �#� 2�,�Ӳ?o��?�:�ד�=���As!�O <O3O��rO]OoO�O�O��O�O�O�O_�� :Z#S8_J_\_n_ �_�_�_�_�_�_�Y_ !ooEo0oioTo�oxo�o�o�I�� 3> [��`h�g A�e�g ��bBk!t�1C�`0�.t��=#�
��N�nk(EuK���QuLE@��eeu=�D��qu��;��=ʁu8I��u��/It$ �$�m5�@rI���uF��3�uBQOGO��x��t��+���E��.���Q���$�{��a�(4$�m��%�7�>�E���B�<~w����8E�=y��;�j��ar���х>��݅��?s ���B�H�g!s >���B A@��?E��qJ��b�@�sF���3Fs�"��E�~�b��vC���C�B��AB������j!AAo!,k!�Bpp#B6q���f!u�@u�@�s @p0@�u�:p7 3�	�	��l�c�u���`�.pݑ Bo C��?���g ݯ��`�?�33���a:�o-�?��a��c� ������������ڿ��?Ls�S�c~�8< ��0����B����� ̻p0%rk�a��8/x���
��<� >�-2��nπ�ߤ϶���e����߾�P��J������� �����V�A����@� ��)qݑ��)r��� �·������	��c�� �oI��+�y����O� a���ڑ��)rk v��l�1��_FCCOORD 32 `!�?����� ��r���
� =�d&�J| ���/��*/� ]//2/�/F/�/j/�/ �/�/�/#?�/�/J?? }?0?R?�?f?�?�?�? �?�?�?CO�?OjO,O �OPOrO�O�O�O�O�O __�Oc__8_�_L_ �_p_�_�_�_o�_�_ >o$oo�o6oXo�olo �o�o�o�o7�o ^D2�Vx�� ���$��W�
�<� ~�d�R�Ïv���ꏬ� �Џ�D��w�*�\� ����r�㟖���
�̟ =���d�&���J�|� ���������د*�� ]��2���F���j��� ޿Ŀ��#�ֿ��J�� }�0�RϤ�f��ϊϼ� ������C����j�,� ��P�r��߆��ߪ��� ����c��8��L� ��p���������� >�$����6�X���l� ��������7�� ^D2�Vx�� ���$�W
< ~dR�v��� /��D//w/*/\/ �/�/r/�/�/�/
? 3��$CC_FSI�W ����>1� K  6M81Y< w?�?�4