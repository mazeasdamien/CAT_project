��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1RTU4QQ�Rx1R�� � $TIT91� ��� �Td��T0�ThP�T5�V6��V7�V8�V9�W0 �W�WOQ�U�WgQ�U�WU1�W1�W1�W1�W�2�R!SBN_CmF�!@$<!�J� ; ;2�1_CM�NT�$FLAsGS]�CHEK"{$�b_OPTJB� � ELLSETUP  `@�HO8@9 PR�1%x�c#�aREPR�hu0D+�@��b{u[HM9 MN�B;1^6 UTOBJ U��0 49DoEVIC�STI/@��� �@b3�4pBܢd�"VAL�#IS�P_UNI�tp_�DOcv7�yFR_F�@|%u13��A0s�C_WA�t,q�z�OFF_T@N�DEL�Lw0dq�1��Vr?^q�#S?�o`Q"U�t#*�Q3TB��bMO� �OE � [M������REV�B3IL���!XI� v��R  !D��`��$NOc`M�|����ɂ/#ǆ� ԅ��ނ��@Ded p �E RD_E��h��$FSSB6�`K�BD_SE�uAG*� G�2Q"_��2b�� V!�k5p`(��C��00q_ED� �� � t2�$!SL�p-D%$� �#r�B�ʀ_OK1��0] P_C� ʑ0tx��U �`LACI�!��a�Y�� �qCOsMM� # $D
�� ��@���J_\R BIGALLOW�G (Ku2-B�@�VAR���!�AB  � �BL�@� �C ,K�q���`S�p��@M_O]˥���CCFS_UT��0 "�A�Cp'���+pXG��b�0 4�� IMCM ��#S@�p�9���i �_��"t�����M��1 h$�IMPEE_F�s��s�`�� t����D_������D��F�����_����0 T0@L��L�DI�s@�G�� �P��$I�'��%w�CFed X@�GRU@��Mb�N�FLI�\Ì@UI�RE�i42� SW�ITn$`0_N�`S� 2CF�0M� �#u�D��!��Pv`����`J�tV��[ E��.p�`�ʗELBOF� �� ��p`0���3����� F�2T��A`�rfq1J1��z _To!���p��g���G�� �r0WARNM�p#tC�v`�ç`\ � COR-Ur�FLTR��TRA�T9 T%p� $A�CCVq��� ��r�$ORI�_&�ReT��S<���HG�0I���TW��A�UI'�T�M�K�� �202�a1�N�HDR�2��2�2�J; S���3��4���5��6��7��8®�9KD׀
 �2� @� TRQ�$�vf��'�1�<�_U�<�G��Oec  <� P�b�t�53>B_�LLEC��!~�MULTI�4�"u�Q|;2�CHILD���;1���@T� "'�STY92	r��=��)2�������ec# |r056$J� ђ��`���uT�O���E^	EXT�t����2��22Q"�0����$`@D	0�`&��p����� (p�"��`%�ak�����s�@���&'�E�A�u��Mw�9 �% ���TR�� ' L@U#9 ���=At�$JOB���мP.TRIG��( dp������^'�#j�~�-_MO�R�) t$�F�L�
RNG%Q@�TBAΰ �v&r�*`1�t(��0 �x!�0�+P��p�%4��*��@͐U��q�!�;2J�S_R��>�C<J�T8&<J D`5CF9����x"�@?��P_�p�7p+ \@RaO"pF�0��IT�s�0NOM��>Ҹ4s(�2�� @U<PPgў�P8,|Pn��0�1P�9�͗ RA���pl�?C�� �
$TͰ.tMD3�0T��pQU�`�΀+AHlr>�T1�JE�1\�J����PQ��\Q��hQCY�NT�P��PDBG�D̰�0-���PU�6$$Po�|�u�AX�����TAI�sB�UF,�3�A�1. �����F�`PI|�U-@PvWMuXM�Y��@�VFvWSIMQ�STO�q$KEE�SPA��  ?B�BP>C�B�A��/�`�ˏMARG�u2�F�ACq�>�SLEW�*1!0����
�WQ_MCW$0'���p�JB�Ї�qDEC�j�eN"s�V%1� Ħ�CHNR�MPs�$G_@�gD��_�@s��1_FP�5�@TC�fFӓC�� ����qC��+�VK�*���"*�JRx���SE7GFR$`IOh!�0;STN�LIN>�csCPVZ��R�A�D2�� ��r 2��hr�rcb��?3` +^?�� �եq�`��q|`����p�t��|aSIZ#�!� �T�_@%�I��qRS�*s��2y {�Ip{�pTpLF�@��`��CRC����CCTѲ�Ipڈ�a���b��MIN��a1�T����D<iC �C/����!uc�OP4�n j�E�Vj���F��_!uF��N����|a��=h?KeNLA�C2�AOVSCA�@A�Up�r1�4�  �cSF�$�;�Ir ��3�a�05��	 D-Oo%g��,,m�����ޟ�N"RC�6� n���sυ��U��R�0HANC���$LG��ɑDQ�$t�NDɖ��AR۰N��aqg��ѫ�X��ME��^�Y�[PS�RAg�X�AZ�П���:rEOB�FCT��A���`�2t!Sh`0ADI��O��y�s"y�n!@�������~#C�G3�t!��BMPmt@�Y8�3�afAES$���v��W_;�BAS#?XYZWPR��*��m!��	VQU�87/  ƀI@d��2�8\�p_C:T����#1R_L
 � 9K ���C�/�(z�J�LB�$�3�xD��5�FORC��b�_AV;�MOM$*�q�SaԫBP`Ր� y�HBP�ɀE�F�����AYLOAD&$�ER�t&3�2�Xxrp�!u�R_FD��_ : T`I�$Y3��E�&��Ct��[MS�PU
$(�kpD��9 �b�;��B�	EVId�
��!_IDX2$���B@X�X<&v�SY5� %��R_HOPe�<��ALARM��2W�s���0= hb Pnq�`M\qJ@$PL4`A&�M#�$�`���� 8�	���V�]�0���1U�PM{�U��>n�TITu�
1%�![q�BZ_;���? �B pQk��6�NO_HEADE ^az��}ѯ��`􂳃����dF�ق�t���@��@��uCIRT�R�`��ڈL��D�ClB@4�RJ�� �[Q����A�2>���O�R�r��O����T`UgN_OO�Ҁ$����T�����I�VxaCx�PXWOY�z��B��$SKA�DR�ADBT�TRL��C��րfpbD�s��~�DJj4 _��DQ}��PL�qwbWA���WcD�A��A=�2��UMMY9��1!0�+����D;[Q;PR�� 
MМZ���E O�Y1�$�a$8�9��L)F!/_c���0G�G/��p�PC�1H�f/���PENE
A@Tf�I�/��M$��COR`"JH y@ �E$L�#F$#PR���+jp���nq�_D$�qPROSS]�
���R�r�` >u�$TRIG96�PAUS73ltETgURN72�MR:�eU 0Ł0EW$�~�SIGNALA��QR$LA�З5�1�G$PD�H$PDİ�AI�0�A�C�4�C��DO�D�2�!��6GO_AWAY2MOZq�Z�W �DCS��CSCB�g�K Իa#���E+RI�0Nn�T�`$�����FCBPL�@QBGAGE���P��ED`|BD�wA[CD�OF�q�[F0�FoC��MPM�AB0XoC�$FRCIN��2Dk��@��O$NE�@�FD�L8�� L� �����=��Rw�_��P>� OVR10����lҠ�$ESC_|�`uDSBIO��p��pTe�E�VIB�� `s��Z��V��p�SSW��$�VL��:�Lk��X���ѣ�0bQ����USC�P��qA=�	Q��MP1%e@&S*`�(bt`'c5۳ESUd��-cWg&S Wg?cWd����Wd��Wd<.���AUTO$�Ya҃�ac�SB����-d���&SwB[��GB�f_$VOLT�g ���  �GAOD!��q���@:�ORQ�ҀKra�$DH_THE&0�Rgp� <qtnwALPHnt��o��w0 Vp]�$�.�Ra�[��s�5�`r�CQ�#BUD�S� F1M���sV
��;��L�b�tk���BRTHR��L��T`�Z���Vɖ��D)E  �1��2�⋅ ��������kѯ�a� �Tt0V�ꆸ������@̈Я�-�"�N~���sS2����INHB��ILTG0ɡ�T?� �3$�w��E��PqQxQ��TqPe��0Y�AF}�O�ນ��ڗ ��qPڳē����bPܙ���PL?���3���TMOU��ēS��� � ��s�/�S18���O��Aܙ��I����CDqIƑ˩o�STI��գ�O:ҋ�,0���AN��Qg�S��+r�#x$�����w�1_����PRA�P`�vC����MCN�eQe�����VER�S��r�oPIw�F�PåǲШ۷G.�DEN��G>�����F�2H�Ƿ�M�7�F��_�MN�D̠,���@�d�{ƭa����OB����U˱z���DI ���#���3�����A��w�Fx���3�O�N�5��Q��VAL��CR[�_SIZp��b�;Qn�REQ�R�b��]2b���CH q�΂�ڃ�Ռ�����:�n�S_U��X��wW�FLG���wU$CV�iMGP�QδFLXP�923R�u�L��EAL�P-�C	��+rT��W��� �R��c���NDMS�7� ��K>S�P_M'0h�STWv������AL�P���Q����U���U�IAG@,�o��d�U�-�T"	A-`� ���A��� ��H`��Q`��6��Pq_D&��1s��.�P��F�>2�T�� ?7 1A>���#�#L��?`_=i @@>LD�pc���0�FRI�0 `Ѐ��1}Ѳ�IV\1�*�^1�U�P`��a��C�L!W��
`L=S&-c&&S�C.w��  L���!����d�Q$w!�҇��$w��p��
�P�5RSM��P���V0h � r�l�d^2AW�a_TRp�}�8@NS_PE�A����< ��$�SAVG�8�6G]%���CAR �`�!�$���"CRa���$ d�#qE�@��"STD���!Fpo��'QOF0��%��"RC���&RC۠�(F�2A�R#7����%, gMA�Q_�a��
QQ��al2��%u4Ib�r7I�R�9�wQ�7�8M/��!C:pR�  �p�2F<�SDN�a0 �  W2QM P $Mi��s$cA �$C�cm�9���4���AT�0CY_ �N LS!IG1@x'yB��y@@H2Y��NO����SDE�VI�@ O@�$�RBT:VSP0�3�CuT�DBY|�A�	W`3CHNDGD�AP H@GRP�HE iXL�U��VS��Fx2��CL1p �Q6ROp��FB�\]�FEN�@��Sp��ChAR d�@�DOd�PMCS�b�P薇P�R��HO�TSWz42�DMpELE�1/e� D8`�RS T�@���r� hfl��`OL�GHA�Fk�Fs��|�C�A@�T � $MD�LUb 2S@�E ���q�6�q	0�i�c�e
�cJ��	uݢ�#~X5t+w�PTO��� x�bHe DSLAVS�� U  ��INAP �	V�ЊyA_;�wENUAV $R��PC_�q�2 1bLr�wﰦtSHO+� W ���A�a�q��2�r�v�u�vNc_�CF� X`c ,f��r�OG g`E��%D�h�{PC�Iߣi�MA��D�x �AY?�W� p�NT�V	�D�VE�0@�SKI��T�`g?Ň�2�� JZs�! Cpꆻ��f�_SV/ ��`XCLU��H�N��ONL��'�Y�T���OT:eHI_V|,11 APPLY���HI4`;�U�_ML��� $VRF�Y8�	�U�M{IO#C_I���J 1/��2߃O�@X�LSw"`@�$DUMMY4����ڑ�Cd L_�TP���kC��^1CNFf���E��@T�$y� D_#UQ_��ݥ�YPCP��=�� ������aD���� �Y +�
0RT�_;P��uNOC�Cb Z�r�TE ���=�פ DG�@�[ D�P_BA�e`kc�!$��_��H��d���E \�p�Ab=cARGI�!�$���`[ B�S;GNA] ��`U��IGN�Տ��� ���V������ANNUN��&�˳�ExU�J'�ATCH빀�J���4�rA^� <@g�����:c	$Va��������AEF] I�� �_ @@FͲIT>b�	$TOTi �C��O�c�u�M�@N�I�a`tB��c�r��A>���DAY@CLOAD�D\�n��~�� �EF7�+XI�Ra��K����O%��ap�ADJS_R�!@b��>�H2�"[�
 c�%��`�a͠MPI�J��D��A��?�Ac 0@��х�� ��Z�ϡ��Ui ��CTR�L� Yp d��T�RA8 ?3IDLE_PW  �Ѡ��Q��MV�GV_���`c�q�p�;Q@e� 1q$��6`<cTAC-3@��P�LQ�Z�Rz�\ A-u:ɰSW;�A\���/J��`�b�K�OH�(OP9P; �#IRO� �"gBRK��#AB � �O������� _ ���F���`d͠, j@S�oRQDW��MS��P6X�'z��IFEgCAL�� 10^tN��V��豊�V�(0L��CP
��N� 9Yb�0FLA_#�3OVL ��HE���"SUPPO��ޑ\B�L�p��&2X�*$Y-
Z-
W-
��`/��0GR�XZ�q6�$Y2�CO�PJ�SA�X2R��*r�!���:��"�BI�0)�f{ `�@CACHE���c��0�s0LA�Z SUFFI, �C��{Q\���6�o��1MSW�g �8�KEYIMA-G#TM�@S��n�
2j�r��%�OCVsIE��~�h �a�BGL����`�?�P@��@���i��!`STπ!�����������EMAI�`N��`A @Z�'FAU� �j�"{Qa��U�3��� �}�k< $dI#�US�� �IT'��BUF`��DN�B���SUBu$�DC�_���J"��"SAV �%�"k������';�r�P�$�UORD���UP_u �%��8OT�T��_B`��8@LM0l�F4��C7AX@Cv�b��Xu 	��#_G��
c@YN_���lT6���D�E��M��U��T��F��cavC�DI`BEDT)@IC��~�m�rI�G�!"c�&��l`��-�P���FZP n (�pSV� )d\�ρ�����B��o� �����>"$3C_R�IK��kB��hD{p�RfgE.(ADSPd~KBP�`�IIM�# �C�Aa�A��U�G��4�iCM! IP��KC��� �DTH� �S�B2*�T��CHS�3�CGBSC��� ��V�d�YVSP�#[T_DrcCONV�Grc[T� $�Fu F�ቐd�C�0�j1��SC5�e]CM�ER;dAFBCMP;c@ETBcF�\�FU DUi ��+�~�CD�I%P70�2# �EO���qWӏ�SQ��QǀSU���MSS�1ju�4`�T�aAa��A�1r�� "�Й��4$Z!O@s���l�U6�&�2�eP���eCNc�l�x�l�l�iGROU�Wd)��S c�MN�k Nu�eNu�eNpR|b|�i��cH�pi��z
 �0CYC���s�w�c�6�zDEL�_D��RO�a���qVf���v{�O�2���1��t���:R�ua�.#� ��A	L� �1sˢI1¡�DJ0�PB���>aR^�9T�Gbt ,!@���5��aGI1LcR1s3 
��ԠNO��1Au���������P�����Cڠ	�������1��J0�0vH *	�LU�1#J�Q��V 
�[�7Az���z��z�@�z��z�Fz�7w��8w�9w���y���1���1��1��1��1�Ě1њ1ޚ1�2R��2����2��2��U2��2Ě2њ2ޚU2�3��3��3�����3��3��3Ě3*њ3ޚ3�4���bXTF��1w6�.(�0@�f�0�U�0ŷ�e���FDR5�xTU VE��?1���SR���RE�F���O�VM~C)�A2�TR�OV2�DT� R�MXa�IN2���Q�2�'INDp�r�
���0�0�0Gu1��[�G`��r{�D_�[�RIV�P���GEAR~AI%Or�K"N�0��y�p�5`@�a�Z_�MCM� �����U�R�Ryǀ��!?3 ��p?nЋ�?n�ER�vт�H�!�P��zI:�PXq�B�RI0%��#E�TUP2_ { ���#TDPR�%�TBp�����Վ��C��2| T��"�4)��:%	`^B��p�I+FI��� Mc����.�PT���FLU=I�} � ��K UR�c!���B�18SPx E�EMP�p�2u$��S^�?x��qJق0
3VRT����0x$SHO��Lq�6 ASScP=1��PӴBG_���-�����FOcRC:dh�d~)"KFUY�1�2\�2
Ap�1h� p� |��7NAV�a��������S!"��$VgISI��#�SCM4CSE����:0E�V�O��$���G@���$��I��@��FMR2��� �5`�r�@ �� �2�I�9 F��"�_���LIM�IT_1�dC_L�M������DGCL�F����DY�LD����5������� �����u	 T��FS0Ed� P�QC�0$EX_QhQ1i0�P�ajQ3�5��GoQ���� ����RSW�%ON�PX�EBU1G��'�GRBp�@mU�SBK)qO1L�7 ��POY 
)P��P��M��OXta`SM��E�"�a����`_E � �
@��TERMZ%�Nc)ORI�1_ �c%��SMepO��_ ��c%DMA��`�(��c)UP>� �g� -���b����q#� ���G�*� E�LTOQ�p�0�PFIrc�1Y��P�$�$߆$UFR��$��1L0e� OT�Y7�PT4q�k3NS]T�pPAT�q4OPTHJ�a`EG`8*C�p1ART� !5p� y2$2REL�:)ASHFTR1�1��8_��R�Pc�& � $�'@�� ��H�s�1 @I�0�U�R} G�PAYLO�@�qDYN_k���.bp�1|��'PERV�� RA��H��g7�p�2�0J�E-�J�RC����ASYMFLTR��1WJ*7����E �ӱ1�I��aUT�p bA�5�F�5P�PlC��Q1FOR�pMH�I!���W��/&8�0F0�b�H��Ed�� �m2N���5`O�C1!?�$�OP����c��X���bRE�PR.3��1a�F��3e��R��5e�X�1(�e$P�WR��_���@R_`�S�4��et$3UD�Ҹ���Q72 ����$H'�!�`ADDR�fHL!G�2�a�aʛa���R��U�� H��SSC����e`-��e���e��SEE���HSCD���� $���P_�_H B!rP�����_HTTP_��HU�w� (�OBJ�l�b(�$�fLEx3��PWq�� � (���ะ_��T?#�r1S�P��z�KRN�LgHIT܇5��P���P��r������PL��PS�S<�ҴJQUER�Y_FLA 1�qB_WEBSOC��G�HW�1U���`}6PINCPU���Oh��q����d����d�����IHM�I_ED� T ��RH�?$��F�AV� d�Ł��IwOLN
� 8��yR�@$SLiR�$INPUT_�($
`��P�� �ـSLA� ����5�1��C���B��IO6pF_�AS7��$L%�}w%�A��\b.1`�����T@HYķ촑���؁_UOP4� `y�ґ�f@�¤�������`PCC�
`����#���aI�P_ME�񵁗 �Xy�IP�`�U�_GNET�9���Rpĳs�)��DSP(�Op=��BG�p��9M�A��� l�:C�TAjB�pAF TI��-U��Y ޥ�0PS6ݦBUY IDI�r F ��P��q�� �y0�,����Ҥ��NQ�Y R��IRC�A�i� � �ڛy0�CY�`EA �����񘼀�CC�����R�0�A�7QDAYy_���NTVA�����$��5 ���SCAd@��CL����t���𵁛8�Y��2e�o�N_�PCP�q��ⱶ��,�N����
��xr���:p�N� 2� ؀��(ᵁ����xr۠LABpy1��Y ��UNIR�9�Ë ITY듭�$�e�R#�5����R_URL���$AL0 EN��ҭ�t� ;�T��T_U��ABKY_z��2D#ISԐ�C�Jg����P�$���E��g�R��З A�/���J����FLs��7 �Ȁ���
�UJR.� ���F{0G`��E7��J7 �O R$J8I�7���R�d�7��E�8�{�H�APHI�QS��DeJ7Jy8B��L_KE*п  �K��L}M[� � <X��XRl�u���WATCH_VA��o@DўtvFIELc��cy3����4� � o11Vx@��-�CT[�9��m��PLGH���� $��LG_SIZ�t�z�2y�,p�y�FD��Ix��� +!��w�\ ����v��S ���2��p��������\ ���A�0_gCAM]3NzU
RFQ�\vv�d(u�"B��2�p����I��+ �\ ���v�RS���0 } �ZIPDUƣ�p�LN=��ސ �p�z6���f�>sDr�PLMCDAUi�EAFp���TuGqH�R��|�BOO�a?�� C��I��IT+���`��RE���SCR� �s���DI��SF0�`RGIO"$D�����TH("�t|�S�s{�W$�|�X��JGM^'MgNCH;�|�FN��ba&K�'uЅ)UF�(�1@�(FWD�(HL.�)STP�*V�(%�X�(��(RS9HIP�+��C[T�# R��&p:'^9U=q�$9'�H%�C𜓚"Gw)�0PO �7�*��#W}$���)�EX��TUI�%I ���Ï���rCO#C�� *�$S��	�)��B@�NOFAcNA|��Q
�AI|�8�t:��EDCS��c��C�c�BO�HO�GSȅ��B�HS�H(IGN�����!O���D�DEV<7LL���Z���­Ц(�;�T�$��2�p�����*�#A���(�`뀸{�Y��POS1�U2��U3�Q��1R�A�Ш# ��{�PtD�� ��&q)��0�d��V+STӐR�Yl�B@~ ` �$E.fC.k�p<p=fPf��4�ѩ LRТ� �� x�c�p��<�Fp�d/�@!�_ � ���7Lp&���c�{MC7� ���CLDPӐ��TR�QLI#ѽ�ytFAL��,r�5s8�D�5wS�LD5ut5uO�RG��91HrCRESERV���t���t��c�� �� 	u95t5u��PITp��	xq�t�vRCLMC�������q&�M��k�������$DEBUGMAS��ް��?%U8$T@��Ee�g�ޥ�MFRQՔ�� � j�HRS�_RU7��a��A<��k5FREQ� ��$/@x�OVER���n��V#�P�!EFI�%�a��g�8,S���t� \R�ԁ�d�$U�P��?��p�PS�P��	�߃C��͢a��U�\�l�?(P��PMwISC� d@��QRQ��	��TB� � Ȗ0A՘A�X����ؗ�EXC�ESjҧ�M��\���W�����oQ��SC>�P � H��̔_��Ƙǰ]������KHԳK�J� m�B�_K�FLIC�dB��QUIREG3M�O��O˫3�q�ML:�`MGմ �`���T���aNDU�]��>��k�G��Df��INAUT���RSM>�a��@�N�r]3-��p5�PwSTL\�� 4X�7LOC�VRI%��U;EXɶANGuBu����� A���b�������MFO� ����Y�b@�e4�2�k�SUP�eQ�FX���IGG� � ��p�c���cQ6 �dD�%�b|�!`��!`���|��3w�ZWa�TId��p�XPIN[��� t��MD��I��)֟@���H8ݰM��DIA��ӂ��W,!�wQ�1�D��);�O���]��[ 0�CU��VP�(�pu���O!_V���� ���S�X�5������P��0N���P��KES2����-$B� ����ND�2����2_TX�dXTRA�C?�/���M�|q�`�P�v��XҰ�Pt SB�q`�USWCS��Tx��	���PULS��A�NSޔ��R��JOIN��H��~`j�=��b��b�����P=��$��b$���TA����S���S�H�S�E��SCF�aPJ���R��PLQ� ���LO��н�.�������8�p�������RR2���� 1��eA^�q d$��Iΐ�+�G�A2+/� w�PRIN��<$R SW0�"�a/�ABC�D�_J%�¡��_Ju3�
�1SPܠ$e��P��3����`��J/���r��qO8QIF��CS�KP"z{�{�J���QL2LB�Ұ_AZ�r�~E�LQ��OCMP0ೕ�T���RT������1�+���P1���>@�Z�SMG�0��=�JG�`SCyL�͵SPH_�@���%V�� R�TER`  �< A)_�@G1"�A�@c̔�\$DI�
"23�UDF�}!L�W�(VELqIN8�b)@� _BL�@u� �$G�q�$�'�'�%`�<�� ECHZR/�TgSA_`����	E}`<����5�B��1}`_�� �@)5D2d%��A4I��N9�t&R�DH�A�����P$V `�#>A�$��ł�$�Q@�R}ӆ��H �$BELv�|��<!_ACCE�!�c��7/��0IRC_4] ��pNTT��SO$PS�rL� d�/Es��F{�@F 
��9gGCgG36B���_�Q�2�@�A��n�1_MGăDD�A]"łFW�`���3�E�C�2�HDE�KPP�ABN>G��SPEE�B�Q%_pB�QY��Y��11$USE_t��,`Pk�CTReT�YP�0�q P�YN���Ae�V)хQM���ѷ��@O� YA�TINCo�ڱ�B�DՒ8�WG֑ENC�����u�.A�2Ӕ+@INP�OQ�I�Be��$N�T�#�%NT23_�"łIcLO� ł_`��I�œif� œk��? �` ej�C400fMOSI�A���ОA����PERCH  �c��B" �g��c�� lb=�����oU�@�@	A�B(uLeT	~��1eT�ljgv�fTRK@%�AY��"sY� �q�B�u�s۰�]��R�U�MOMq�ՒY�M!P�Ĕ�C�s�C�JR��DUF �BS_�BCKLSH_C �B)����f���St�H���RR��QDCLAL�M-d���pm0��CH�K���GLRTY���d��Y��)�N�d_UM]�ԉC�p�A!�=PLMT� �_L�0��9��E �.� ��#E)�#H� `=��Q3po�xPC�a�xHW�頿EׅCMqCE��@�GCN_,1ND�Ζ�SF�1�iVoR��g<!��0r�n��CATގSH)� ,�DfY��f��7A����܀PAބ�R_	P݅�s_ �v���s����JG�T�]���Y�����TOR�QUaP��c�yPO�U��b��P%�_W �u�t��1D��3C��3�C�IK�IY�I�3F��6�����@VC"�00RQ�t��1���@8ӿ��ȳJRK���,��UpDB M��Up�MC� DL�1BrGRVJ�Cĭ3Cĳ3$��H_��"�j@q�CO1S~˱~�LN��� µ�ĭ0�����u��ʈ�̓��Z���f$�M�Y��؊���>�T�HET0reNK2a3�3hҧ3��CBm�kCB�3C! AS� ���u��ѭ3��m�SB8�3��x�GTS$=QC�����������$DU��Kw�B(�%(��%Qq_��a��x�{�K���b(��\�A`Չ��p�{�{��LPH~�g�Aeg�S µ��������g����(��֚�V��V��0���V��V��V��V���V	�V�V%�H���������G�����H���H��H	�H�H*%�O��O��OV	��UO��O��O��O��UO	�O�O�Fg�����	�����SPBALANCE_-ѶLE��H_`�S�P!1��A��A��PFULCElTl���.:1��UTOy_����T1T2��22N���29`�!@�qnL�=B�3�qTXp�Ov 
A4�INSE9G�2�aREV��`�aDIF�uS91�l8't"1�tpOB.!t�M��w2�9`��,�?LCHWARRCBAB�� ��#�`-�(�Q 5�X�qPR��&8��2�� 
�""���1eROB͠CR�0r5��0p�C�1_���T � x $WEIGH�PFrp$��?3àI�Q�g`IFYQ�@LAGĒRq�S�R �RBI�Lx5OD�p�`V2S�T�0V2P!t�W0 P�01�&1/0�30
�Px�2�QA  2řd^[6DEBUg3L_@z�2�MMY9&E� Nz�Drp$D�_A�a$�0��O� ���DO_:@A.1� <B0�6��m�Q�B�2�0ND-cdH_p`�P�3O�� �� %��T`"a��T/!�4)@�TICKh3| T1"1@%�C ��@N͠�XC͠R?��Q�"�E�"|�E8@PROMP�S�E~� $IR���Q��R;pZRMA�I)��Q�R4U_r0�2S; �q�PR8�C�OD�3FU�Pd6I�D_[�vU R!G�_SUFFu� �l3�Q;Q�BDO`�G �E�0�FGRr3 �"�T�C�T�"�U�"�UPׁ�T8D�0�B0Hb �_FI�19*cO�RD�1 50�23�6V�+b�Q1@$Z;DT}U	 �1;E��4 *:!L_�NAmA�@�b�EDEF_I�h�b�F�d�E �2�F�4�F�c�E�e�FISP��PAKp�Ds"�C�d��44בi�B�2D�"�It�3D��O#OBLOCKE z��S�O�O�Gq�R�PUM�U�b�T�c�T�e �T!r�R�s�U�c�T�d �R�6�q�S� ���U �b�U�c�S�Z��X�@�P` t�@qe�)@W��x���s����TE�<D�( }l1LOMB_���ɇ0V2VIS;�I�TYV2A��O�3A�_FRI��a SIq�QR�@��@R�3�3V2W��W��4����_e��QEAS^3�Rϡ��_�[p:R��4�5�6_3ORMULA_Iz����THR^2��EGtg�30f��<8�5COEFF_O�A�	 ��A��GR�^3S�g0BCAnO/C$ܐ�]3me�1GR�P� � � �$�p�YBX�@TM�~w���u�B�s��bCE�R, Tttsd�0� M �LL�TSpS~�_SVNt�ߐ���0q����0� ���SETUsMEA�*P�P��W0�1+b/0�� � h��   @ڐo�l�o�cqz��b��@cqq`tP� G��R�� Q\p*q[p趻>�c NPREC�>at�5@MSK_�$|�� PB11_USER�e"�p{ ���VEL�� �{ 0�$Ō!I]`�w�MT�ACFG����  �@@ O�"NORE-0l@o�V�SI.1�d��6�"�UXK�fP!��DE��� $KEY�_�3�$JOG��0SV������!��}�SW�"�a\a4S�ՐT|�GI�p`�| ^�� 4 ph��'d2�!XYZc����31�_ERR#�� 8Ԡ�AfP�V�d��1����$BUF��X����wMOR|�� HB0CUd�lA�!��GQ\axB�,"!a$� ����a��u��?�G�~�� � $S1IՐ���VO��T��0OBJE_��A�DJU)B��ELA�Y���%�DR�OU�.`=ղВQ0b=���T���0���;BDIR���; I�"0GDYNW�2��T���"R���@�0�"�O�PWORK���},%@SYSBUy���SOP��ޑ��U�; P�pN�<�P�A�t�>�"��OP��PUd!0�`!��^l�IMAGw�B0�y�2IM�Õ�IN�e�d��RGOVR!D��-��o�Pq��@0��J�Os���"L�p�Ba���o�PMC_QEe`���1Ny M� A�21�2T���SL�_��� � $OVSL�ǫ�?q�`"��2�" -�_��k �P��k�Pu���2�C� �`�Ź���/_ZER�D��w$G�� 2=���� @*���%MO~PRI��� 
�JP8+��=!/�L���ح�T� �0AT�US��TRC_T���sB��}fs��9s�1Re`��� DFAm����L���"��00a� ޱ��XEw{�����C0vcUP��+p	qPXPȝj�43 �e��PG\���$S�UBe�%�qe9J?MPWAIT z�}%LO��F�A�R�CVFBQ�@x"�!R��� �x"ACC� R�&�B�'IGNR_{PL9DBTB�0Pqy!BWbP�$w��Uy@�%IGT�PI���TNLN�&2R���rL�NP��PE�ED \HADO!W�06�w��E[q4�jO!�`SPDV!� LbAz�`�07��3UNIr��0"!R��LYZ`� o}�PH_PK���e�RETRIE�9{�q�/�0'PFI"�� �G`�0D� 2�g�DBG�LV�#LOGSIYZ��EqKT�!U��2VDD�#$0_T�G��MՐCݱ��|@eMR�vC}�3�CHECK�0���0O�V!�k��I��LE(!��PA�rpT�2K�W�@IP�2V!� h $ARIBiR� c�a/�qO�P8�ӐATT�� 2�IF|@z�Aq4S�3�UX����PLI�2V!� $g���I�TCHx"[�W �A�S9�wSLLB�V!�� $B�A�DYs��BAM�!���Y9�PJ5Ƚ�Q��R6�V�Q_KGNOW�Cb��U��#AD�XV��0D�+i?PAYLOAt��BIc_��Rg�RgZOc�L�q��PLCL_�� !7��b�Q�B��d���fF�iC�֠�js��d�I�hR�ؠ�g�ҢdB����JL��q_J�a���AND��Ĳ.t�b�a�L!q�PL0AL_ �P�0���Q�րC��DNcE���sJ3CpWv� TPPDCK������P��_ALPHgs�sBaE��gy|��K�|1�� � ����HoD_1Oj2ydDP�AR�*��;�&�^��TIA4U�5U�6��MOM��a����n���{�Y�B� AD�a���n���{�PUB��R��҅n�҅{�/�2�Wp��W �  �PMsbT� �@xQ���� e$PI��81�@�TgJ��niJ�IV�Id�Ir��[��3!��>!��r�Ӫ�U3HIG�SU3�%�4 얎4�%� ���"�����!
��!�%SAMP ���^��_��%�P4s ю���[ 	� ��3 ���0���&���@����^��Sp��H&0	�IN�SpB�����뤕"��6��6�V�GAMM�SyI�� #ETْ��;�D�tA�;
$ZpIBR!62]IT�$HIِ_��H����˶E��ظAҾ���LWͽ�
���@7���rЖ,0�qC�%�CHK��" �~I_A�����Rr �Rqܥ�Ǚ��ԥ��ɾWs �$�x �1���I7RC�H_D�!� RN{��#�LE��ǒ!�,��x���90MSWsFL�$�SCR((G100��R@��3]B ��ç��a����َ0���PI3A9�MET�HO����%��AX�H�XX0԰62ESRI��^�3��R�0$u	��pF{�_���I?ⲣ1�L�L�_�a�OOP����wᜲ���APP:���F����@{���أRT�V�OBp�0T����;��� 1�I��� ���r���RA�@MG�A1���SSV�-��P_@CUR�g�;�GRO[0S�_SA�Q��Y�#NO�pC!"�tY� �Zolox�������!bX����&�DO�1A�� �A����Х��A���A`"�WS�c L"|h�*�� � �ãYLH�qܧ��S rZ�]B�o�=�q(�õq_�C1��'M_W���g���c�M� �`Vq��$p�x1o�3"�PMJ�,�� �'A� 9��!Wi:�$�L WQ|ai�tg�tg�tg{t� �N`���S���SpX�0O�sRqZp��P� *�� ���M������������@��X��� ��@BL�q_~R� |�q#(Y� ���&n��&{�Y�Z��'0�&t��Q�� !��"N0�� ��&P#Q��PMON_QU�c� � 8�@Q�COU��%PQTH��HO�^0HYSf:PES�R^0UEI0tO�@O|T�  �0�PGõz�RUN_TO�K�0ْ.�'� PE`�5C��A�<�INDE�ROGGRAnP� 2g��NE_NO�4�5I�T��0�0INFO�1� �Q�:A���'�OIB� (��SLEQݖFAѕ�F@�6�@OSy�T�� 4�@ENAB|��0PTION.S%0ERVE���G���wFGCF�A� @bR0J$Rq�2����R�H�O�G��EwDIT�1� �vR�K�ޓʱE�sNU0W*XAUTu�-UCOPY�ِN\����MѱNXP\[qƯPRUT9� _RN��@OUC�$G��2�T&��$$CL�`?0��&�������� �P�Sܛ@�X�PX=K�QIRTU��_��PA� _WRK �2 e�@ 0  �5�Q�MoYhJo|m �|l	�`�m�o��`��o�o�f�e�l}��aI[ct'`BS��*� 1�Y� <7�� �����&�8�J� \�n���������ȏڏ ����"�4�F�X�j� |�������ğ֟��� ��0�B�T�f�x��� ������ү����� ,�>�P�b�t�������켿srCC��LMT�?0���s  d�ѴINڿ�дPR_E_EXE��)��Ƅ0jP��za'`D�V��S�@e)��%select?_macro�����kϤ�qtIOCNV�VB�� ��P��U�Sňw���0V 1]4kP $$p��a0�|�`?���߰ >�P�b�t߆ߘߪ߼� ��������(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L ^p�������� ��$�ѰLAR�MRECOV �^�����LMD/G �Ь��LM_IF ���d!TPIF�-157 Men�u cannot� be disp�layed  (�TCP) ) O0���� d�9��K�]�o��, 
; �	 ����>TELEOP ~ǘLINE 0Ǒ�AUTO ABO�RTEDǘJOI�NT 100 %�����$���1���A��������ж�ȯҦ��ѰNG?TOL  @ʛ�A   ��Ѱ�PPINFO �� f�L�^�p����  ������ k���ۿſ�����5���Y�C�iϏ�%��� ү����������'߀9�K�]�o߁ߓߙ�P�PLICATIO�N ?t���|�Ha�ndlingTo�olǖ 
V9.40P/17�~��
8834ؒ���F0�	�549���������7DF�5�О�ǓNone���FRA�� �69��_ACoTIVE1�  ��� �  ��ސMO�D��������CH?GAPONL�����OUPL[�1	��� >�B�T�f����CUREQ 1]
��  Tp�p�ծ��������l��� ����������i3�l�p���^H��A�t
HTTHKY� FXv|�� *<N`���� ����//&/8/ J/\/�/�/�/�/�/�/ �/�/�/?"?4?F?X? �?|?�?�?�?�?�?�? �?OO0OBOTO�OxO �O�O�O�O�O�O�O_ _,_>_P_�_t_�_�_ �_�_�_�_�_oo(o :oLo�opo�o�o�o�o �o�o�o $6H �l~����� ��� �2�D���h� z�������ԏ��� 
��.�@���d�v���0��������TO������DO_CLEA�N���E�NM  �� p������ɯۯv�DSPDgRYRL���HI��o�@��G�Y�k�}��� ����ſ׿�������MAX��,�呿��=�X,�<�9�<���PLUGG,�-�9���PRC��Bm�"q�6�(ϗ�O���^�SEGF�K�� �� �m��G�Y�k�}�8������LAP$�7� �������+�=�O�a�s����� �T�OTAL_ƈ� �U�SENU$�1� �������RGDI_SPMMC�d��C�O�@@�1�O�"�D��-�_STRING 1��
�M��S���
��_ITE;M1��  n��� ������ $6H Zl~��������I/O SIGNAL���Tryout� Mode��I�npNSimul�ated��Ou�t`OVER�R!� = 100���In cyc�lT��Prog� Aborj��~JStatus���	Heartbe�at��MH F�aul��Aler�!/!/3/E/W/�i/{/�/�/�/  (���(����/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO�/WORИ�~A�/ XO�O�O�O�O�O __ $_6_H_Z_l_~_�_�_�_�_�_�_�^PO ���"`�KoEoWoio {o�o�o�o�o�o�o�o /ASew��bDEV%n�p9o ����#�5�G�Y� k�}�������ŏ׏������1�C�PALT�-j��OD����� ��ȟڟ����"�4� F�X�j�|�������į֯X�GRIB���� ���6�H�Z�l�~��� ����ƿؿ���� π2�D�V�h�z�����R �-��&���������� "�4�F�X�j�|ߎߠ� �������������PREGn�W���0� ~������������ � �2�D�V�h�z���������$�$AR�G_~@D ?	������  	$�$	[]��$:	��SBN_CONFIG�X�WqRCII�_SAVE  �$zm��TCEL�LSETUP �
%  OME�_IO$$%M�OV_H� ��R�EP��#��UTOoBACK� 	�tFRA:\�D� .D�z '�`�D�w� ��s  2�5/11/29 �20:26:16D�;D���#//h��C/j/|/�/�/�/�/D�X/�/?? (?:?L?�/p?�?�?�? �?�?�?g? OO$O6O HOZO�?~O�O�O�O�O��O�O���  c_�F_\ATBCK?CTL.TM�)_�;_M___q_8INI�m��j~CMESSAG� �Qz >�[ODE_D� ��j�XO�p�_@PwAUS6` !�� ,,		� ; :oHg.ohoRoto vo�o�o�o�o�o�o`@*<v��d~`TSK  mxw}_CUPDT�P�Wd�p�VXWZD_ENB�Tf
�v�STA�U�u��X�ISX UNT 2��vwy � 	 �������g1��i�0gK5h�D�R����D�z�������F� ��jc �D� �', Q� �Ir�������,�n/�MET��2@���y PQ�?�fU�??�?W�P�>�f�?U~�?�N�>ca�A=��=��<��d<z���>i5�SC�RDCFG 1vY ��� ����%�7�I�pD�Q�	ܟ�� ����ϯ��Z��~� ;�M�_�q�������6���FGR9��p�_Գ�PNA� 	�FѶ_ED�P1���� 
 �%=-PEDT-¿ �R�v���Es� -(FE�D�;9/��>���  ����2 �����B� ����{� ����j�����3��#�  �G�Y���G�ߠ�6�����4������Yހ���Z�l������5 K������Y�t���&�8���\���6��d ��Y�@����(��7�S0wY�@w��f���8�W��{�IZ��C/��2/���9{/��//LZݤ/?V/h/�/�/��CR���?�? Tn?�? ?2?�?V?԰~!�NO_DEL��ҲGE_UNUS�E޿дIGALL�OW 1� �  (*SY�STEM*
�	�$SERV_GR�[�@`REG�Eq$�C
��@NUM�J<�C�MPMU?@
��LAYK�
�PMPAL�P>UCYC10 N3^�P!^YSULSU`_�M5Ra�CLo_~�TBOXORI�E�CUR_�P�MPoMCNVV�P�10I^�PT4DL�I�p�_�I	*PR�OGRA�DP�G_MI!^Ko]`AQL+ejoTe]`B�o��N$FLUI_RESU9W�o�O�oF�dMR�N�@�<�? �;M_q��� ������%�7� I�[�m��������Ǐ ُ����!�3�E�W��2BLAL_OUT� �K���WD_ABOR:PcO���ITR_RTN � �$�빸�NO�NSTO�� �lHCCFS_UT�IL �̷C�C_AUXAXI�S 3$� h�}�j�|�����ƽCE?_RIA_I`@��נ��FCFG $�/�#���_LIM�B2�+� �� � M	��B\���$� �
Ԡ��)�Z�%%�/�����[������ ���!������L��(
5�����P}A�`GP 1H�����A�S�e�w�j6�CC� C7��UJ��]��p�����_�� C������U���������é�U̩�ձ�ߩ���������;���PC�k�����������*��������ɱ���������� D_� D!�!е!�!� ��&?��HE@ONFqIpC�G_P�P;1H� +EH� �ߟ߱����������C�KPAUS�Q1H�ף b�S� H�A��e������ ��������E�+�i� {�a���A?Iץ��MؐNFO 1���� ��3��$4�@k��?��@i*:��]/H��r���
=q�* �D�C�Ҭ��D
�1���@�G���Y�hPb�O� �� ��LLECT_��!�����EN�+`�ʒ���NDEַ#�/��1234567890�"�A��/ҵHw��#)j��< i{��;��/� �/`/+/=/O/�/s/ �/�/�/�/�/�/8?? ?'?�?K?]?o?�?�?@�?�?O�?��$�� ��IO #&��"S▒O��O�O�O`GTR�2'DM(��^�?�NN��(oM Z��_M[OR)q3)H��7� �U3��Y�_�_�_�_�_P�[bR�kQ*H�,S�I?<�<Ѡ<cz�KFd����P,�� ;ϒo�o�o˿�o�oœh�UY@E�oS� �sja.�PDB.���4�cpmidbg03��Рs:��>uq�pz��v  E��>x��}.���}�`��|�<�m!gP���t��~f��������@ud1:��?��XqDEF �-��zC)*�c�O�buf.txt�J��|K�[`�/DM��>���R�A���MCiR20_{RCdX���hS21�����G���CzA�d4�A�"R�A�A�=.�?��A�<� A%B���\B��GB�Ԗ�A���B�OB����D]^Dc���D���C@�j�D��Db�Ӱ���Ufg23DLQD�	>z�!� 2���}��yc
�@x�9� C�Ĵ  �D4G�E����  E%q�F�?� E�p�u��F�P E��f�F3H ���GM��Ъ5�>��33��?�xnt9�q@�Q5�����RpA?a��=L�/�<#�QU�@,��Cϒ���RSMO?FST +i���^��P_T1Ɠ4DM�A =ք�MOD�E 5dm�@��X	Q�M;��%���?���<��M>��Ͷ�TEKSTc�2i�`�R�Q6�O�K�CN�AB���n� 8��\�n�mCdB���Cp�p�����p:d�QS ��� �٨����4�I7>����>B8m5$�R�T_c�PROG %j%��d�1�h@�NUSER��x�K�EY_TBL  �e�����	
��� !"#�$%&'()*+�,-./(:;<=>?@ABCc��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������>�������������������������������������������������������������4A8�L�CK��F�y��ST�AT��2�X�_A�LM�����_AU_TO_DO�E�~FDR 3:i�2hi�US�x��i�$g��A� �����T *g�2� bf�� /�/9/;�*pm�P/ z/�~/h/�/�/�/�/ �/?"=�G?Y?k?/ |?�?L/�?�?�/�?�? OO�?*O@OvO�O6? �O�O�O~?�O	_�?*_ $_BOD_6_p_~_T_�_ �_�_�_�Oo)o;o�O Loqo_�o�o�_�o�o �o�o�o�oFXo ��No���o� ���@�N�$�b� x�����n����� �A��b�\�z�|�n� ������ʟ���(�֏ O�a�s������T�ʯ į��֯����2� H�~���>���ɿۿ�� �ϼ�2�,�J�L�>� xφ�\Ϛϰ����Ϧ� �1�C��T�y�$Ϛ� �߲ϴߦ�������� �N�`�߇���V� ����������� H�V�,�j�������v� ����$I��j d���v���� �0��Wi{& ��\����� /&/�:/P/�/�/F �/�/�/��/?�:? 4?R/T?F?�?�?d?�? �?�? O�/'O9OKO�/ \O�O,?�O�O�?�O�O �O�O�O
_ _V_h_O �_�_�_^O�_�_�O
o o"_$ooPo^o4oro �o�o�o~_�o	�_ ,Q�_rl�o�~ �����&�8��o _�q���.����dڏ ԏ��� �.��B� X�����N�ǟٟ럖� ��!�̏B�<�Z�\�N� ����l���������� /�A�S���d���4��� ��¯Ŀ�����Կ� (�^�p���ϩϻ�f� ���Ϝ���*�,�� X�f�<�zߐ����߆� ���#���4�Y��z� t�ߔ��������� ��.�@���g�y���6� ����l����������� (6J`��V� �����)��J DbdV��t� ��/�7/I/[/ l/�/<�/�/��/�/ �/?�/?0?f?x?&/ �?�?�?n/�?�?�/O O2?4O&O`OnODO�O �O�O�O�?__+_�? <_a_O�_|_�O�_�_ �_�_�_�_ o6oHo�O oo�o�o>_�o�ot_�o �oo�o0>R h��^o����o �1��oR�L�jl�^� ����|���Џ��� ?�Q�c��t���D��� ��ҏԟƟ ���"� 8�n���.�����˯v� ܯ���"��:�<�.� h�v�L�����ֿ迖� �!�3�ޯD�i���� �Ϣ��ϖ����ϴ��� �>�P���w߉ߛ�F� ����|�����
���� 8�F��Z�p���f� ��������9���Z� T�r�t�f��������� �� ��GYk� |�L������� �*@v�6 ���~�	/�*/ $/BD/6/p/~/T/�/ �/�/�/�?)?;?� L?q?/�?�?�/�?�? �?�?�?�?OFOXO? O�O�ON?�O�O�?�O �OO__@_N_$_b_ x_�_�_nO�_�_o�O oAo�Obo\oz_|ono �o�o�o�o�o(�_ Oaso��To� ��o�����2� H�~���>��ɏۏ� ���2�,�J�L�>� x���\���������� �1�C��T�y�$��� ����������į� �N�`��������V� ��ῌ������� H�V�,�jπ϶���v� ���߾�$�I���j� d߂τ�v߰߾ߔ��� ���0���W�i�{�&� ���\����������� �&���:�P�����F� ������������: 4R�TF��d� �� ��'9K�� \�,����� ���
/ /V/h/ �/�/�/^�/�/�
? ?"/$??P?^?4?r? �?�?�?~/�?	OO�/ ,OQO�/rOlO�?�O~O �O�O�O�O�O&_8_�? __q_�_.O�_�_dO�_ �_�O�_�_ o.ooBo�Xo�otc�$CR_�FDR_CFG �;re~�Q
UD1:�W:�TJ�d  �`�\��bHIST 3<�rf  �`  w?�R@tUAtBtC�PpUDtEtItgq�potw�_��bI�NDT_EN6p~�T�q��bT1_DO  1�U�u�sT2��w�VAR 2=�g�`qh_r C���R�d4���d�m[��RZ�`S�TOP��rTRL?_DELETNp�t� ��_SCRE�EN re�r_kcsc�rUw��MMENU 1>~��  <�\%�_��T��R��S /�U���e�w�ğ���� ��џ�	�B��+�x� O�a�����������ͯ ߯,���b�9�K�q� ������࿷�ɿ�� ��%�^�5�Gϔ�k�}� �ϡϳ��������H� �1�~�U�gߍ��ߝ� ��������2�	��A� z�Q�c������� ����.���d�;�M� ��q�������������YӃ_MANUA�L{��rZCD�a�?�y�rG ����R�f"
�"
?�|(��PK�WGR�P 2@�yaqB1� � s��� ��$DBCO�pR�IG���v�G_E�RRLOG A���Q�I[m ��NUMLIM��s��u
�PXWORK 1B�8���//�}�DBTB_�� !C%�ap�S"� ��aDB_AWAYz��QGCP �r�=�ןm"_AL(�F�_�Yz���p�p�vk  1D� , 
��/"�/%?/(_M�pqw,�@�=5ONTIM6����t�_6�)�
�0�'MOTN�ENFpF�;REC�ORD 2J�� �-?�SG�O� �1�?"x"!O3OEOWO �8_O�O�?�OO�O�O �O�O�O(_�OL_�Op_ �_�_�_A_�_9_�_]_ o$o6oHo�_lo�_�o �_�o�o�o�oYo}o 2�oVhz��o� �C�
��.�� R��K��������Џ ?��ߏ�*�����+� b�t�㏘�����Ο=� O�����:�%���p� ߟ񟦯��O�ǯ�]� �����H�Z����� ����#�5����ϩ��i"TOLEREN�Cv$Bȿ"� L���� CSS_CC�SCB 2K�\0"?"{ϰϟ� ��7��
����@�R� d�3߈ߚ�"�x��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy���� �������R�LL]�La��m1T#2 C��C��F�^ +A�C�pC���#�0�� 	 A����B���?�  �$�����\0袰�0��B� �`#s�K/]/o/�ϓ/�/�/s/�/�/���ʈ�̍5�οRr���o;�&;Ȧ�/��/`?;
�@��O?�?�?�?�Ȏ0AF��?{F�A OO�7�1���9M	AB
AZOdBAE�9�$O�O�O�Oi:P��`^�@0�DJCA�� @��
qX-.
[#_   M?�>O�ڴ�q_�_�_�_:W�A<o:[@<ǲ/o�/�_+o`Poboto�eACHC�jV�WB$�Dz�cD�`�a=/�o�oo�oHW�a.+!��2=t�,yD��YqC��I?�-t�s� js�w�yj���� ���Q���@`� �$�����A����B މ�o��'�9��_]� o�N���r���ɟ۟_��B�ʄ��YZ>`���@'BO�B�e�@�Vz�?RW�:C�l�R�0d�v����� `_ м¯���
���̯9� ,�]�o��� �H����� ٿ뿊��ƿ3�E�W� iϬ���$ϱ����� � �����/�A�S߶�w� V�h߭ߌ��S���ߐ�_�f	��H�?� Q�~�u������� �����D��-�g� q�������������
 @7Icm�8�߾�  ��� ��)M@qd v������� //I/P�m/�v/�/ �/�/�/�/�/�/?3? *?<?i?`?r?�?^/�? �?�?�?�?O/O&O8O JO\O�O�O�O�O�O�O|�O�g	  Q��P�s ��PC4p*p�pp6U6P\C9p/p�� ]V^PM]�6P�:P�>P�VJ_+�^P�bP�fP�VLr]v��Tp Q
k� ��_oo�id1Q&oNo ;o_co�oˏUUA   �o�k1Q@�  �o�k�b�]����Up( �� 1��6�1C���C�cPfL��?#��c>�{��2�`�cP�@@�d�,�r�`B�cP>�s�q;C��p����b�t�<�o?�PH?�)S�B�tq0�q�p�r�`B���eDIC�&�Q�4( �o�z�UU�5�=���Bd�=�^�R?T�:C�HQ�-R��?����C����B�F��b��`ځ`  �?�p���U�[?����}t��$���$�DCSS_CLL�B2 2M���p�P�^?�NS�TCY 2N����   �������ʟ؟��� � �2�D�Z�h�z��������¯ԯ��SA�D�EVICE 2O��!�$��4&V� h�������˿¿Կ� ��
�7�.�[�R�ϑ���ϵ�����4(A�HN?DGD P��*��Cz�A�LS 2Q��_�Q�c�u߇���߽߫���?�PARAM RP��1��`�&�RBT 2T��� 8�P<C�'p �qi�l��s@"�R��(qI�ʹX��0�pB CW  ��B\x�N��`�Z����%��)� ��X�j��p����zq��I���B �(s,�F� �p�V��q���b��B ��4&c �S�e� l�4+����H1~ޡ���D�C��$Z��b���A�,� 4�u@�X�@��^@w����]B���B��cP%��C4��C3:^C4��nЬ ��p8�-�B{B���A���� l���C�C3��JC4jC3���yn+�3 Dff 2�A PB W4+@:�]o�W �����/�/ P/'/9/K/]/o/�/�/ �/�/?�/�/�/?#? 5?�?Y?k?�?�?�o�? �?O�?6O!OZOlOWO �O�Es�?�?�?�O�O _�O�OL_#_5_G_Y_ k_}_�_�_�_ o�_�_ �_oo1o~oUogo�o �o�o�o�owO D /Aze����O �o�o
��o��R�)� ;���_�q��������� �ݏ�<��%�r�I� [�m��������ǟٟ &�8��\�G���k��� ����گů����� F��/�A�S�e�w�Ŀ ������ѿ����� +�x�O�aϮυϗϩ� ������,���b�t� ﯘ߃߼ߧ������ ���:��C�U߂�Y� k����������� 6���l�C�U�g�y� ���������� ��	 -?Q���� ���@+d vQ������ ��*///%/r/I/ [/�//�/�/�/�/�/ &?�/?\?3?E?�?i? {?�?�?U�?�?"O4O OXOCO|OgO�O{� �?�O�?�O�O0___ f_=_O_a_s_�_�_�_ �_�_o�_oo'o9o Ko�ooo�o�o�o�o�o �O:%^I�������H�$D�CSS_SLAV�E U����	���z_�4D  	��A�R_MENU V	� �j�|�������ď�BY�� ��~�?�SHOW 2W>	� � �b�a G�Q�X�v��������� П֏���� @�:� d�a�s���������� ߯��*�$�N�K�]� o�������̯ɿۿ� ��8�5�G�Y�k�}� �϶�����������"� �1�C�U�g�yߠϝ� ���������	��-� ?�Q�c��s����� ��������)�;�M� t�������������� ��%7Ip�m ���������� !3ZWi�� �J����// DA/S/e/��/��/ �/�/�/�/?./+?=? O?v/p?�/�?�?�?�? �?�??O'O9O`?ZO �?�O�O�O�O�O�OO �O_#_JOD_nOk_}_ �_�_�_�_�O�_�_o 4_.oX_Uogoyo�o�o �o�_�o�o�ooBo ?Qcu���o:����CFG MX)�3�3q5p��FRA:\�!�L+�%04d.WCSV|	p}�� �qA g�CHo�zv�	����3q�����́܏� �|��4��JP�����qp1� �R�C_OUT Y���C��_�C_FSI ?~i� .� ������͟����� >�9�K�]��������� ίɯۯ���#�5� ^�Y�k�}�������ſ �����6�1�C�U� ~�yϋϝ��������� �	��-�V�Q�c�u� �ߙ߽߫�������� .�)�;�M�v�q��� ����������%� N�I�[�m��������� ��������&!3E ni{����� ��FASe �������� //+/=/f/a/s/�/ �/�/�/�/�/�/?? >?9?K?]?�?�?�?�? �?�?�?�?OO#O5O ^OYOkO}O�O�O�O�O �O�O�O_6_1_C_U_ ~_y_�_�_�_�_�_�_ o	oo-oVoQocouo �o�o�o�o�o�o�o .);Mvq�� �������%� N�I�[�m��������� ޏُ���&�!�3�E� n�i�{�������ß՟ ������F�A�S�e� ��������֯ѯ��� ��+�=�f�a�s��� ������Ϳ����� >�9�K�]φρϓϥ� ����������#�5� ^�Y�k�}ߦߡ߳��� �������6�1�C�U� ~�y����������� �	��-�V�Q�c�u� �������������� .);Mvq�� ����% NI[m���� ����&/!/3/E/ n/i/{/�/�/�/�/�/��/�/3�$DCS�_C_FSO ?����71 P ? ?T?}?x?�?�?�?�? �?�?OOO,OUOPO bOtO�O�O�O�O�O�O �O_-_(_:_L_u_p_ �_�_�_�_�_�_o o o$oMoHoZolo�o�o �o�o�o�o�o�o%  2Dmhz��� ����
��E�@� R�d���������ՏЏ ����*�<�e�`� r���������̟��� ��=�8�J�\�����|��?C_RPI4>F?�������3?��&�o����� >SLү@d������%� 7�`�[�m�Ϩϣϵ� ���������8�3�E� W߀�{ߍߟ������� �����/�X�S�e� w����������� �0�+�=�O�x�s��� ���������� 'PK]o��� �����(#5 Gpk}����� Q���/6/1/C/U/ ~/y/�/�/�/�/�/�/ ?	??-?V?Q?c?u? �?�?�?�?�?�?�?O .O)O;OMOvOqO�O�O �O�O�O�O___%_ N_I_[_m_�_�_�_�_ �_�_�_�_&o!o3oEo noio{o�o�o�o�o�o �o�oFASe�������>�N�OCODE Z�U��?�P�RE_CHK �\U��pA �p?�< ��pU�x]�o�U� 	 <Q� �������ۏ�Ǐ� #����Y�k�E����� {�şן��ß���� C�U�/�y�����s��� ӯm���	���?�� +�u���a�������ɿ �Ϳ߿)�;��_�q� K�}ϧϝ������ω� ��%����[�m�Gߑ� ��}߯��߳����!� ��E�W�1�c��g�y� ������������A� S�-�w���c������� ������+=a sM_����� �'�]o	 ������/ #/�G/Y/3/e/�/i/ {/�/�/�/�/?�/? C?9Ky?�?%?�?�? �?�?�?	O�?-O?OO KOuOOOaO�O�O�O�O �O�O�O)_____q_ K_�_�_a?�_�_�_�_ o%o�_Io[o5oGo�o �o}o�o�o�o�o�o �oEW1{�g� ��_����/�A� �M�w�Q�c������� ���Ϗ�+���a� s�M���������ߟ� ��'���3�]�7�I� �����ɯۯ���� ���G�Y�3�}���i� ��ſ��������1� C���+�yϋ�eϯ��� ����������-�?�� c�u�Oߙ߫߅ߗ��� �����)��M�_�U� G���A�������� �����I�[�5���� k������������� 3EQ{q�� �]����/A ewQ���� ���/+//7/a/ ;/M/�/�/�/�/�/� �/?'??K?]?7?�? �?m??�?�?�?�?O �?5OGO!O3O}O�OiO �O�O�O�O�O�/�O1_ C_�Og_y_S_�_�_�_ �_�_�_�_o-oo9o co=oOo�o�o�o�o�o �o�o__M_�o k�o����� ���I�#�5���� k���Ǐ��ӏ��׏� 3�E��i�{�5c��� ß�����ӟ�/�	� �e�w�Q�������ѯ 㯽�ϯ�+��O�a� ;��������Ϳ߿y� ���!�K�%�7ρ� ��mϷ��ϣ������� ��5�G�!�k�}�W߉� �ߩ������ߕ��1� ��g�y�S���� ��������-��Q� c�=�o���s������� ������M_9 ��o���� �7I#mY k������!/ 3/)/i/{//�/�/ �/�/�/�/�/?/?	? S?e???q?�?u?�?�? �?�?OO�?%OOOE/ W/�O�O1O�O�O�O�O __�O9_K_%_W_�_ [_m_�_�_�_�_�_�_ o5oo!oko}oWo�o �omO�o�o�o�o1 UgAS��� ���	����Q� c�=�����s���Ϗ�o ������;�M�'�Y� ��]�o���˟���� ۟�7��#�m��Y� �����������!� 3�ͯ?�i�C�U����� ��տ�������	� S�e�?ωϛ�uϧ����Ͻ������$�DCS_SGN �]	�E��-����29-N�OV-25 20�:38 ��N�27�_�x�x� [}�t��q�т�x���ك�JѨ�EƼÞ� ��ǖ��  1�HOW �^	� �x�/�VERSI�ON =��V4.5.2��E�FLOGIC 1�_���  	������C��R�%�P�ROG_ENB � ��:�{�s�U?LSE  X���%�_ACCLI�M�����d���WRSTJNT��E��-�EMO�|�zя�$���INIOT `2�����OPT_SL ?�		�	�
 	�R575��]�74jb�6c�7c�50���1���C���@�TO  L��� �]V�DEX��dE��x�PATH ;A=�A\k�}��HCP_CL?NTID ?�:� D�ռ���IAG_GRP �2e	�����z�	 @� � 
ff?aG���B�  �2��/�8[I@�c�ς!�7@��z�@^�@�
�!��mp�2m15 8901234567�����  ?���?�=q?���
?޸R?��Q�?��?������(�?Ǵz���x�@�7  A_�Ap !�7A�88_�B4�� ��L�x��
�@�@���\@~�R@x�Q�@q�@j��H@c�
@\���@U�@Mp��//'$�; |�O)H��@Ct }>d 9��@4�_/\)@)� #t {@��/��/�/�/�/P'?�̗�?���_ ?�}p�?u?on{?s ?\�Q�? ?2?D?V?�h8�
=?����0w5�z�H?�p�h��?^�R�?�?�?�?�?h8�U�t0���@�?��0�;@&O 8OJO\OnOP'�$_� _Y_k_�O?_�_�_�_ �_�_s_�_�_1oCo!o goyoo�o��Bj"� ��2{1�@"?����f�t0�d"5!=�
u4V��u"��B3t�A>u��?@�[q��@`,=q��=b��=�E�1>�J�>�n��>��H"<�;o �z�s�q���� �x�C�@<(��Uz� 4��� ����A@x�? *�o��m*�P�b�� �tn���2���Ώ�����i>J��&��bN2�"��G��N��o@�@v���0����@ffr!�l ��33���({��"C�� ƒ�I�CH�)C.dBت"8"����'���"~��A?�&"K����pf�B��@�p�������p���?}Wͽ�r�������@�~Ᵹ-M���Cu=TG���}�)D��C�Ҭ�D�xО������3���N�T������1��@�G���Y�@Rs"� ���ǿ���ֿ�����<O3[>���P�_�Ǿ��J���#�!�o���CT_CONF_IG f��>|�egY���STBF_TTS��
����О�}���1�MAU�����ҿMSW_CF��g��  # ��OCV7IEW��h!�-���s߅ߗߩ߻� �ߟ�a�����,�>� P���t������� ]�����(�:�L�^� �������������k�  $6HZ��~ ������y  2DVh���`����v�RC�	i���!�0./S/�B/w/f/�/�/�/��S�BL_FAULT� j*6��!GP�MSK���'��TD?IAG k��-�������U�D1: 6789?012345I2��=1���%P\υ?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�Od696ħI�r
t?�O|�TR'ECP"?4:
B44_ [7M[s?p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�O�O�O�o�7�UMP_OPT�IO=��.�aTR�����)uPME���Y_TEMP�  È�3B�C�gp�B�QtUN�I����gq�YN_?BRK lL�7�?EDITOR�a�a�@�r_
PENT �1m)  ,�&TPSNAP�^P ��l&MTP�G�p��TEL3EO+�f�&�/�����z�����ۏ ����5��Y�k�R� ��v���ş���П� ���C�*�g�N�v��� ���������ޯ���?�Q���EMGDI_STAzuV�gq��uNC_INFO� 1n!��b����X���������n�1o!� ��o���
�
�d�oU�g�y� �ϝϯ���������	� �-�?�Q�c�u߇ߙ� �߽��� u����
�� *�B�*�P�b�t��� �����������(� :�L�^�p��������� 2�������9�C Ugy����� ��	-?Qc u�������� //1;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?��?�?�?O)/O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�?�?�_ �_o�_3O=oOoaoso �o�o�o�o�o�o�o '9K]o�� ��_�_����+o 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y��������ӟ ���	�#�-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� �7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߹��� �������%�/�A�S� e�w��������� ����+�=�O�a�s� �������������� �'9K]o�� ������# 5GYk}�	�� ����/1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?��?�?�?�? /O)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�? �_�_�_�_O�_!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew��_�_��� �o�+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o���� ���ɟ۟���#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� ���߹���������� %�7�I�[�m���� �����������!�3� E�W�i�{��߇����� �����/AS ew������ �+=Oas ����������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?���?�? �?�?��?OO1OCO UOgOyO�O�O�O�O�O �O�O	__-_?_Q_c_ u_�?�_�_�_�_�?�_ oo)o;oMo_oqo�o �o�o�o�o�o�o %7I[m�_u� ���_���!�3� E�W�i�{�������Ï Տ�����/�A�S� e��������u�� ����+�=�O�a�s� ��������ͯ߯�� �'�9�K�]�w����� ����ɿ�����#� 5�G�Y�k�}Ϗϡϳ� ����������1�C� U�g߁��ߝ߯���ۿ ����	��-�?�Q�c� u����������� ��)�;�M�_�y߃� ������������ %7I[m�� �����!3 EWq�c����� ����////A/S/ e/w/�/�/�/�/�/�/ �/??+?=?O?i{ �?�?�?�?��?�?O O'O9OKO]OoO�O�O �O�O�O�O�O�O_#_ 5_G_�?s?}_�_�_�_ �?�_�_�_oo1oCo Uogoyo�o�o�o�o�o �o�o	-?Qk_ u����_��� ��)�;�M�_�q��� ������ˏݏ��� %�7�I�cQ������ ���ٟ����!�3� E�W�i�{�������ï կ�����/�A�[�� �$ENETM�ODE 1p����  
k�k�f�����j��OATCFG �q�����Ѵ��C���DAT�A 1rw�Ӱ�.��*	�*��'�9�K�]�l�dlύ�e��ϻ�������� �'ߡϳ�]�o߁ߓ� �߷�1���U����#� 5�G�Y����ߏ��� ��������u��1�C� U�g�y������)��� ����	-����c�u�����j�RPOST_LO��	t�[
׶#5�Gi�RROR_P-R� %w�%L��XTABLE  w�ȟ�����RSEV_NUM� ��  ����  �_AUT�O_ENB  ����X_NO5! �uw���" W *�x �x �x 	�x + +w �/�/�/�Q$FLTR=/O&H�IS#]�J+_A�LM 1vw� e�[x,e�+�/�Q?c?u?�?�?�?�/_\"W   w�v!����:j�TCP_V_ER !w�!x޻?$EXT� _R�EQ�&�H)BCSsIZKO=DSTKhI�f%�?BTOL�  ]Dz�"��A =D_BWD��0�@�&�A���CDI�A wķ���]�KSTEP�O�Oj�>POP_DO�Oh��FDR_GRP s1xw��!d 	�?x�_��yPs�Y�Q�'�M"����l��T� ����VyS�_�]��TB CA��߅Az�m]A^���_`���@՚��_�[Go2oWo�}oho�o�o�o�]@\��G?�"�?k��)>���n
 F@c�`�bX.��o(2�o�oZ�E~i|A@`�t@'S33�uh}@�q� g��yPq��|yP�G�  @�Fg��fC�8RL��}?�  h��6�X�����875t���5���5`+���~X���>�� �y���_�|:� ��͓FEATUROE y���@���Handl�ingTool ��]Engl�ish Dict�ionary�4�D St��ard���Analog� I/O>�G�gle ShiftZ��uto Soft�ware Upd�ate�mati�c Backup����ground� Edit ��C_ameraU�FY��CnrRndIm����ommon �calib UI���nˑ�Monoitor$�tr�?Reliabn���DHCP �[�at�a Acquis�3�\�iagnos���R�v�ispla�yΑLicens�Z�`�ocument Viewe?��^�ual Che�ck Safet�y��hance�d���s�Fr�ܐ�xt. DI�O /�fi��@�e�nd�Err>�L(��\�4�s[�rP�K�� �@
�FCTN /Menu��vZ����TP In��faycĵ�GigE־��Đp Mask� Exc�g=�H�T԰Proxy �Sv��igh-wSpe�Ski��� Ť�O�mmuni�c��onsV�ur໰��q�V�ײcon�nect 2��n{crְstru!�$�ʴ�eۡ��J��X��KAREL Cmod. L�ua�~��Run-Ti<��Env�Ȟ�el u+��s��S/W��ƥ���r�Book�(System)�
�MACROs,~M�/Offseu��p�HO���o�u�MR�8�4���MechStop+�t����p�im�q���x�R������odo�witc�h�ӟ�.��4�O�ptmF��,�fi�l䬳�g��p�ul�ti-T�Γ�P?CM fun�Ǽ��o��������Regeie�rq���riݠ�F���S�Num �Sel��/�:� Adjua�*�W�q�h�tatu��ߪ��RDM Robo}t�scove'���ea��<�Fre�q Anlyq�Rem��O�n5�����ServoO�!��?SNPX b-�v�;SN԰Cliܡ?r�Libr&�_��Q ��q +oJ�t���ssag��X�@ 0����	�@/Iս��MILIB��P� Firm���Pλ�AccŐ͛TPsTXk��eln���������orq}uo�imula=�4�|u(�Pa&���ĐX�B�&+�ev.̸��ri��TU�SB port ��iPf�aݠ&R� EVNT� n?except�����%5��VC�rl�c���V���"�%4q�+SR SCN�/gSGE�/�%UI	�?Web Pl��>���A43��ۡ��ZDT Applj�<
�{1EOAT�����&0?�7Gridp�񾡬=�?iR�"�.5� F���/גRX-10iA/L�?�Alarm Caouse/��ed(��All Smoo�th5���C�sciyi+�V�Load�ΌJUpl�@w�to�S ��rityA_voidM(�s7�1t�@�ycn��0���_�CS+���g. c��XJo� ��-T3_H�.RX��U����Xcollabo����RA�:�.9�D��in���N�RTHI
�On��e Hel����ֿ������1trU�ROS Eth$��A� �����;,�G �B�,|HUpV�%�W�3t ԰�_iRS�ݐ��64MB DRsAM�o�cFRO8���L8F FlD���d��2M �A:�opm�bԕex@V�
�sh�qD��wce�u��p��|tyn�sA�
�%�Ar����J��^�.v� P)Q/sbS�`���8O�N��mai��U����R�q�T1��^FC+Ԍ%̋Fs�9�ˌk̋��Typ߽FC%�hױV�N Sp�ForްK��Ԇ��lu!����cp�P'G j�֡�RJ�[L`Sup"}���֐f��crFP��lu� ��al�����r��i�
q�4@�ް�uest,IMPLE ׀6*|H�Z���c0�BTeap(�|���$rtu���V�9HMI�¤��wUIFc�pono2D�BC�:�L�y�p� ��������ʿܿ	� � �?�6�H�u�l�~ϫ� �ϴ���������;� 2�D�q�h�zߧߞ߰� �������
�7�.�@� m�d�v������� �����3�*�<�i�`� r��������������� /&8e\n� �������+ "4aXj��� �����'//0/ ]/T/f/�/�/�/�/�/ �/�/�/#??,?Y?P? b?�?�?�?�?�?�?�? �?OO(OUOLO^O�O �O�O�O�O�O�O�O_ _$_Q_H_Z_�_~_�_ �_�_�_�_�_oo o MoDoVo�ozo�o�o�o �o�o�o
I@ Rv����� ����E�<�N�{� r�������Տ̏ޏ� ��A�8�J�w�n��� ����џȟڟ���� =�4�F�s�j�|����� ͯį֯����9�0� B�o�f�x�����ɿ�� ҿ�����5�,�>�k� b�tφϘ��ϼ����� ���1�(�:�g�^�p� �ߔ��߸������� � -�$�6�c�Z�l�~�� �����������)� � 2�_�V�h�z������� ��������%.[ Rdv����� ��!*WN` r������� //&/S/J/\/n/�/ �/�/�/�/�/�/?? "?O?F?X?j?|?�?�? �?�?�?�?OOOKO BOTOfOxO�O�O�O�O �O�O___G_>_P_ b_t_�_�_�_�_�_�_ oooCo:oLo^opo �o�o�o�o�o�o	  ?6HZl�� �������;� 2�D�V�h�������ˏ ԏ���
�7�.�@� R�d�������ǟ��П �����3�*�<�N�`� ������ï��̯��� �/�&�8�J�\����� ������ȿ�����+� "�4�F�Xυ�|ώϻ� ����������'��0� B�T߁�xߊ߷߮��� ������#��,�>�P� }�t��������� ����(�:�L�y�p� �������������� $6Hul~�����  ?H552���21R785�0J614AwTUP'545'�6VCAMC�RIbUIF'2�8cNRE52�VR63SCH�LIC�DOC�V�CSU86�9'02EIOC��4R69VEgSET?UJ7U�R68MASK^PRXY{7OCO#(3?+ �&3j&J6%53��H�(LCHR&O�PLG?0�&MH�CRS&S�'MCS�>0.'552MD�SW+7u'OPu'M�PRv&��(0&PCMzR0q7+ 2l� �'51J51�8�0JPRS"'69�j&FRDbFRE�QMCN93�&SNBA��'SHLBFM1G�8�2&HTC>TMsIL�TPA�oTPTXcFELF�� �8J9�5�TUTv'95�j&UEV"&UEC�R&UFRbVCC�
XO�&VIPnFC;SC�FCSG���IWEB>HTT>R6��H;RV�CGiWIGQWIP�GS�VRCnFDGvu'H7�7R66J�5'R�8R51*
(6�(2�(5V�)J8�86�L=I%� �84g662R�64NVD"&R�6�'R84�g79ڎ(4�S5i'J7�6j&D0�gF xR�TSFCR�gCR�Xv&CLIZ8IC�MS�Sp>STY:nG6)7CTO>���7�NNj&ORqS�&C &FCB��FCF�7CH>F�CR"&FCI�VF�C�'J�PO7GBfMv�8OLaxENDS&�LU�&CPR�7L�WS�xC�STxT�E�gS60FVmR�IN�7IHaF �я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� !3EWi{� ������ /ASew��� ����//+/=/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]? o?�?�?�?�?�?�?�? �?O#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �_�_�_�_�_	oo-o ?oQocouo�o�o�o�o �o�o�o);M _q������ ���%�7�I�[�m���������Ǐُ��  H55�2��21�R7�8�50�J61�4�ATUP7�5�457�6�VCA�M�CRI��UI�F7�28��NREv�52v�R63�wSCH�LICƚ�DOCV�CSU��8697�0F�E�IOCǛ4�R6=9v�ESETW�u��J7u�R68�M�ASK�PRXY���7�OCO��3�W����6�3�J6�5�536�H$�LC�HƪOPLGW�0^�MHCRǪS���MCSV�0��55�F�MDSW���OP��MPR���6��06�PCM��R0`E˓�F���6�51f��51��0f�PRSv��69�FRD���FREQ�MCN��936�SNBA�כ%�SHLB�M�E��ּ26�HTC�V�TMIL�6�T{PAV�TPTX��#ELړ�6�8%�#���J95��TUTv��95�UEV��wUECƪUFR���VCCf�O��VI�P��CSC��CS�Gƚ$�I�WEBnV�HTTV�R6՜���S���CG��IG���IPGS'�RC���DG��H7��RK66f�5�u�R��WR51f�6�2�I5v�#�J׼��6���LU�5�s�v�4��6�6F�R64�NV�D��R6��R84֦79�4��S5n�J76�D0u�FRTS&�CR�CRX��CLI&�e�CMSV�sV��STY��6�CT�OV�#�V�75�NN��ORS����6�F�CBV�FCF��C�HV�FCR��FC-IF�FC��J#�˵G
M��OL�E�NDǪLU��CPUR��Lu�S�C$��StTE�S60n�FVRV�IN��IH���m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s�@��������͏ߏ��STD�LANG���0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰����RBT
�OPTN������'�9�K� ]�o�����������DPN	���)� ;�M�_�q��������� ������%7I [m����� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	-?Qcu� �������� )�;�M�_�q������� ��ˏݏ���%�7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w� ��������ѿ���� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� ������1�C�U�g� y���������������@	-?Qc�f�������9�9��$FEAT�_ADD ?	����  	�#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������DEMO y?   �L� B�T߁�xߊ߷߮��� ��������G�>�P� }�t��������� ����C�:�L�y�p� �������������� ?6Hul~� �����; 2Dqhz��� ��� /
/7/./@/ m/d/v/�/�/�/�/�/ �/�/?3?*?<?i?`? r?�?�?�?�?�?�?�? O/O&O8OeO\OnO�O �O�O�O�O�O�O�O+_ "_4_a_X_j_�_�_�_ �_�_�_�_�_'oo0o ]oTofo�o�o�o�o�o �o�o�o#,YP b������� ���(�U�L�^��� ��������ʏ��� �$�Q�H�Z���~��� ����Ɵ����� � M�D�V���z������� ¯ܯ��
��I�@� R��v���������ؿ ����E�<�N�{� rτϱϨϺ������ ��A�8�J�w�n߀� �ߤ߶��������� =�4�F�s�j�|��� ����������9�0� B�o�f�x��������� ������5,>k bt������ �1(:g^p ������� / -/$/6/c/Z/l/�/�/ �/�/�/�/�/�/)? ? 2?_?V?h?�?�?�?�? �?�?�?�?%OO.O[O ROdO�O�O�O�O�O�O �O�O!__*_W_N_`_ �_�_�_�_�_�_�_�_ oo&oSoJo\o�o�o �o�o�o�o�o�o "OFX�|�� �������K� B�T���x�������ۏ ҏ����G�>�P� }�t�������ןΟ�� ���C�:�L�y�p� ������ӯʯܯ	� � �?�6�H�u�l�~��� ��Ͽƿؿ����;� 2�D�q�h�zϔϞ��� �������
�7�.�@� m�d�vߐߚ��߾��� �����3�*�<�i�`� r������������ �/�&�8�e�\�n��� ��������������+ "4aXj��� �����'0 ]Tf����� ���#//,/Y/P/ b/|/�/�/�/�/�/�/ �/??(?U?L?^?x? �?�?�?�?�?�?�?O O$OQOHOZOtO~O�O �O�O�O�O�O__ _ M_D_V_p_z_�_�_�_ �_�_�_o
ooIo@o Rolovo�o�o�o�o�o �oE<Nh r������� ��A�8�J�d�n��� ����яȏڏ���� =�4�F�`�j������� ͟ğ֟����9�0� B�\�f�������ɯ�� ү�����5�,�>�X� b�������ſ��ο�� ��1�(�:�T�^ϋ� �ϔ��ϸ������� � -�$�6�P�Z߇�~ߐ� �ߴ���������)� � 2�L�V��z���� ��������%��.�H� R��v����������� ����!*DN{ r������� &@Jwn� ������// "/</F/s/j/|/�/�/ �/�/�/�/???8? B?o?f?x?�?�?�?�? �?�?OOO4O>OkO bOtO�O�O�O�O�O�O�__0]   'XF_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o o&o8oJo\ono�o�o �o�o�o�o�o�o" 4FXj|��� ������0�B� T�f�x���������ҏ �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ����������
��.�  /�)�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?V?h?z?�?�? �?�?�?�?�?
OO.O @OROdOvO�O�O�O�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|� �������� 0�B�T�f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�\�n� ���������������� "4FXj|� ������ 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<N `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������P ��$�4�8�+� N�`�r߄ߖߨߺ��� ������&�8�J�\� n����������� ���"�4�F�X�j�|� �������������� 0BTfx�� �����, >Pbt���� ���//(/:/L/ ^/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?l? ~?�?�?�?�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�o&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�`�r����������� ����&8J\ n������� �"4FXj| �������/ /0/B/T/f/x/�/�/ �/�/�/�/�/??,? >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO ^OpO�O�O�O�O�O�O��O __$_6Y�$F�EAT_DEMO�IN  ;T��fP�<PNTIND�EX[[jQ�NPI�LECOMP �z����Q�iRIU�PSETU�P2 {�U~�R�  N �Q��S_AP2BCK� 1|�Y  #�)7Xok%�_8o<P�P&oco9U�_�o o�oBo�o�oxo�o 1C�og�o��, �P�����?� �L�u����(���Ϗ ^�󏂏�)���M�܏ q������6�˟Z�؟ ���%���I�[��� �����D�ٯh���� ��3�¯W��d���� ��@�տ�v�Ϛ�/� A�пe����ϛ�*Ͽ� N���r���ߨ�=��� a�s�ߗ�&߻���\� �߀��'��K���o� ��|��4���X����� ��#���G�Y���}�� ����B���f������1�Y�PP�_ 2>�P*.VR8���*��������l PC���OFR6:�2�V�TzPz�w�]PG���*.Fo/��	�:,q�^/�STMi/ �/ /�-M/�/�H�/?�'?�/�/g?�GIFq?�?�%��?D?V?�?�JPG �?O�%O�?�?oO�
#JSyO�O��5C�O�MO%
JavaS�cript�O�?C�S�O&_�&_�O %�Cascadi�ng Style SheetsR_���
ARGNAMOE.DT�_��� �\�_S_�A�T�_�_>�PDISP*�_���To�_�QLaZoo�CLLB.ZIXwo2o$ :\�a\�o��i�AColla�bo�o�o
TPEINS.XMLƱ_:\![o�QCu�stom Too�lbarbiPA?SSWORDQo��?FRS:\�d�B`Passwor�d Config ���/��(�e��� �����N��r��� ��=�̏a������&� ��J���񟀟���9� K�ڟo�������4�ɯ X��|���#���G�֯ @�}����0�ſ׿f� �����1���U��y� �ϯ�>���b���	� ��-߼�Q�c��χ�� �߽�L���p��ߦ� ;���_���X��$�� H�����~����7�I� ��m���� �2���V� ��z���!��E��i {
�.��d� ���S�w p�<�`�/� +/�O/a/��//�/ 8/J/�/n/?�/�/9? �/]?�/�?�?"?�?F? �?�?|?O�?5O�?�? kO�?�OO�O�OTO�O xO__�OC_�Og_y_ _�_,_�_P_b_�_�_ o�_oQo�_uoo�o �o:o�o^o�o�o) �oM�o�o��6 ��l��%�7�� [����� ���D�ُ h�z����3�,�i� �������ßR��v�������$FIL�E_DGBCK �1|������ < ��)
SUMMA�RY.DG!�͜�MD:U���ِ�Diag Sum�mary����
C?ONSLOG��n����ٯ���Con�sole log����	TPACC�N�t�%\������TP Accou�ntin;���F�R6:IPKDM�P.ZIPͿј
��ϥ���Exception"�ӻ���MEMCHECKЏ�������-�Me�mory Dat�a����&n )��RIPE�~ϐ��%ߴ�%�� Packet L:����L�$�c���S�TAT��߭�� %A�Sta�tus��^�	FTAP����	��/��mment TB�D2�^� >I)ETHERNEw��
�d�u�﨡Et�hernJ�1�fi�guraAϩ��DCSVRF&����7����� verify all:���� 4��DIFF/��'���;�Q�diff��r�d���CHG01������`A����it�2���270���fx�3���I ��p�VTR�NDIAG.LS�u&8���� �Ope��L� ��n�ostic��T�)VDEV�DAT�������Vis�Dev�ice�+IMG@��,/>/�/:�i$�Imagu/+U�P ES/�/FORS:\?Z=���Updates OListZ?��� �FLEXEVEN���/�/�?���1 ?UIF EvM�M����-vZ)CRSENSPK�/�˞�\!O���C�R_TAOR_PE�AKbOͩPSRB?WLD.CM�O͜�E2�O\?.�PS_ROBOWELS���:GIG��@_�?|d_��GigE�(�O��N�@�)>UQHADOW__D_�V_�_��Shad�ow Chang�e����dt�RRCMERR�_�_�_�oo��4`CFG �Erroro ta�ilo MA��k�CMSGLIB goNo`o�o|R�e��z0�ic�o�a�)�`ZD0_O�os��7ZD�Pad�l{ �RNOTI��Rd���Not�ific����,�AG��P�ӟt��� ������Ώ]����� (���L�^�폂���� ��G�ܟk� ����6� şZ��~������C� د�y����2�D�ӯ h��������¿Q�� u�
�ϫ�@�Ͽd�v� Ϛ�)Ͼ���_��σ� ߧ�%�N���r�ߖ� ��7���[�����&� ��J�\��߀���3� ����i����"�4��� X���|������A��� ��w���0��=f �����O�s �>�bt �'�K���/ �:/L/�p/��/�/ 5/�/Y/�/ ?�/$?�/ H?�/U?~??�?1?�? �?g?�?�? O2O�?VO �?zO�OO�O?O�OcO �O
_�O._�OR_d_�O �__�_�_M_�_q_o o�_<o�_`o�_mo�o %o�oIo�o�oo�o 8J�on�o��3 �W�{�"��F� �j�|����/�ď֏�e������0��$F�ILE_FRSP�RT  ��������?�MDONLY �1|S�� 
� �)MD:_�VDAEXTP.�ZZZ1�⏹�ț�6%NO B�ack filey ���S�6P�� ���>��K�t����� '���ί]�򯁯�(� ��L�ۯp������5� ʿY�׿ Ϗ�$ϳ�H� Z��~�Ϣϴ�C��� g���ߝ�2���V��� cߌ�߰�?�����u� 
��.�@���d��߈����C�VISBCK�q�[���*.VD�����S�FR:\���ION\DAT�A\��v�S�V�ision VD ���Y�k����y� ��B�����x���1 C��g���,� P����?� Pu�(��^ ��/��M/�q/ �/>/�/6/�/Z/�/? �/%?�/I?[?�/??�?2?D?�?9�LUI�_CONFIG �}S����;O $ �3v�{S� ;OMO_OqO�O�O�I#@|x�?�O�O�O__ %\�OH_Z_l_~_�_'_ �_�_�_�_�_o�_2o DoVohozo�o#o�o�o �o�o�o
�o.@R dv����� ���*�<�N�`�r� �������̏ޏ��� ��&�8�J�\�n���� ����ȟڟ쟃���"� 4�F�X�j�������� į֯����0�B� T�f�����������ҿ �{���,�>�P�b� ���ϘϪϼ�����w� ��(�:�L�^��ς� �ߦ߸�����s� �� $�6�H���Y�~��� ����]������ �2� D���h�z��������� Y�����
.@�� dv����U� �*<�`r ����Q��/ /&/8/�\/n/�/�/ �/;/�/�/�/�/?"? �/F?X?j?|?�?�?7? �?�?�?�?OO�?BO TOfOxO�O�O3O�O�O �O�O__�O>_P_b_ t_�_�_/_�_�_�_�_ oo�_:oLo^opo�o|�o$h  x�o��c�$FLUI_�DATA ~�����a�(a�dRESUL�T 3�ep� �T�/w�izard/gu�ided/ste�ps/Expert�o=Oas���������z��Continue with Gpance�:�L�^� p���������ʏ܏� � �b-�a�e�0 �0`��cl�a?��ps� ��������ҟ���� �,�>�P��0ow��� ������ѯ����� +�=�O�a�?�1�C�U�=e�cllbs�ֿ �����0�B�T�f� xϊϜ�[��������� ��,�>�P�b�t߆߀�ߪ�i�{��ߟ�]�e�rip(pſ-�?� Q�c�u������� ������)�;�M�_� q���������������@������`�e��#pTimeUS/DST	���� ���!3E�?Enabl(�y �������	/P/-/?/Q/�b�`)�/M_q24| �/�/??)?;?M?_? q?�?�?Tf�?�?�? OO%O7OIO[OmOO �O�Ob/t/�/�/Z�~"qRegion�O 5_G_Y_k_}_�_�_�_��_�_�_�America!�#o5oGo Yoko}o�o�o�o�o�o�o��Ay�O�O3�O�_qEditor �o����������+�=� � To�uch Pane�l rs (rec_ommenp�)K� ������Ə؏���� �2�D�|�%���I[qacces oܟ� ��$�6�H��Z�l�~�����Co�nnect to� Network ��֯�����0�B�@T�f�x�����x��@!��}����,!��s �Introduct!_4�F�X�j�|ώ� �ϲ���������� 0�B�T�f�xߊߜ߮�0�������� ɿ ��"�i�{��� ������������/� A� �e�w��������� ������+=�H�3��+�O� ����� 2 DVhz�K��� ���
//./@/R/ d/v/�/�/Yk}�/ �??*?<?N?`?r? �?�?�?�?�?�?��? O&O8OJO\OnO�O�O �O�O�O�O�O�/_�/ 1_�/X_j_|_�_�_�_ �_�_�_�_oo0oBo S_foxo�o�o�o�o�o �o�o,>�O_ !_�E_����� ��(�:�L�^�p��� ��So��ʏ܏� �� $�6�H�Z�l�~���O ��s՟���� �2� D�V�h�z�������¯ ԯ毥�
��.�@�R� d�v���������п� ���ş'�9���`�r� �ϖϨϺ�������� �&�8���\�n߀ߒ� �߶����������"� 4��=��a��Mϲ� ����������0�B� T�f�x���I߮����� ����,>Pb t�E��i���� (:L^p� ������� // $/6/H/Z/l/~/�/�/ �/�/�/����/? �V?h?z?�?�?�?�? �?�?�?
OO.O�RO dOvO�O�O�O�O�O�O �O__*_<_�/?? �_C?�_�_�_�_�_o o&o8oJo\ono�o?O �o�o�o�o�o�o" 4FXj|�M___ q_��_���0�B� T�f�x���������ҏ �o���,�>�P�b� t���������Ο��� ��%��L�^�p��� ������ʯܯ� �� $�6�G�Z�l�~����� ��ƿؿ���� �2� �S��w�9��ϰ��� ������
��.�@�R� d�v߈�G��߾����� ����*�<�N�`�r� ��Cϥ�g���ύ�� �&�8�J�\�n����� ������������" 4FXj|��� �������-�� Tfx����� ��//,/��P/b/ t/�/�/�/�/�/�/�/ ??(?�1U?? A�?�?�?�?�? OO $O6OHOZOlO~O=/�O �O�O�O�O�O_ _2_ D_V_h_z_9?�?]?�_ �_�?�_
oo.o@oRo dovo�o�o�o�o�o�O �o*<N`r ������_�_�_ �_#��_J�\�n����� ����ȏڏ����"� �oF�X�j�|������� ğ֟�����0�� ��u�7�������ү �����,�>�P�b� t�3�������ο�� ��(�:�L�^�pς� A�S�e��ω��� �� $�6�H�Z�l�~ߐߢ� ���߅������ �2� D�V�h�z������ ���������@�R� d�v������������� ��*;�N`r ������� &��G	�k-�� ������/"/ 4/F/X/j/|/;�/�/ �/�/�/�/??0?B? T?f?x?7�?[�? �?�?OO,O>OPObO tO�O�O�O�O�O�/�O __(_:_L_^_p_�_ �_�_�_�_�?�_�?o !o�OHoZolo~o�o�o �o�o�o�o�o �O DVhz���� ���
���_%o�_ I�s�5o������Џ� ���*�<�N�`�r� 1������̟ޟ�� �&�8�J�\�n�-�w� Q���ů������"� 4�F�X�j�|������� Ŀ�������0�B� T�f�xϊϜϮ���� �������ٯ>�P�b� t߆ߘߪ߼������� ��տ:�L�^�p�� ���������� �� $������i�+ߐ��� ���������� 2 DVh'���� ���
.@R dv5�G�Y��}�� �//*/</N/`/r/ �/�/�/�/y�/�/? ?&?8?J?\?n?�?�? �?�?�?��?�O� 4OFOXOjO|O�O�O�O �O�O�O�O__/OB_ T_f_x_�_�_�_�_�_ �_�_oo�?;o�?_o !O�o�o�o�o�o�o�o (:L^p/_ ������ �� $�6�H�Z�l�+o��Oo ��sou����� �2� D�V�h�z������� ����
��.�@�R� d�v���������}�߯ ����ٟ<�N�`�r� ��������̿޿�� �ӟ8�J�\�nπϒ� �϶����������ϯ ��=�g�)��ߠ߲� ����������0�B� T�f�%ϊ������� ������,�>�P�b� !�k�Eߏ���{����� (:L^p� ���w���  $6HZl~�� �s�������/��2/ D/V/h/z/�/�/�/�/ �/�/�/
?�.?@?R? d?v?�?�?�?�?�?�? �?OO���]O/ �O�O�O�O�O�O�O_ _&_8_J_\_?�_�_ �_�_�_�_�_�_o"o 4oFoXojo)O;OMO�o qO�o�o�o0B Tfx���m_� ����,�>�P�b� t���������{oݏ�o ��o(�:�L�^�p��� ������ʟܟ� �� #�6�H�Z�l�~����� ��Ưد����͏/� �S��z�������¿ Կ���
��.�@�R� d�#��ϚϬϾ����� ����*�<�N�`�� ��C���g�i������ �&�8�J�\�n��� ���u��������"� 4�F�X�j�|������� q�������	��0B Tfx����� ����,>Pb t������� /����1/[/�/ �/�/�/�/�/�/ ?? $?6?H?Z?~?�?�? �?�?�?�?�?O O2O DOVO/_/9/�O�Oo/ �O�O�O
__._@_R_ d_v_�_�_�_k?�_�_ �_oo*o<oNo`oro �o�o�ogOyO�O�O�o �O&8J\n�� �������_"� 4�F�X�j�|������� ď֏�����o�o�o Q�x���������ҟ �����,�>�P�� t���������ί�� ��(�:�L�^��/� A���e�ʿܿ� �� $�6�H�Z�l�~ϐϢ� a���������� �2� D�V�h�zߌߞ߰�o� �ߓ��߷��.�@�R� d�v��������� ����*�<�N�`�r� �������������� ��#��G	�n�� ������" 4FX�|��� ����//0/B/ T/u/7�/[]/�/ �/�/??,?>?P?b? t?�?�?�?i�?�?�? OO(O:OLO^OpO�O �O�Oe/�O�/�O�O�? $_6_H_Z_l_~_�_�_ �_�_�_�_�_�? o2o DoVohozo�o�o�o�o �o�o�o�O_�O%O _v������ ���*�<�N�or� ��������̏ޏ��� �&�8�J�	S-w� ��cȟڟ����"� 4�F�X�j�|�����_� į֯�����0�B� T�f�x�����[�m�� ��󿵟�,�>�P�b� tφϘϪϼ������� ���(�:�L�^�p߂� �ߦ߸������� ￿ ѿ�E��l�~��� ����������� �2� D��h�z��������� ������
.@R �#�5�Y��� �*<N`r ��U�����/ /&/8/J/\/n/�/�/ �/c�/��/�?"? 4?F?X?j?|?�?�?�? �?�?�?�??O0OBO TOfOxO�O�O�O�O�O �O�O�/_�/;_�/b_ t_�_�_�_�_�_�_�_ oo(o:oLoOpo�o �o�o�o�o�o�o  $6H_i+_�O_ Q����� �2� D�V�h�z�����]o ԏ���
��.�@�R� d�v�����Y��}ߟ 񟵏�*�<�N�`�r� ��������̯ޯ𯯏 �&�8�J�\�n����� ����ȿڿ쿫���ϟ �C��j�|ώϠϲ� ����������0�B� �f�xߊߜ߮����� ������,�>���G� !�k��Wϼ������� ��(�:�L�^�p��� ��S߸�������  $6HZl~�O� a�s����� 2 DVhz���� ����
//./@/R/ d/v/�/�/�/�/�/�/ �/���9?�`?r? �?�?�?�?�?�?�?O O&O8O�\OnO�O�O �O�O�O�O�O�O_"_ 4_F_??)?�_M?�_ �_�_�_�_oo0oBo Tofoxo�oIO�o�o�o �o�o,>Pb t��W_�{_��_ ��(�:�L�^�p��� ������ʏ܏��� $�6�H�Z�l�~����� ��Ɵ؟꟩��/� �V�h�z�������¯ ԯ���
��.�@��� d�v���������п� ����*�<���]�� ��C�EϺ�������� �&�8�J�\�n߀ߒ� Q������������"� 4�F�X�j�|��Mϯ� q��������0�B� T�f�x����������� ����,>Pb t�������� ����7��^p� ������ // $/6/��Z/l/~/�/�/ �/�/�/�/�/? ?2? �;_?�?K�?�? �?�?�?
OO.O@ORO dOvO�OG/�O�O�O�O �O__*_<_N_`_r_ �_C?U?g?y?�_�?o o&o8oJo\ono�o�o �o�o�o�o�O�o" 4FXj|��� ����_�_�_-��_ T�f�x���������ҏ �����,��oP�b� t���������Ο��� ��(�:����� A�����ʯܯ� �� $�6�H�Z�l�~�=��� ��ƿؿ���� �2� D�V�h�zό�K���o� �ϓ���
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� ������������ ��#���J�\�n����� ������������" 4��Xj|��� ����0�� Q�u7�9��� ��//,/>/P/b/ t/�/E�/�/�/�/�/ ??(?:?L?^?p?�? A�?e�?�?�/ OO $O6OHOZOlO~O�O�O �O�O�O�/�O_ _2_ D_V_h_z_�_�_�_�_ �_�?�?�?o+o�?Ro dovo�o�o�o�o�o�o �o*�ON`r �������� �&��_/o	oS�}�?o ����ȏڏ����"� 4�F�X�j�|�;���� ğ֟�����0�B� T�f�x�7�I�[�m�ϯ ������,�>�P�b� t���������ο��� ��(�:�L�^�pς� �Ϧϸ����ϛ����� !��H�Z�l�~ߐߢ� ����������� �߿ D�V�h�z������ ������
��.����� �s�5ߚ��������� ��*<N`r 1������ &8J\n�?� �c������/"/ 4/F/X/j/|/�/�/�/ �/�/��/??0?B? T?f?x?�?�?�?�?�? ��?�O�>OPObO tO�O�O�O�O�O�O�O __(_�/L_^_p_�_ �_�_�_�_�_�_ oo $o�?EoOio+O-o�o �o�o�o�o�o 2 DVhz9_��� ���
��.�@�R� d�v�5o��Yo��͏� ���*�<�N�`�r� ��������̟��� �&�8�J�\�n����� ����ȯ��я����� �F�X�j�|������� Ŀֿ�����ݟB� T�f�xϊϜϮ����� ������ٯ#���G� q�3��ߪ߼������� ��(�:�L�^�p�/� ���������� �� $�6�H�Z�l�+�=�O� a��������� 2 DVhz���� ����
.@R dv������� ����/��</N/`/r/ �/�/�/�/�/�/�/? ?�8?J?\?n?�?�? �?�?�?�?�?�?O"O ��/gO)/�O�O�O �O�O�O�O__0_B_ T_f_%?w_�_�_�_�_ �_�_oo,o>oPobo to3O�oWO�o{O�o�o (:L^p� �����o� �� $�6�H�Z�l�~����� ��Ə�o珩o��o2� D�V�h�z������� ԟ���
���@�R� d�v���������Я� ����׏9���]�� !�������̿޿�� �&�8�J�\�n�-��� �϶����������"� 4�F�X�j�)���M��� �߅�������0�B� T�f�x������� ������,�>�P�b� t���������{��ߟ� ����:L^p� ������  ��6HZl~�� �����/�� ��;/e/'�/�/�/�/ �/�/�/
??.?@?R? d?#�?�?�?�?�?�? �?OO*O<ONO`O/ 1/C/U/�Oy/�O�O_ _&_8_J_\_n_�_�_ �_�_u?�_�_�_o"o 4oFoXojo|o�o�o�o �o�O�O�O	�O0B Tfx����� ����_,�>�P�b� t���������Ώ��� ���o�o�o[��� ������ʟܟ� �� $�6�H�Z��k����� ��Ưد���� �2� D�V�h�'���K���o� Կ���
��.�@�R� d�vψϚϬϾ�Ͽ�� ����*�<�N�`�r� �ߖߨߺ�y��ߝ��� ��&�8�J�\�n��� �������������� 4�F�X�j�|������� ����������-�� Q������ ��,>Pb !�������� //(/:/L/^// A�/�/y�/�/ ?? $?6?H?Z?l?~?�?�? �?s�?�?�?O O2O DOVOhOzO�O�O�Oo/ �/�/�O_�/._@_R_ d_v_�_�_�_�_�_�_ �_o�?*o<oNo`oro �o�o�o�o�o�o�o �O_�O/Y_�� �������"� 4�F�X�o|������� ď֏�����0�B� T�%7I��mҟ �����,�>�P�b� t�������i�ί�� ��(�:�L�^�p��� ������w��������� $�6�H�Z�l�~ϐϢ� ���������ϻ� �2� D�V�h�zߌߞ߰��� ������
�ɿۿ�O� �v��������� ����*�<�N��_� �������������� &8J\�}?� �c�����" 4FXj|��� ����//0/B/ T/f/x/�/�/�/m�/ ��/�?,?>?P?b? t?�?�?�?�?�?�?�? O�(O:OLO^OpO�O �O�O�O�O�O�O _�/ !_�/E_?	_~_�_�_ �_�_�_�_�_o o2o DoVoOzo�o�o�o�o �o�o�o
.@R _s5_��mo�� ���*�<�N�`�r� ������gȍޏ��� �&�8�J�\�n����� ��c��џ���"� 4�F�X�j�|������� į֯������0�B� T�f�x���������ҿ �������ٟ#�M�� tφϘϪϼ������� ��(�:�L��p߂� �ߦ߸������� �� $�6�H���+�=ϟ� a���������� �2� D�V�h�z�����]��� ������
.@R dv���k�}������$FMR2_GRP 1���� �C4  B��	 ��9K6/F@ a@�6�G�  �Fg��fC�8R�y?ǀ  ��66��X���875t���5���5`{+�yA�  /�+BH�w-%@S339%�5[/l-6@6!�/xl/�/�/ �/�/?�/&??J?5?�G?�?k?�?��_C_FG �TK��?�? OO�9NO {
F0FA� K@�<RM_CHKTYP  ��$&� ROM�a@_MINg@������@�R XS�SB�3�� 7�O���C��O�O�5TP_DEF_OW  ���$WIRCOM�f@_�$GENO�VRD_DO�F̾�E]TH��D dzbUdKT_ENB7_{ KPRAVCu��G�@ �Y �O�_�?oyo&onI* �QOU�NAIRI<�@��oGo�oX�o�o��C�p3���O:��B��+sL�i�O�PSMT���Y(�@
t�$�HOSTC�21���@�5 kMC��R{����  27.0z0�1�  e� ]�o�������K�ď֏���������	anonymous!� O�a�s����� �4��������D�!� 3�E�W�i��������� ï柀�.���/�A� S���课�П���� Ŀ����+�r�O�a� sυϗϺ������� ��'�n��������� ��ڿ����������F� #�5�G�Y�k���υ� ����������B�T�f� C�z�g��ߋ������� �����	-P��� ��u������ (�:�<)p�M_q ��������/ $ZlI/[/m//�/ ����//�/D!? 3?E?W?/?�?�?�? �?�/�?./OO/OAO SO�/�/�/�/�?�O? �O�O__+_r?O_a_ s_�_�_�O�?O�_�_�oo'o�t�qENT� 1�hk P!\�_no  �p\o �o�o�o�o�o�o�o �o:_"�F� j�����%�� I��m�0���T�f�Ǐ ��돮��ҏ3���,� i�X���P���t�՟�� ៼�
�/��S��w� :���^�������������ܯ=� �QUI�CC0J�&�!1�92.168.1'.10c�X�1��v�8��\�2�ƿؿ9��!ROUTER�:��!��a���PCJOG��e�/!* ��0��U�?CAMPRT�϶�c!�����RTS����x� !So�ftware O�perator PanelU߇����7kNAME !~Kj!ROBO�����S_CFG 1��Ki ��Auto-st�arted�DFTP�Oa�O�_�� �O����������E_� .�@�R�u�c�	����� ������cN:�L�^�; r���R������ ��%H�[ m���jO|O�O �O4!/hE/W/i/{/ �/T�/�/�/�/�// �//?A?S?e?w?�?� ���??�?</O+O =OOO?sO�O�O�O�O �?`O�O__'_9_K_ �?�?�?�?�O�_�?�_ �_�_o#o�OGoYoko }o�o�_4o�o�o�o�o f_x_�_g�o� �_�����o�� -�?�Q�tu������ ��Ϗ�(:L^`� 2��q����������� ݟ���%�H�ʟ[� m����������� � ί4�!�h�E�W�i�{� ��T���ÿտ�
�� ��/�A�S�e�w����_ERR �����ϗ�PDUSIZW  �^6�����>��WRD ?�(����  guestƀ��+�=�O�a���S�CD_GROUP� 3�(� ,��"�IFT��$PA��OMP�� n��_SH��ED��w $C��COM���TTP_AUTH� 1��� <!�iPendan�m�x�#�+!KAREL:*x���KC�������VISION SET��(����?�-�W�R���v������������������G�CT_RL ���a��
�FFF�9E3��FR�S:DEFAUL�T�FANU�C Web Server�
tdG� ���/� 2D�V��WR_CON�FIG ���������ID�L_CPU_PC�� �B���� ;BH�MIN���~�GNR_IO�������ȰHMI_EDIT ���
 ($/C/��2/ k/V/�/z/�/�/�/�/ �/?�/1??U?@?y? d?�?�?./�?�?�?�? OO?OQO<OuO`O�O �O�O�O�O�O�O__�;_�NPT_SI�M_DO�*N�STAL_SCR�N� �\UQTPMODNTOL�Wl[�RTYbX�qV\�K�ENB�W����OLNK 1�����o%o7oIo[o�moo�RMASTE���Y%OSLA�VE ��ϮeRAMCACHE�o��ROM�O_CFG�o�S�cUO'��b?CMT_OP�  "��5sYCL�ou� _ASG 1����
 �o��� ����"�4�F�X��j�|����kwrNUMj����
�bIP�o��gRTRY_CNx@uQ_UPD�Êa��� �bp�bA��n��M��аP}T{?��k ��._ ������ɟ۟퟈S�� �)�;�M�_�q� ��� ����˯ݯ�~��%� 7�I�[�m�������� ǿٿ�����!�3�E� W�i�{�
ϟϱ����� ���ψϚ�/�A�S�e� w߉�߭߿������� ��+�=�O�a�s�� �&���������� ��9�K�]�o�����"� �������������� GYk}��0� ����CU gy��,>�� �	//-/�Q/c/u/ �/�/�/:/�/�/�/? ?)?�/�/_?q?�?�? �?�?H?�?�?OO%O 7O�?[OmOO�O�O�O DOVO�O�O_!_3_E_ �Oi_{_�_�_�_�_R_ �_�_oo/oAo�_�_ wo�o�o�o�o�o`o�o +=O�os� ����\n�� '�9�K�]��������ාɏۏi�c�_ME�MBERS 2��:�  � $:� ����v���1���RCA_ACC 2���  � [}�M 4|�� ;� �_� )5�l�l�%l���� ����� {���a�BUF�001 2�n�=� ��??�  ��=�=��  �>>��V��=8=8���=�=����?H?H.�V>(�>(.��
���=��=�  �@��@�N�VK0K�0  � **���@
���@��@m��j��u0u~]��8=�=���_x?�?؆��J�;����8H����oxX�XM������K�L��8��Mu�08�<x�T7�M�7���u0��g��u0c��@���u0��(�4�B�N��[�i�v򤄪���򤷢���������Z���z�z��z�*z�Vu0?��5@��=�=ZU��I����V���������X�%X�����ߙ2��� �"�4�F�X�j�|��� ����ĭ��ءڡࡍ� ������������� 	���������!��� )���1���9���A��� I���Q���Y�����i� ��q���y������҉� �ґ��ҙ��ҡ��ҩ���Ϳ߿�3���l� �l���"��*�� 2�l�9�>�B�>�J�>� R�l�Y�^�b�l�i�n� r�n�z�n��n��l� �����������l� �����������T�ƣ ��Ѡ��٢��l���� ����������� ��!�/���1�?���A� O���Q�_�����i�w� ��y��ӎ򉲗ӎ� �ӎ�Ў�[������� ��������������~a�CFG 2�n�G 4��l�l��<l�47%�a�H�IS钜n� ��� 2025-�11-29l� 珚�������l�;g� � % ��� /i�B���r� ������// K]J/\/n/�/�/�/ �/�/�/�/#/5/"?4? F?X?j?|?�?�?�?�? �/?�?OO0OBOTO fOxO�O�O�?�?�?�O �O__,_>_P_b_t_ �_�O�O�_�_�_�_o o(o:oLo^oL	��[ m�o�o�o�o�o�!3!: c��2
l�d��-Zq�_�_< �������� +��_t�s������� ��͏ߏ���L�^� K�]�o���������ɟ ۟�$�6�#�5�G�Y� k�}�������ů��� ����1�C�U�g�y� ����ԯ������	� �-�?�Q�c�u�coue �Ѐo�o�o��������"�4�F�X�!o�  ��}Ӳ�Ŀa������� ����,�>�P�ߙ� �ߘ���������� �(�:�q��p����� ���������� I� [�HZl~��� ���!3 2D Vhz����� 
//./@/R/d/�v/�/�/��u`I_C�FG 2��� �H
Cycle� Time�B�usy�Idl��"�min�+�1Up�&��Read�'D�ow8? 2��#Count�	ONum �"����<��~�qaPROmG�"�������)/softp�art/genl�ink?curr�ent=menu�page,1133,1�/OO/OAO�3b5leSDT_ISOLC  ���� �@�.J23�_DSP_ENB�  vK0�@IN�C ��M�Ä@A�   ?�  =���<#�
�A>�I:�o �A_`_���O<_�GOB�0�C�C5�FVQG_�GROUP 1��vK<Zq<���C��_D_?��?�_��Q�_o.o@o@�_dovo�o�o�,_�NYG_IN_AU�TOcT�MPOSR�E^_pVKANJI_MASK v�Hq�RELMON ��˔?��y_ox�@����.6r�3��7��C���u�o�DK�CL_L�`NUM��@�$KEYLO�GGING������Q�E�0LANGU�AGE ���~��DEFA�ULT ����LGf�!��:2����x�@{�80H � ���'0�� +
������GOUF� ;��
��(�UT1:\��  �-�?�Q�h�u����������ϟ�����(�g4�8i�N_DISP ��O8�_��_��LOCTOL����Dz|�A�A���GBOOK ����d�1
�
�۠X����#�5�G�Y�`i���3{�W�	��@쉞QQJ¿Կ1���_BUFF 2�NvK ���25�
�ڢVB&�7 C�ollaborativ�=�OΗώ� �ϲ���������'�� 0�]�T�fߓߊߜ��?DCS ��9�B �Ax�����%�-�?�|Q���IO 2���� ���Q� ������������ �*�<�N�b�r����� ����������&�:e�ER_ITMsNd�o����� ��#5GYk }����������hSEV��M.dTYPsN�c/pu/�/
-�aRST5����SCRN_FLW 2�s��0��� �/??1?C?U?g?�/�TPK�sOR"��NGNAM�D��~�N�UPS_ACR� ��4DIGI�8~+)U_LOAD[P�G %�:%T_NOVICEt?���MAXUALR�M2��1���E
LZB�1_P�5�0 ��4y�Z@CY��˭�O�+���ۡ�D|PP 2]�˫ ��	R/ _
_C_._g_y_\_�_ �_�_�_�_�_�_oo ?oQo4ouo`o�o|o�o �o�o�o�o)M 8qTf���� ���%��I�,�>� �j�����Ǐُ���� �!���W�B�{�f� ������՟����ܟ� /��S�>�w���l��� ��ѯ��Ư��+���O�a�D���p���RHD�BGDEF ��E�ѱO��_LDX�DISA�0�;c�M�EMO_AP�0E� ?�;
  ױ��3�E�W�i�{ύ���ϱ�Z@FRQ_C_FG ��G۳�A ��@��Ô�<��d%�� ������Bݯ�K���*i�/k� **:tҔ�g�y�ߔ��� �����������J� ���Es�J d������,(H���[���� �@�'�Q�v�]����� ����������*�NPJISC 1��9Z� ������ܿ������	Zl_MSTR �#-~,SCD 1�"��{����� ���//A/,/e/ P/�/t/�/�/�/�/�/ ?�/+??O?:?L?�? p?�?�?�?�?�?�?O 'OOKO6OoOZO�O~O �O�O�O�O�O_�O5_  _Y_D_i_�_z_�_�_ �_�_�_�_o
ooUo @oyodo�o�o�o�o�o �o�o?*cNl�MK���;�љ$MLTAR�M���N��r� ��հ��İM�ETPU��zr���CNDSP_A�DCOL%�ٰ0�C�MNTF� 9�F�Nb�f�7�FSTLqI��x�4 �;�ڎ�s����9�PO�SCF��q�PR�PMe��STD�1ݶ; 4�#�
v��qv�����r��� �����̟ޟ ��� V�8�J���n���¯������9�SING_CHK  ���$MODA����t�{�~2�DEV �	�	MC:>f�HSIZE��zp��2�TASK �%�%$1234?56789 ӿ��0�TRIG 1�; lĵ�2ϻ�0!�bϻ�YP�����H�1�EM_IN�F 1�N�`�)AT&FV0�E0g���)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ��2��H6� ^���Rφ��A�߶� q�������� ��5� �����ߏ�B߳��� ��������1�C�*� g��,��P�b�t��� ���R�?���u 0��������� ������M q�� �Z���/�%/ ��[/ 2�/�/ h�//�/�/�3?�/ W?>?{?�?@/�?d/v/ �/�/O�//OAOx?eO ?�ODO�O�O�O�O_��NITORÀG �?z�   	�EXEC1~s&R2*,X3,X4,X5,X���.V7,X8,X9~s 'R�2�T+R�T7R�TCR �TOR�T[R�TgR�TsR��TR�T�R�S2�X2��X2�X2�X2�X2��X2�X2�X2�X2*h3�X3�X37R2��R_GRP_SVw 1��� (��=�ĝ<Ŧ��=�9P�w�������jc�a���_D�B���cI_ON_DB<��@�>zq  �2p��S;Y�1u�2p�>w+�ZpyZpzY��@?N   �rp]p�@yq$�rY�-ud1�����8��PG_JOG ��ʏk�
�2��:�o�=���?����0�B��~\�n��������0H�?��C�@�ŏ׏����  ������qL_NAME �!ĵ8��!�Default �Personal�ity (fro�m FD)qp0�R�MK_ENONL�Y�_�R2�a 1��L�XLy�8�gpl d�� ��şן�����1� C�U�g�y��������� ӯ���	��n�
�<� N�`�r���������̿޿� :��)� ;�M�_�qσϕϧϹ� ��������%�7�I� [�m�ߑߣߵ����� �����!�3�E�W�i� {������������ ��/�A�S�e�w��� ������������+��<�Sew� ������^��A�a��B�Bw��Pf�� ����/!/3/E/ W/i/{/�/�/�/�� �/�/??/?A?S?e? w?�?�?�?�?�?�?�? �/�/+O=OOOaOsO�O �O�O�O�O�O�O__�'_9_&O�S���x_�]�rdtS���_�] �_�_�W�����S"oe_8oXoa ��qo goyo�o�o�o�o�ouP��p"|����	`@[oUgy8qK�A\�p���s� A �P�y@h�Q�Q��"����Tk\$���  ��P�PE~�xC�  �I� @oa�<o��p�������@ߏ
f�Q,������0���PCr� �� 3r �.� @D7�  A�?�G�-��?.I�.@I��A����  ;�	�lY�	 �X  ������� �,� � �����uPK��o�����]K���K]�K	�.��w�r_	�<���@
�)�b�x1�����I�Y�����T;fY��{S���3�����I�>J���;Î?�v�>��=@��'���E��Rѯע�Z���wp��u�� �D!�3��7pg�  �  ��9�͏W���	'� �� u�I� ?�  ��u���:�È��È=���ͱ���@���ǰ�3��{3��E�&���N�pC�  �'Y�&�Z�i�b�@f�i�n�C����I��C����b���r���`����B �p�Ŕq���}ر�.DzƏ<ߛ�`�K�p�ܖ����������А 4�P����.z��d � �Pؠ?��ff�_��	�� 2p>�P���8.f�t�C>L���U���(.��P���٨���������� x��;e��m��KZ;�=�g;�4�<<a����%�G��3�|���p?fff?ذ�?&S���@=0e�?��q��y�r N�Z���I���G���7� ��(�����!E0 iT�����x��F�p���#�� D��w��� ����//=/(/ a/L/�/p/��/�p� 6�/Z#?�/ ?Y?k? }?��?�?>?�?�?�? �?�?1O�����KD�y�{CO�OO�O��ɃذO�O�O�O�y����J��}�DD1���.�D��@�AmQa���9N,ȴA;��^@��T@|j�@$�?�V��>�z�ý���=#�
>\�)?��
=�G}�-]�{=����,��C+�ןBp���P��6���C98R����?N@��(���5-]G�p��Gsb�F�}��G�>.E�V�D�Kn����I�� F�W��E��'E����D��;n����I��`E����G��cE�vmD���-_�oQ_ �o�o�o �o$H 3X~i���� �����D�/�h� S���w��������я 
���.��R�=�v�a� s�����П����ߟ� �(�N�9�r�]����� ����ޯɯۯ���8� #�\�G���k������� ڿſ���"��F�1� C�|�gϠϋ��ϯ����������P(�Q343�] �����Q�	�x9�Oߵ53~�mm��aҀ5Q�߫�a�Ǔ����ߵ1��������1��U�C�(y�g��%P�P���!�/��'���
���.������4�;�t� _��������������� :%��/�/d������� �7%[I�m���027� � B�S@J@�CH#PzS@�0@ZO/1/@C/U/g/y/�-�#���/�/�/�/�/�3?��3�� @�3��0�0�13��5
 ?f?x?�?�? �?�?�?�?�?OO,Op>OPO�Z@1 �������c/�$MR�_CABLE 2�ƕ� ��TT�����ڰO���O �Y�@���C_���_ O_u_7_I__�_�_�_ �_�_o�_�_oKoqo 3oEo{o�o�o�o�o�o �o�o�oGm/�K!�"���O�����ذ�$�6����*Y�** �COM� ȖI�����"43�%% �2345678901���� ��Ï��R� � !� �!�
���Mnot sent b���W��TE�STFECSAL?GR  eg)
!�d[�41�
k�������$pB����������� 9UD1�:\mainte�nances.xsmlğ�  C:��DEFAU�LT�,�BGRP {2�z�  ����%  �%!1s�t cleani�ng of co�nt. v�il�ation 56
��ڧ�!0�����+B��*�����+���"%��mech���cal che{ck1�  �k�!0u�|��ԯ�����Ϳ߿�@���rollerS�e�w�ū��m�ϑϣϵ�@��Basic q�uarterly�*�<�ƪ,\�)�;�0M�_�q�8�MJ���� "8��� ����� �����+�=�C�g�ߋ����߹��������@�Overhau��6���?� x� I�P����}���������� $n������aI l�ASew���� �� �+= O�s����� ��/R�9/�(/ ��/�/�/�/�//�/ �/N/#?r/G?Y?k?}? �?�/�???�?8?O O1OCOUO�?yO�?�? �O�?�O�O�O	__jO ?_�O�Ou_�O�_�_�_ �_�_0_oT_f_;o�_ _oqo�o�o�o�_�oo ,oPo%7I[m �o��o�o��� �!�3��W���� ����ÏՏ�6���� l����e�w������� ��џ�2��V�+�=� O�a�s������ͯ ����'�9���]� ������⯷�ɿۿ� ��N�#�r���YϨ�}� �ϡϳ������8�J� �n�C�U�g�yߋ��� �������4�	��-� ?�Q��u������ߞ� ��������f�;��� ������������� ��P���t�I[m ������: !3EW�{� �� ���// lA/��w/��/�/�/�/�/X*�"	 X`�/?.?@?�)B a/ o?�?�?�?�?�?�?�? �?O#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_��_�_�_�_�_	oo"� Џ!?�  @�! M?HoZolo��&4o�o�o�o�(�*�o** F�@ i!k&�`o'9��o]o���� �/^&�o����� /�A�S�e���#��� ��я�����+�q� ����7�������k�͟ ߟ��I�[���K�]� o���C�����ɯ���o$�!�$MR_HIST 2�g%}#�� 
 \7"�$ 23456789013�;���b2�90/����[��� ./����ǿٿF�X� j�!�3ρϲ���{��� ������B���f�x� /ߜ�S����߉��߭� �,���P��t��=����$�SKCFM�AP  g%�&��b
�� �����ONREL � �$#������E�XCFENB�
8����&�FNC-���JOGOVLIM��d#�v���KEY��y���_PA�N������RUN�i�y���SFSPDTYPM�����SIGN��T1�MOTk����_�CE_GRP 1�g%��+�0�o w�#d���� ��&�6\ �7y�m��� /�4/F/-/j/!/t/ �/�/�/{/�/�/�/?��+��QZ_EDI�T
����TCOM_CFG 1���a0�}?�?�? 
^1�SI �N����?�?���?$O�����?XO78T_A�RC_*�X�T�_MN_MODE�
�U:_SPL�{O;�UAP_CP�L�O<�NOCHE�CK ?�� �� _#_5_G_ Y_k_}_�_�_�_�_�_��_�_oo��NO_?WAIT_L	S76> NTf1����%z��qa_ERRH2�������?o�o�o�o��OGj�@�O�cӦm| 4|��GA@g��A�����PF������W�-�`���<���?����)��n�bPA�RAM�b����vHO��w
�.�@� = n�]�o�w�Q� ����������Ϗ�)���w�[�m� ������ODRDSP��C8�OFFSET_CARI0�Oǖ�DISԟœS_AΖ@ARK
T9OPEN_FILE���1T6�0OPTION_IO����K��M_PRG %���%$*����'�WmO��Nsq�ǥ�� ���u����	 �����Ӧ�����R�G_DSBL  �����jN���R�IENTTO�f��C�����A ���U�@IM_DS����r��V��LCT �{mP2ڢ�3̹���dҩ��_PEX��@���RAT�G �d8��̐UP Sװ�:����Sϰe�Kωϗ��$�r2�G�L�XL;Ț�l㰂� ������'�9�K�]� o߁ߓߥ߷�������@���#�5�G���2�� v�������������e�B�T�f� x��������������� ,>Pbt� ������ (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? �q1�~?�?�?�?�?�?��?�?O O2ODO�yA�a�m?~N��~O�O�P�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�O�Oo $o6oHoZolo~o�o�o �o�o�o�o�o �_ oVhz���� ���
��.�@�R�0d�QOES������
B�d�ӏ�ʏ� �������Y�D�}�0��r���������ԟ ڟ���p���=�M��q�	`��������c�:�o�¯ԯ�����A�  P�k�C�C�ڰ"ڰ����O��/  ���-���~)�C�  �t� k���g�����Կ��ѿ�
�5���^:�ĳ�OU���� �� ��H��n�� o� ^�\�� @D�  p�?��v�\�?:px�:qC�4r�p�(��  ;��	l��	 ��X  ������� �,? � ��������Hʪ�����H���Hw�_zH�����8�B���B�  �Xѐ�`�o�*��3�	���t�>u���fC{�����:pB\�
��Ѵ9:qK�t�� ����$����*��� DP��^��b�g  �  �h������)�	'� � ���I� � � ��'�=��q�����t�@��@��!�b��^;b�t��U�(�N��r�  '���E�C�И�t�C��И��ߗ���jA�@!�����%�B�� ���,���H:qDz �k�ߏz���w�����А 4P��D�:uz:���	f�~�?�ff'�&8� ]�mb�8:p��>L��H���$�(:p�P���	������:� �x�;e�m"��KZ;�=g;�?4�<<���E/�Tv��b���?offf?�?&� �)�@=0�%?��%`9��}!��$� x��/v��/f'��W,? ?P?;?t?_?�?�?�? �?�?�?O�?(OOLO �/�/�/EO�OAO�O�O �O�O_�O_H_3_l_ W_�_{_�_�_1��_A� ��eO+o�ORooOo�o �o�oK/�o�omo�o@*'`+�,�zt���CL�H��}?�����
������u����#D1�/n�t��p�qޜ�@I�h~,���A;�^@���T@|j@$��?�V�n�z��ý��=#��
>\)?���
=�G�����{=��,���C+��Bp�����6��C98R���?}p���(��5���G�p�Gsb��F�}�G�>�.E�VD�K�L����I��� F�W�E���'E���D���;L����I���`E�G���cE�vmD���\�՟��ҟ���/� �S�>�w�b������� ѯ�������=�(� :�s�^���������߿ ʿ�� �9�$�]�H� ��lϥϐϢ������� ��#��G�2�W�}�h� �ߌ��߰�������� 
�C�.�g�R��v�� �������	���-�� Q�<�u�`�r������� ������'M�=(�34�]O!����8h~�%3�~�m����5qQ������<�!���  �`N�r��	eP@"P��Q�_/V�/9/$/]/H)����c/j/�/�/�/�/�/ �/�/!??E?0?i?T?�"&�_�_�?�?�8� �?�?O�?OBO0OfO TO�OxO�O�O�O�Oy2f?_  B��p,Y�$QCHR�z�p@�N_`_r_�_�_�_�]c�O�_�_oo�+o?�Bc� @*d4�QqJc�D
 2o �o�o�o�o�o�o %7I[m��oa� �����c/��$PARAM_MENU ? ��  �DEFPU�LSE��	WAITTMOUT�{�RCV� �SHELL_WR�K.$CUR_S�TYL�p"�OsPT8Q8�PTBM��G�C�R_DECSN�p�V<������ �����-�(�:�L��u�p��������qSS�REL_ID  ���̕USE�_PROG %��z%���͓CCR��pޒ��s1�_HO�ST !�z!6�s�+�T�=���V��h���˯*�_TI�ME�rޖF��pGDEBUGܐ�{͓�GINP_FLM3SK��#�TR2�#�WPGAP� ��_�b�CH1�"�TYPE�|�P����� ���0�Y�T�f�x� �ϜϮ���������� 1�,�>�P�y�t߆ߘ� �߼�����	���(��Q�L�^�p��%�WO�RD ?	�{
 �	PR�p#�MAI��q"SU�d���TE��p#��	91���COLn%��!���L�� !���F�d�TRA�CECTL 1�v �q �_� �#��|��_�DT Q� ���z�D � 7�La��k` ������������� 1CUgy�� �����	- ?Qcu���� ���//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�O__ /_A_S_e_w_�_�T� �_�_�_�W�� �Uoo*o<oNo`oro �o�o�o�o�o�o�o &8J\n�� �������"� 4�F�X�j�|������� ď֏�����0�B� T�f�x���������ҟ �����,�>�P�b� t���������ί�� ��(�:�L�^�p��� ������ʿܿ� �� $�.�oP�b�tφϘ� �ϼ���������(� :�L�^�p߂ߔߦ߸� ������ ��$�6�H� Z�l�~�������� ����� �2�D�V�h� z��������������� 
.@Rdv� ������ *<N`r��� ����//&/8/ J/\/n/Dϒ/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6H Zl~����� ��� �2�D�V�h��z����������$P�GTRACELE�N  ��  �������Ά_UP ������������΁_CFG ����烸�

���*�*�D�O���>O�  �O���DEFSPD e�������΀�H_CONFIG� ���� �����dĔ�݂ 	��ǑP^�a�㑹�ۂ΀IN�TROL ��=�8^����PE��೗����*�ÑO�΀L�ID���	T�L�LB 1ⳙ ���BӐB4��O� 䘼�����Q� << ��?������ �M�3�U���i����� ����ӿ��	�7�T�Ϣk�b�tϡ�诚���������S�GRP� 1爬���@�A!���4I����A �Cu��C�OCjVF�/��Ȕa�z���ÑÐ�t��ޯ�s���´�ӿߨ�B �����������A��S�&�B34�`_������j�� ��������	�B�-����Q���M�������  Dz����.��� ��&L7p[� ������6�!Zh)w
V�7.10beta�1*�Ɛ@�*��@�) @�+�A Ē?���
?fff>�����B33A��Q�0�B(��A���AK��h ����//'/9/
P�p*�W�ӑ�n/��/�%���R�f?h����*��� P2�LR��/�/�/�/��/H?�Ĕ�I�u �&:���?��x?�?A����P!\3 Bu�B���?�5BH�3[4b��o��4��[4R5��/B\3x3Dx�?@YO�?aOkO}O�<<� R@��O�C�O�O�O�O��DA�X�KNOW_�M  Z�%�X�SoV 賚ڒ ���_�_�_?�_�_��_o����W�M+�鮳� ��	<�3#���_�o�\~=��
]bV4�@u��u��e�o�l�,�X�MR+��JmT�3?��W�1C{�OADBANFWDL_�V�ST+�1 1����P4C��� [��i/����� ?�1�C���g�y����� ���ӏ�*�	��`�?�Q�c��w2�|Va��up�<ʟ���p3 ��Ɵ؟Ꟃw4��+�=��w5Z�l�~�����w6����ѯ㯂w7  ��$�6��w8S�e�Xw����wMAmp�������OVLD � ��yo߄rP�ARNUM  ��{+þ�?υqSCH�� �
��X���{s��UPDX�)ź�|�Ϧ�_CMP_@`����p|P'yu�E�R_CHK����yqbb3��.�RS8pp?Q_MOm���_}ߥ�_RES_G�p쩻
�e��� ��0�#�T�G�x�k�}� �������������������������:� Y�^���Y�y������� �������������� ��R�6UZ�ӥ��u����V 1���FvpVa@k�p���THR_INR�p��(byudMA�SS Z)MN�GMON_QU?EUE �uyvTup\!��N�UZ�qNW��END��߶EXE�����BE���OPT�IO��ۚPROGRAM %z�%��~ϘTA�SK_I��.OCFG �z+�n/^� DATACc�+�1#s2ae?"? 4?F?X??|?�?�?�?��?o?�?�?OO�/IWNFOCc��-�� �?wO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_:GFD���, 	��!��K�_�!�)fN!fECNB��0m��Pf2Yo�khG�!2�0k �X,		d�=���·o���e�a$��pd��i�i�g_E?DIT ��/%�7����*SYS�TEM*upV9.�40107 cr7�/23/2021� A��Pw���PRGADJ_�p  h $X|[�p $Y�xZ�xW�xқtZқt?SPEED_�p�p�$NEXT_C�YCLE�p���q�FG�p ���pALGO_V� �pNYQ_F�REQ�WIN_�TYP�q)�SIuZ1�O�LAP�r�!�[��M+����qC?REATED�r��IFY�r@!NAM��p%h�_GJ�S�TATU��J�DE�BUG�rMAIL�TI����EVE<U��LAST������tELEM� �� $ENAB<�rN�EASI򁼁�AXIS�p$P�߄�����qROT�_RA" �rMAX� ��qE��LC�A�B
���C D_L9VՁ`�BAS��`��1�{���_� ��Y$x���RM� RB��;�DIS����X_cSPo�΁�� �u|�P� | 	�� 2 \�AN�� �;����8�Ӓ�� �0�PAYLO��3�V�_DOU�qS���p��tPREF� �( $GRID*�E
���R����Y�  �pOTO|ƀ�q  �p℄!�p��k�OXY�� � $L��_PO|�נVa.�SRV��)����DIRECT_1T� �2(�3(�4(�U5(�6(�7(�8����F��A�� �$VALu�GRGOUP����qF�_� !���@!�������RAN泲���R��/���TOTA��F���PW�I=!%�REGEN#�8����� ��/���ڶnTzЉ���#�_S����8�(��V[�'���4���GRE��w���H��D������V_H��DAY:3�V��S_Y�Œ~;�SUMMAR���2 $CON?FIG_SEȃ����ʅ_RUN�m�C|�С�$CMPR��P�DEV���_�I�ZP�*��q��ENHANCE�	�
���1���'INT��qM)b�q��2K����OVR6o�PGu�IX��;���OVCT�����v�
 4 ����a�>���PSLG"�� \ �;���?�1���SƁϕc�U�����Ò�4��U�q]�Tp�� (`�-��rJ<�Oz� CK�IL_MJ�b��VN�+��TQn�{�N5���C�UL�ȀD�V(�C6�P_h�຀@�MW�V1V��V1d�2s�2d�3*s�3d�4s�4d���'�	�������p	�I=N	VIB1qp1�B 2!pq/,3 3,4 4,�p?� �;��A���N��������PL��TOR�r3�	��[�SA�V��d�M�C_FOLD 	$SL���Պ�M,�I��L� ��pL�b��KEEP_HNADD	�!Ke�UCCOMc�k��
�lOP���pl��.lREM�k��P΢���U��ek�HPW� KS�BM��ŠCOLL�AB|�Ӱn��n��+�IT�O��${NOL�FCALX� �DON�rZ���o ,��FL�>��$SYNy,�M�C=����UP�_DLY�qs"DGELA� ����Y(��AD��$TAB�TP_R�#�Q�SKIPj% ����OR� �E�� P_��� �)���p 7��%9��%9A�$:N� $:[�$:h�$:u�$:���$:9�q�RA��� X�����MB>�NFLIC]��0�"�U!�o���NO_�H� �\�< _SW�ITCHk�RA_�PARAMG�� ��p��U��W�J��:Cӣ�NGRLT� OO�U�����8X�<A��T_Ja1F��rAPS�WEIG=H]�J4CH�aDcOR��aD��OO���)�2�_FJװ���sA0�AV��C�HOB.�.��l�J2�0�q$�EeX��T$�'QIT���'Q�pG'Q-�GߐR�DC�m" � ��<��
R]��
H�<��RGEA��4��U�FLG`g��H���ER	�SPC�6R�rUM_'P��2�TH2No��@Q 1  ��0�����  D q�وIi�2_P�2�5cS�ᰁ+�L10_CI��pe� �pk����U ՖD��zaxT�p�Q(�;a��c��޲+��i���e��` P>`DESIGRb$�VL1:i1Gf�c�g;10�_DS��D��wp
`FPOS11�q l�pr��xL1C/#AT�B��9U
WusIND��}��mqCp�mq`B	�HO�ME�r `aBq2GrM_q���S 	a�q3Gr�@�� ��$��w4GrG�Y�k�}�����6�5Grď֏�����6�6GrA�S�e��w����� �?t7Gr��П�����`!@s8Gr;�M�_��q�������S �q ` �@sM��P���<K@��! T`M�L�M�IO��m�I��:2�OK _OPy���� »Q�2�pWEG" 7�x EQA�E � #s%Ȳ$wDSBo�GNA�b�� C�P2�_aSw232S�$ �iPr��xc�ICE<@�%�PE`2� @IT���P�OPB7 1�F7LOW�TRa@2��U$�CUN��`�A�UXT��2Ѷ�ER�FAC3İUU�w�,�SCH��'% t<_9�E���A$FREEF'ROMЦ�A�PX q�UPD"YbA�3PT.�pEEX0����!�FA%bҲ���RV�aG� &�  ��E�" 1�AL�  �+�jc�'��D�  2& ��S\PcP(
 ' �$7P�%�R�24� ��T�`AXU���DSP���@�W���:`$��RNP�%�@��z��K��_MIR������MT��AP����P"�qD�QSY�z������QPG7�B�RKH���ƅ AXI�  ^��i�����1 ����BSO�C���N��DUM�MY16�1$S�V�DE��I�FS�PD_OVR7d9� D����OR��֠N"`��F_����@�OV��SF�RU�N��"F0�����U�F"@G�TOd�LC�H�"�%RECOV��9@�@W�`&�ӂ�H��:`_0�  }@�RTINVE��.8AOFS��CK�KbFWD������1B,��TR�a�B �FD� ��1= B1pBL� �6� A1L�V��Kb����#��@+<�AM:��0��j��_M@ ~�@h���T$X`x ��T$HBK���F���A�����PPA�
��	����~��DVC_DB�3�@pA�A"��X1`�X3`��S�@��`�0��Uꣳ�h�CABPP
R�S #���c�B�@���GUBCPU�"��S�P�` R��11)ARŲ�!?$HW_CGpl�11� F&A1Ԡ@8p��$UNITr�|l e ATTRIr@�y"��CYC5B�C�A��FLTR_2_FI������z2bP��CHK_���SCT��F_e'F1_o,�"�*FS�Jj"CHA�Q�'91Is�82RSD����1���_Tg�`�L i�EM�NPMf�T&2 8p&2- �6�DIAGpERAI�LACNTBMw�L�O@�Q��7��PSı�� � ��PRRBSZ`�`BC4�&�	��FUN5s��RIN�PZaߠ�0�7Dh�RAH@���`�� `C�@�`C�Q�C�BLCURuH�DA0�K�!�H�HDAp�aA�H�C�ELD�������C��jA�1�CTI�BUu�8p$CE�_RIA�QJ�AF� P��>S�`DUT�2�0C��};OI<0DF_LC�H���k�LMLF�aH�RDYO���RG��@HZ0��ߠ�@�UM�ULSE�P�'3.iB$J��J�����FAN_ALM��dbWRNeHA#RD��ƽ�P��k@!2aN�r�J�_}��AUJ R+4�TO_SBR��~b�Іj�e 6?A�cMPIN�F��{!�d�A�cREG�NV��ɣZ�5D��NFLW%6r$M�@� ��f� ��0 h'uCM4NF�!�ON	 e!e�#�(b*r3F�3��h	 ���q)5�$�g$Y�r��u�|_��p*$ �/��EG������qAR��i���2�3�u�@<�wAXE��ROB��7RED��WR��c�_���SY`��q� :?�SI�WRI���vE STհ�ӭ d���%Eg!��t8��^a"��B����9�3� �OTO�a���ARY��ǂ�1�����FIE���$LI�NK�QGTH���T_������390���XYZ����!*�OFF������ˀB��,B`l���e���m�FI� ���C@Iû�,B��_J$�F�����S`����3-!$1�w0��d�R��C��,�DU��r��3�P�3TUR`!XS.�Ձ�bXX�� ݗFL�d���pL��0���34���� +1)�K��M��5�5%B'��ORQ�6��fC㘴��0B�O;�D�,������aN�OVE��rM�� ���s2��s2��r1���`0���0�g /�AN=! �2�DQ�q���q�} R�*��6����s��V����ER��jA	�2E���.�C��A���0���XE�2Ӈ�A��AAX��F��A�N!�S� �1_��Q_Ɇ�^ʬ�^� ��^��0^ʙ�^ʷ�^�1&�^ƒP[ɒPkɒP {ɒP�ɒP�ɒP�ɒP �ɒP�ɒP�����ɪ ��R>�DEBU=#�$8ADc�2����
�A!B�7����V� <" 
��i�q��-! ��%��׆��׬��״� ���1�י��׷�JT���DR�m�LAB��8ݥ9 FGRO� ݒ=l� B_�1�u� ��}��`����ޥ��qa��AND�����qa� �Eq��`1��A@�� �NT$`��c�VEL�1��m���1u���QP��m�NA[w�(�CN1� ��3�줙� �SERsVEc�p+ $@@�d@��!��PO�
�� _�0T !���򗱬p, w $TRQ�b�
(� -DR2�,+"P�0_ .� l"@!�&ERR���"I� q���~TOQ����L�p]�e����0G��%��� � RE�@ /� ,��/I -��R�A� 2. d��&�"  0��p$&��2tPM���OC�A8 1 � pCOUNT����FZN_CFG2 4B �f�"T�:#��Ӝ� ��^�s3 ���M:0�R�qC@��/�:0�FA1P��?V�X�����r����� �P:b�pHE�Lpe4 }5��B_BAS�c�RSR�f @�SH�!QY 1�Y 2|*U3|*4|*5|*6|*e7|*8�L!RO�����NL�q �AqB���0Z ACK��[INT_uUS`8�Pta9_PU�>b%ROU��PH@�h9#�u`w�9�TPFWD_KAR��ar RE���PP��A]@QUE�i&��	�f�>`QaI`��9#�j38r��f�SEME��6t��PA�STY43SO�0�DI'1�`p���18�rQ_TM�c�MANRQXF�E�ND�$KEY?SWITCHj31�:A�4HE	�BEA�TM�3PE�pLEP��1��HU~3F�4�2S?DDO_HOeMBPO:a0EF���PRr��*�v�uC��@O�Qo �OV_�Mϒ��Eq�OCM����7��p8%HK��q5 D��g�U�j�2M�p�4R��FwORC�cWAR�����:#OM�p G6 @�Ԣ�v`U|�EP�p1�V'p�T3�VM4�� �p#O�0�L�R7��hUNLiOE0hdEDVaq �Q�@d8 <p�AQ9�l1MSUP�G�UaCALC_�PLANcc1��A�YS1�@�9 � X`��P �q�;a�թ�w��2��j�M�$P�㣒�fyt$��rSC�M�pm�q ���aPq��0�tYzZzCEU�Q�b�� T!��Hr�pPv��NP�X_ASf: 0�g ADD��$�SIZ%a$VA���MULTIP��"��pq�PA�Q; � $T9op�B$���rS��j!C~ �vOFRIF�2S�0��YT�pNF[DODBUX�B��u&�!���#CMtA�Е���x������ 	�SZ >��< � �p��TEg�����$SG%L��T��X�&{��x�㰀��STMTe��ЃPSEG�2��ByW���SHOW؅n�1BAN�`TPO�@��gᣥ������ mV�_G�= ���$PC���O�F�B�QP\�SP�0A�&0^�, VDG���>� �cA00�����P���P���P����P��5��6��7*��8��9��A��b`����P��w᧖S`��F����h���1��v�h��י1�1�1��1��1�1%�12�1�?�1L�1Y�1f�2���2��2��2ʙ2�י2�2�2��2��2�2%�22�2�?�2L�2Y�2f�3���3��3��3ʙ3
י3�3�����U3�3%�32�3߹U3L�3Y�3f�4��U4��4��4ʙ4יU4�4�4��4�U4�4%�42�4߹U4L�4Y�4f�5��U5��5��5ʙ5יU5�5�5��5�U5�5%�52�5߹U5L�5Y�5f�6��U6��6��6ʙ6יU6��6�6��6�U6(�6%�62�6߹U6L�6Y�6f�7��U7��7��7ʙ7יU7��7�7��7�U7(�7%�72�7߹�7L�7Y�7f��V��`_UPD��? ��c 
�V����@ x $gTOR�1T�  �caOP �, ZQ_7�RE^��� J��S�sC�A��_Ux�p��RYSLOA"A � �u$�v���w�@���@��bVALUv10�6�=F�ID_L[C:�HI5I�R$FI�LE_X3eu4$��C��SAV��B� hM �E_BL�CK�3�ȁ�D_CPU��p��p5�hz��@S2R C � PW���� 	�!LAށS�R�#.!'$RUN�`G@%$D!'$�@G%e!$e!'%HR03$� �'$��T2Pa_LI��RD  � G�_O�2�0P_E�DI�R@�T2SPD�#E�"i0ȁ|�p	�
�DCS9@�G)F � 
�$JPC71q�� S�:C;C9$M�DL7$5P>9T�C�`@7UF�@?8S� ?8COBu �@�#T|�L�G�P;;԰ 9:;TAOBUI_�!L�HGb��% FB3�G$�3A�sR�LL�B_AVAI�B �� �2�!��I $n� SEL� NẼ.�@RG_D N��Ta��>ESC�PJS �1/AB�PT�R�	�2_M]`L�Kc \M f/QL_�R�FMj��PGi�U9R��6��PS_�P�\� �p�EE7B�TwBC2�eL ����``�`b$�!FT��P'T�`TDC�g�� BPLp�sNU;WT�H��qhTgtWR��2$�pERVE�.S�T;S�Tw�R_A�CkP MX -$�Q�`.S�T;S�P�U@�`IC�`LOW&�GF1�QR2g�`��p�S�ERTI�A�d^0iP�PEkD�EUe�LACEM&zCC#c�V�BrppTf�edg�aTCV�l�adgTRQ�l�e�j@|�Scu��edcu�J7�_ 4J!��Se@qde�Q2�0���1��PRcuPJKlvVK@<�~qcQ~qw�spJ0�l�q�sJJ�sJJ�sAAL�s�p�s�p�vd���r5sS�`N1�l �p�k�`5dXA_́9A��1BCCF�BN =`M GROU ���bh�NPC0sD�R�EQUIR�R� E�BU�C�Q�6g0 �2Mz��Pd�QS�GUO�@�)AP�PR0C7@� 
$:� N��CLO� ǉ�S^U܉Se
Q�@A.�"P �$PM]P�`8�`sR�_MGa!��C���+��0�@,�B{RK*�NOLD*�SHORTMO�!Hm�Z��JWA�SP�t p`�sp`�sp`�sp`�s(p`�A��7��8sQ!|�QTQ� m���R.Q�cQ�PATH�*� �*��X&����P�NT|@A��"p��� �IN�RU�C4`a��C�`UM��Y
`�)p��>��Q��cP���p��PA�YLOAh�J2LN& R_Am@�L ������+�R_F�2LSHR�T/�L�O���0���>���ACRL0z�p�y�ޤsR9H5b$H+����FLEX��� BJVR P��_._��_�_� BJ�US�0:�_�Vd`0�G��_`tQd`�_�_lF1G� �ũ�o0oBoTofoxo��E�o�o�o�o�o�o �o ����wz3lt�����3EWF�^zT!��X�'qju�� uu~�W؁���p�u �u�u�u������(�T �P5�G�Y��' AT��l�pE�L0�_B��s�J�Svz�JEW�CTR7B�`NA��d�HAN/D_VB�����TUO@`+�`T�SW��V� $$M��e G��AV�Qs�De�oA@A��@�	$�A5�G�AU�Ad�� 6�T�G�DU�Dd�PD�G/ -STI�5V�5Ng�DYF ��+� x����P&�G�&�A�@�lw�o�Q�k�P�� ����ʕӕܕ�RJUW 7 ��� ��3%�?!AS�YMT�(�m�T�Vp*�o�A�t�_SH� ~������$����Ưد�J񬢐�#39\"���_VI��`8|�q0V_UNIrS�4��.�Jmu�2��2 A��4X��4�6a�pt� ������&E_��������E��CH( X� ̱���T-Oc�PP�VsSvD�US�RU�P�����z@�D�A}@_5�U��P�EyAa��RPROG�_NA��$�$�LAST���CA�Ns�ISz@XYZ_SPu�DW]R@Ͱb,VSV@�E1QENc���DCUR�H�Tޜ�HR_T��Y�tQ9S�d��OƓT  �uP?�Z) ��I�!A�D�� �Q���#�S���� �3��vP [ � ME�O��R#B�!T�PPT0F@1�a-�1�̰� h1a�%iT0� $�DUMMY1��o$PS_��RF���% $lfװFL�A*�YP�bc?$GLB_TI �Up�e`ձ#�LIF(!�\����g`OW��P��eVOL#qLb �a_2��[d2[`����b�P�cZ`T�C��$BAUD,v��cST��B�2g`�ARITY0sD_[WAItAIyCJ�2�OU6�ZqyyT�LANS�`�{S�SyZc��BUF_�r��fиx�PyyCHK]_�@CES��� +JO`E�aA�x�bUBYT���� �r�.�.� ��aA���M�������Q] �Xʰ����ST����SBR@M21�_@��T$SV_cER�b����CL�`ʐ�A1�O�BpPGL�h0EW(!^ 4 �$a$Uq$�q$W�9�A��@R��"ՁUم_� "��D$GI���}$ف q^҄�(!` L�\.��"}$F�"E6��NEAR��B$�F}��TQ" J��@R� a7�?$JOINTa�)�y:�ՁMSET(!b  +�Ec�2�^��Se�Ĕ^�(!c�k  ��U�?���LOCK_FO@�� �PBGLV��GmL'�TE�@XM��N�EMP��:�K��b�$U�؂a�#2_���q�`<� 4�q�^��CE/�?���� $KARb�M>�STPDRA܀�����VECX�����I�Uq�av�HE�T�OOL���V��R�EǠIS3��6L��ACH̐m b^Q�ONe[d3���I�dB�`@$RAIL__BOXEa���gROB�@D�?���?HOWWAR0Aa�<i`-�ROLMtb���$�*���T��`����O�_FU�!��HTML58QS�� �&Հ�(!d��& �@��(!e���������B Ӄ}p(!f 	t��m�^a��t��VB�PO��AIPE�N���O����q�|�AORDED��m �z�XT`��A)�RPMO�P go D �`OB� ����ǯ�Uc�`��� ��SYS��ADR���pP`U@^  hs ,"��f$A���E��E��pPV�WVA�Qi �c �@ق�UPR�B>�$EDI�Ad�_VSHWRU�z�ƀ�IS�Uq�pND��P7���G�HEAD��! @���!i�KE�UqO`CP)P��JM�P��L�U;�RAC�E�Tj���IjL�S��C��NE�<����TICK!eMKQ:���HNr��k @���HWC���P�FF��`STYleB+�LO�aD�[�C�l3�
�@�F%�$A��D=��S�!$�1�p a�e�q�e9Pv �FSQU��#�LO�b_1TERC�`"�TS?�m 5���R�m@3����ܡ�O`	c IZ�d�A�eha�qtb}��hA}pP~r��_DO��B�X�pSSQ�SAXI�q��v�bS�U�@TL���REQ_ܠ��ET���`�CJY%��FY'��Af�\!\d9x�P ��  �R$$nl-�w �����c
��uV
Qh(�A ���dC`�A�� 	�Y��D��pH�E"�	CC�C���/�/�/	4!SSC��` o h5�D1Smడ[`SP�@�AT� 
R��L���XbADDR�s$�Hp� IF�Ch�_2CH���pO����- ��TUk�Ir �p��CUCph�V
��I�Rq�4���c
��
K�
�0]!���P'r \z�D����|,K� P�"CN��*�CƮ��!�TXSCREE��s�Pp@��INA˃<�4�Dp"�����`t T� ���b����O Y6������U4h�RR��������R1�T�QUE��u# �j �qz`Ś��'RSML��U����V�1tPS_��6\� �1�9G\���C��2�@4 2��0O�v�R��&F�AMTN_FL*�`Q��W�~ ��BBL_/�9WB`�Pw ����B5O ��BLE"�Cxg�R"�DRIGHt�RD��!CKGR�B`�ET���G�AWIDTHs���RB��a��r �UI��EYհRx d�ʰ�����`y�BACKЍ��>U���PFO܉�QWLAB�?(��PI��$UR�m�~P��P�PHy1 y 8 $�PCT_��,"�R�PRUpP�s5�C_�RO%!Jt�zV�ȇ�pU�@r�SR ���LUM�S��� ERVJ��SP|��T{ � " �GE�Rh� �¯�LIPAeE��)^g@�lh�lh�ki5ik6ik7ikpP`�Z�x����$u1��p�Q� zQUSR�ل| <z��PU�2�a#2�FOO 2�P�RI*m9�[�@pT�RIPK�m�U�NDO��})� ��Yp��y����0i�����p ~�Rp�qG ��T���-!�rOS2��vR��2�s�CA�����ro�$�1i�UIaCA���p�3Ib_�sOFFA�*D@���Ob�r�a5�L�t��GU���Ps��������+QS�UBo� ��E_�EXE��VeуsW]O� �#��wF��WAl�p΁fP=
 V_DB��NRSRT�pO�V☖����3OR/�5�RAU@6�TK���y__���� |j ��OWNj�34$GSRC�0`���DA�<��_MPFI����ESP��T�$0�� c��g��Pp�z�E!G� `%�ۂ34J�n��COP��$���p_���/�+�6���CT�Cہ�ہ�X��DCS��P�4�COMp�@�;��Oo�=��b�K�^�/�VT�qU'���Y٤Z���2���@p�w#SB�����2�\0˰_��M8��%!]�DIC#��sAY�3G�PEE�@T�QS�VR1���eQL�� a��P�D  ��f�z��f�> ����6�9!A�t�b# �~L2SHADOW���#ʱ_UNSCA�d�׳OWD�˰DG�DE#LEGAC�)�q'�VC\ C>��� v����だm�RF07���7�d`C2`7�DRIVo���ϠC�A]�(��` ���MY_UBY�d?Ĳ��s��1�� $0�����_ఆ����L��BM�A$n�DEY	�EXp@,C�/�MU��X��,���0US����;p_R@"1�0p#�2�G�PACIN*���RG��c�y�:�y��sy�C/�RE�R"!�qsBq�y�D@� L 
!�G�P�"��Tp�	R�pD@�&P�Px1Q���	.���RE��SMWq�_Ar�u@+�{�Oq�AA/�3�h�EZ�U���� ��p�HK���P�J��_/�Q0{�EA�N��ۀ2�2�0�MwRCVCA� �:`GORG��Q�dR	��8L�����REFoG�� ���!�+`	�p��������<���q�_ ����r��� S�`C���Ú�W��@D� ���0�!��#q�š�O�U����?� ��Վ2�J@0� 1�*p����0 �UL�@��CO̷0)��� NT �[i�Z�Qf�af% L飏��Q���a�VIAچ�� �ÀHD7 6P�$JO�`oB��$Z_UPo��2Z_LOW��$�QxiBn��1$EP �s�y�� 1!f � � 1¦4� m5�PA�A �oCACHG�LO�w�В�1B���CJn�I#F^��Tm�����$HO2�32{��Uÿ2O�@����Ro��=a��ƐVPx��X@A"_SIZG�K$Z$�F(�G'���C�MPk*FAIo�G���AD�)/�McRE���"P'GP�0�е�9�ASYNB;UFǧRTD�%�$�P!�COLE_2D�_4�5W�sw�~�U�ӍQO��%ECCU��VEM��v]2�VIRC�!5�#�2�!_>�*&�pWp���AG	9R�XYZ@�3�W���8��4d+Qz0T"��IM�1�6�2P�GRABqB�q��;�LERD�9C ;�F_D��F��f50MH�PE�R_�[���l�JRLAqS�@��[_GEb� �H൑~23�E�T����"���b��I��D�ҙ6m�BG_L3EVnQ{�PK|Л6,\q��GI�@N\P4�A��P��!g�dr��S� �NRTZLʁc�Ų��#a��c"!D�qDE����Xа�X���Җ1��
d��pzZ���d�c���D4q��̫��2pT��U&��[ $�ITPr9pp[Q��ՓV�VSF$�d�  fp/�fгUR��ZSMZu9�dr��ADJ`C�v� ZDVf� D�X�AL� � 4 P�ERIKB$MS7G_Q3$Q!o%[���p'��dr:g�qxQ� �XVR\t���B�pT_\��R
_�ZABC"�����Sr���
W��aAC�TVS' � �� $|u�0�cCgTIV�Q!IOu�s&D�IT�x�D�Vϐ
x�P��4�!���pPS����� �#��!���q!L�STD�!�  �_�ST��a�aq�CHx�� L-�@��u��Ɛ*���P GN�A#�C�!q�_F�UN�� ���7ZIPu��HR��$L���XZMPCF"��`bƀ�r�X�ف��LNK��
�Ł�0#�� �$ !��ބCMCMk�C8�C"�����P{q $J8�2�D6!>�O�H�i��T�i�2�����M���U9X�1݅UXE1Ѡ� �1C���Y���������˗7�FTFG>���n��_�Z���X��j��l�Ā��YD�'@ � 8n�R�� Uӱ$HEI3GHd�:h?(! 'v��T���� �c Gd��qp$B% x� E��SHIF��hRVn�F�`�HpC� 3�(�8H`O� ѡ�C��+%D	�"��CE�pV�19���P�HERs� � �,! M�c�u�
�$�POWERFL S �p|����|��p�RG�`  ������_�A�  ��?�p����pd��NSb �����?�  Bz|� �l�  <@�|��%���˃���8�ŵ�� 2ӷ��� 	H��l&����>���A� |��t$���*��/�� **:@���p�ϥ��͘���F������ɘ�� |�����5������� %ߟ�I�[߉�ߑ�� ����������w�!�3� a�W�i��������� ��O����9�/�A��� e�w�������'���� �=O}s �������k 'UK]��� ���C/��-/#/ 5/�/Y/k/�/�/�/? �/�/?�/?�?1?C? q?g?y?�?�?�?�?�? �?_O	OOIO?OQO�� 	 �O�O�O_ �E��3_���O`_�O�_��_÷PREF �Ӻ�p�p
��I?ORITY 4�|�d���p����pSPL`z����WUT�VqÈ�gODU~����Y�_?�OG��Gx���R��,fHIBqO�y�|kTOENT �1��yP(!A�F_t�`�o�g!�tcp�o}!�ud�o)~!�icm�0bXY�̳�k �|�)�� �����p� ���u����� �N�5�r�Y��������̏�����*/c̳�ӹ���E�W�|�>�+^�F��/��4����|��,�7�A��_,  ��P�����%�|�'���Z@��h�z�����|���ENHANCE S	#�7�A9�d��<���  �,f�T�
�_�S����POSRTe�rb�@�U���_CARTR�EP�Pr|brSKS�TAg�kSLGS6�`�k����@�Unothing������Ϳ>��P�b�To��TEMPG ?isϨE/��_a_seibanm_��i_�����0� �T�?�x�cߜ߇ߙ� �߽�������>�)� N�t�_������� ������:�%�^�I� ��m�����������  ��$H3lWi ������� D/hS�w���uϪ�VERS�I�P=g  disable���SAVE �?j	2670H�705��k/!`�m//*�/ 	�(H%b�O�+�/�Se? 6?H?Z?l?z:%<�/�?4�*'_j` 1
�kX �0ubuE�?xOqG�PURGE��1Bp`�ncqWF<@�a�TӒ*fW�`]Daa��WRUP_DELAY z�f�B_HOT %?e�'b��OnER_NORMAL�HGb�O%_�GSEMI_*_i_��QQSKIP�3.��3x��_��_�_ �_�]?eo+goKo]o oo5o�o�o�o�o�o�o �o�o5GYi �}������ �1�C�U��y�g��� ������я����-��?�7%�$RACF�G �[ќ�3��]�_PARAMr�Q3y��S @И�@`�G�42Cj۠��2��CbFzB�B]�BTIF����J]�CVTMOUړ����]�DC�R�3�Y ���Q>�g�@���B�@��jx��S��{�����5�C����0�_��\�� ;e�m����KZ;�=g;�?4�<<���f@8����� �5� G�Y�k�}�������ſ�׿���xURDIO_TYPE  �V��5��EDPRO�T_a�&,>��4BHbCEސS�v�Q2c� ��B�ꐪϸ���ϐ� ���&�ݹ�W�V_~� o����߱������� ��A�O�m�r���9� ������������� �=�_�d������� ����������'I� Nm����� ����#EJi +k����� �//4/F//g// �/y/�/�/�/�/�/	? +/0?O/?c?Q?�?u? �?�?�?�?�??;?,O���S�INT 2��I���l�G;� �jO|K��鯤O�f�0 �O�K�?�O�?_ __N_<_r_X_�_�_ �_�_�_�_�_�_&oo Jo8ono�ofo�o�o�o �o�o�o�o"F4 j|b����������B�O�EFPOS1 1"�?  xO�� o×O����ݏ鈃��� Ϗ0��T��x���� 7���ҟm�������� >�P����7������� W��{�����:�կ ^����������S�e� �� ��$Ͽ�H��l� �iϢ�=���a��υ� � ߻����h�Sߌ� '߰�K���o���
�� .���R���v��#�5� o����������<� ��9�r����1���U� ����������8#\ ����?��u ��"�FX� ?���_��/ �	/B/�f//�/%/ �/�/[/m/�/?�/,? �/P?�/t??q?�?E? �?i?�?�?O(O�?�? OpO[O�O/O�OSO�O wO�O_�O6_�OZ_�O ~_�_+_=_w_�_�_�_ �_ o�_Do�_Aozocf�2 1r�o.o ho�o�o
o.�oR �oO�#�G�k �����N�9�r� ���1���U������� ���8�ӏ\���	�� U�����ڟu�����"� ���X��|����;� į_�q������	�B� ݯf����%�����[� ��ϣ�,�ǿٿ� %φ�qϪ�E���i��� ����(���L���p�� ��/�A�Sߍ������ ��6���Z���W��+� ��O���s������ ��V�A�z����9��� ]���������@�� d��#]��� }�*�'`� ��C�gy� �&//J/�n/	/�/ -/�/�/c/�/�/?�/ 4?�/�/�/-?�?y?�? M?�?q?�?�?�?0O�?�TO�?xOO�O�o�d3 1�oIO[O�O_ �O7_=O[_�O__|_ �_P_�_t_�_�_!o�_ �_�_o{ofo�o:o�o ^o�o�o�o�oA�o e �$6H�� ���+��O��L� �� ���D�͏h�񏌏 �����K�6�o�
��� .���R���퟈���� 5�ПY�����R��� ��ׯr��������� U��y����8���\� n�������?�ڿc� ����"τϽ�X���|� ߠ�)�������"߃� nߧ�B���f��ߊ��� %���I���m���,� >�P���������3� ��W���T���(���L� ��p�����������S >w�6�Z� ���=�a�  Z���z/ �'/�$/]/��//�/@/�/�O�D4 1�Ov/�/�/@?+?d? j/�?#?�?G?�?�?}? O�?*O�?NO�?�?O GO�O�O�OgO�O�O_ �O_J_�On_	_�_-_ �_Q_c_u_�_o�_4o �_Xo�_|ooyo�oMo �oqo�o�o�o�o�o xc�7�[� ���>��b�� ��!�3�E����ˏ� ��(�ÏL��I���� ��A�ʟe������ �H�3�l����+��� O���ꯅ����2�ͯ V����O�����Կ o�����Ϸ��R�� v�Ϛ�5Ͼ�Y�k�}� ����<���`��τ� ߁ߺ�U���y��� &���������k�� ?���c������"��� F���j����)�;�M� ��������0��T ��Q�%�I�mx��/�$5 1�/ ���mX��� P�t�/�3/� W/�{//(/:/t/�/ �/�/�/?�/A?�/>? w??�?6?�?Z?�?~? �?�?�?=O(OaO�?�O  O�ODO�O�OzO_�O '_�OK_�O�O
_D_�_ �_�_d_�_�_o�_o Go�_koo�o*o�oNo `oro�o�o1�oU �oyv�J�n �������u� `���4���X��|�ޏ ���;�֏_������ 0�B�|�ݟȟ���%� ��I��F�����>� ǯb�믆������E� 0�i����(���L��� 翂�Ϧ�/�ʿS��  ��LϭϘ���l��� ��ߴ��O���s�� ��2߻�V�h�zߴ��  �9���]��߁��~� ��R���v����#�	6 1&���� �����������}� ��<��`��� �CUg��& �J�n	k�? �c��/��� 	/j/U/�/)/�/M/�/ q/�/?�/0?�/T?�/ x??%?7?q?�?�?�? �?O�?>O�?;OtOO �O3O�OWO�O{O�O�O �O:_%_^_�O�__�_ A_�_�_w_ o�_$o�_ Ho�_�_oAo�o�o�o ao�o�o�oD�o h�'�K]o �
��.��R��v� �s���G�Џk�􏏏 ���ŏ׏�r�]��� 1���U�ޟy�۟��� 8�ӟ\������-�?� y�گů����"���F� �C�|����;�Ŀ_� 迃������B�-�f� ϊ�%Ϯ�Iϫ���πߣ�,���P�6�H�7 1S����I��� ��������3���0� i���(��L���p� �����/��S���w� ���6�����l����� ��=������6� ��V�z�  9�]���@ Rd���#/�G/ �k//h/�/</�/`/ �/�/?�/�/�/?g? R?�?&?�?J?�?n?�? 	O�?-O�?QO�?uOO "O4OnO�O�O�O�O_ �O;_�O8_q__�_0_ �_T_�_x_�_�_�_7o "o[o�_oo�o>o�o �oto�o�o!�oE�o �o>���^� ����A��e� � ��$���H�Z�l���� �+�ƏO��s��p� ��D�͟h�񟌟��� ԟ�o�Z���.��� R�ۯv�د���5�Я�Y���}�c�u�8 1��*�<�v���߿� �<�׿`���]ϖ�1� ��U���y�ߝϯ��� ��\�G߀�ߤ�?��� c����ߙ�"��F��� j���)�c������ �����0���-�f�� ��%���I���m���� ��,P��t� 3��i��� :���3�� S�w /��6/� Z/�~//�/=/O/a/ �/�/�/ ?�/D?�/h? ?e?�?9?�?]?�?�? 
O�?�?�?OdOOO�O #O�OGO�OkO�O_�O *_�ON_�Or___1_ k_�_�_�_�_o�_8o �_5ono	o�o-o�oQo �ouo�o�o�o4X �o|�;��q ����B���� ;�������[���� ���>�ُb�����!��������MASK +1 �������~ΗXNO  ݟ����MOTE  ����S�_CFG !Z���N�����PL_RANGV��N������OWER� "��Ϡ��S�M_DRYPRG7 %���%W���եTART #�Ǯ�UME_PR�O���q���_EX�EC_ENB  y����GSPDJ�쌰����TDB̯���RMп��IA_OPTION��և����NGoVERS���`�řI_AIR7PUR�� R�+�\��ÛMT_֐T �X���ΐOBOT�_ISOLC���������u�����N�AME8��H�ĚOB_CATEG��ϣ,��S�[�.�O�RD_NUM ?�Ǩ��H?705  N�����ߺ�ΐPC_TI�MEOUT�� x�ΐS232s�1$���� LT�EACH PEN�DAN��o�������V�T�Ma�intenanc�e ConsN��&�M�"B�P�No Use6�r�8����������̒��NPQO$��Ҋ�"���/CH_LM�Q����	a�,�!UD�1:��.�RՐVA3ILw��粥*�_SR  t� ����5�R_INT7VAL���� ����V_DATA_GRP 2'����� D��P �������	��� ���B0R Tf������ /�/>/,/b/P/�/ t/�/�/�/�/�/?�/ (??L?:?p?^?�?�? �?�?�?�?�?O O"O $O6OlOZO�O~O�O�O �O�O�O_�O2_ _V_ D_z_h_�_�_�_�_�_ �_�_o
o@o.oPovo�do�o��$SAF�_DO_PULS�W�[�S���i�SCA�N�������SC�à( �!����
S�S�
���Ķ�q�q�qN� �L^ p���5���� ��$��+�"�r2M�qX�dM�h�rJ�	t/� @��@������ʋ|��� r �ք��_ @N�T ��'�9�K�X�?T D��X��� ������ɟ۟���� #�5�G�Y�k�}�����x��䅎������Ǧ  "�;G�oR� ���p�"�
�u��D�i���q$q�  � ���uq��\� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z����珈������ ������g�;�D�V� h�z���������������(�Ӣ0�r�i�y� ��$�7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/?r�+?=?O?a? s?�?�?�?�?�?8��? OO'O9OKO]OoO�O ��$�r�O�O�O�O 	__-_?_Q_c_u_�_ �Y�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4@FXj|�c�路 g�������0� B�T�f�x���������ҏ������:�.Ҧ��y�3�	��	123456�78��h!B!�� \��p0����Ο�� ���(�:�@��c� u���������ϯ�� ��)�;�M�_�q��� ��R���ɿۿ���� #�5�G�Y�k�}Ϗϡ� �����ϖ�����1� C�U�g�yߋߝ߯��� ������	��-���Q� c�u��������� ����)�;�M�_�q� ��B���������� %7I[m� �������! 3EWi{��� ����////� S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?D/�?�?�?�?�? OO'O9OKO]OoO�O@�O�O�O�O�O*��� �O	_�E�?5_G_Y_�yCz  A��z_   ��x2�r� }��)�
�W�  	�*�2�O�_�_ o$o"l�#\��_ho zo�o�o�o�o�o�o�o 
.@Rdv� ���Mo���� *�<�N�`�r������� ��̏ޏ����&�8��J��X #P$P�Q�R<�u� k��Q  ������S�P����Q�Qt  ЌPÙ۟�P(� `�,b����]�PFl��$SCR_GRP� 1*!+�!4� � ��,a �U	 v��~������d���%����ɯ���h]���P�D1� D�7n��3��Fl
C�RX-10iA/�L 234567W890�Pd� r���Pd�L ��,aC
1o��������[ ¶~�+fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@�R�d�t�?��H�~����m��ϴ����������,a��1���U��[�G�imXhuP,[�}��P0���B�  BƠߞҷԚ�9A�P��  @1`��暡@����� ?����H����ښ�F?@ F�`A�I� @�m�X��|����� ������������:�0%�7�I�[�B�i��� ��������������- Q<u`��En �ٯ���W�P�"+f@_�5��1`b���x����ͣ�O�,dA����ߒ��Fa�,a ��#!"/4/E-!pZ(f/x/G/ (�P�!(� �/�/�/��/�/?#9b����S7�س�M�ECLVLw  ,a��ݲ��Q@f1L_DE�FAULTn4b1��1`�3HOTSTR�=��2�MIPOWERF�m0pU�5�4WF�DO�6 �5L�E�RVENT 1+�u1u1�3 L!DUM_EIP#?�5H�j!AF_�INE�0SO,d!�FT)O�NIO�O!����O ��O�O!�RPC_MAI�N�O�H��O>_SV�IS_�I�-_�_!OPCUf�_�W�y_�_!TP&�PPU�_<Id�_"o�!
PMON_POROXY#o?Feo�no�R<o8Mf]o�o!�RDM_SRV�o<Ig�o!RȠ�"=Hh�oR!
�PM�o9LiA�!RLSYNC���y8��!R3OS(O��4�6��!
CE�PMTC�OM7�?Fk%���!=	K�CONS��>G�lq�Ώ!K�WA'SRC�o?Fm���;!K�USB�=H�n	�f�!STM�0��;JoU����O֟��c����CICE_�KL ?%K �(%SVCPRG1��G�1���c�N�#G3o�t�6�4����"6�5��į6�6��6�7��6���W�R�	9_�d�3���6� 9���6�a�ܿ6���� 6���,�6�ٯT�6�� |�6�)���6�Q���6� y���^����^�ʿD� ^��l�^�ϔ�^�B� ��^�j���^����^� ��4�^���\�^�
߄� ��2���6��/��� �V��<�'�`�K��� o������������� &J5nY�� ������4 F1jU�y�� ���/�0//T/ ?/x/c/�/�/�/�/�/ �/�/??>?)?P?t?�_?�?
�_DEV �I�MC�:�84���4GRP 2/E�0+��bx 	� 
 ,@�?O�� ODO+OhOOOaO�O�O �O�O�O�O�O__@_ R_9_v_]_�_�_O�_ �_�_o�_*ooNo`o Go�oko�o�o�o�o�o �o&8\�_Q �I������ �4�F�-�j�Q����� ��ď���Ϗ��u B�T�;�x�_������� ҟ����ݟ�,��P� 7�t���m�����ί� 7����(�:�!�^�E� ����{�����ܿÿտ ���6��Z�l�Sϐ� 篅���}������ � �D�+�h�z�aߞ߅� ���߻�������� R��v��o����� �������*��N�`� G���k����������� k�8��\nU �y����� �	F-jQ�� �����// B/T/;/x/_/�/�/�/ �/�/�/?�/,??P?p7?I?�?�3d ��6	t?�?�?�?�?O�?�)O8K%�8O]O����vA"AvE�O�G ~O�O�O�O�O�O
YJO /_rI�O\_J_�_n_�_ �_�_�__o@_�_4o "oXoFo|ojo�o�_o �oo�o�o0T Bx�o��oh�d ���,��P��w� �@�����Ώ��ޏ� �(�j�O������p� ����ʟ��ڟ �B�'� f��Z�H�~�l����� Ư������د�� � V�D�z�h����ſ� ������
��R�@� vϸ���ܿf��Ͼ��� �����Nߐ�uߴ� >ߨߖ��ߺ����� � V�|�M��&��n�� �������.��R��� F���V�|�j������� ���*���B0 Rxf����� ��>,Nt ���d���� //:/|a/s/*/L/ &/�/�/�/�/�/?T/ 9?x/?l?Z?|?~?�? �?�?�?,?OP?�?DO 2OhOVOxOzO�O�OO �O(O�O_
_@_._d_ R_t_�O�O�_ _�_�_ �_oo<o*o`o�_�o �_Po�oLo�o�o�o 8zo_�o(�� ������R7� v �j�X���|����� �*��N�؏B�0� f�T���x�����՟� �������>�,�b�P� ��ȟ���v��ί� ��:�(�^�����į N�����ܿʿ�� � 6�x�]Ϝ�&ϐ�~ϴ� ��������>�d�5�t� �h�Vߌ�z߰ߞ��� ���:���.���>�d� R��v�������� ���*��:�`�N��� �����t������� &6\�����L ������"d I[4|�� ���<!/`�T/ B/d/f/x/�/�/�// �/8/�/,??P?>?`? b?t?�?�/�??�?O �?(OOLO:O\O�?�? �O�?�O�O�O _�O$_ _H_�Oo_�O8_�_4_ �_�_�_�_�_ ob_Go �_ozoho�o�o�o�o �o�o:o^o�oR@ vd����� 6�*��N�<�r�`� �����Ϗ�������� &��J�8�n�����ԏ ^�ȟ��؟ڟ�"�� F���m���6�����į ��ԯ֯��`�E��� �x�f���������п &�L��\���P�>�t� bϘφϼ�����"Ϭ� ߨ�&�L�:�p�^ߔ� �ϻ��τ������ � "�H�6�l�ߓ���\� �����������D� ��k���4��������� ����
L�1C�� ��d�����$ 	H�<*LN` ����� �/ /8/&/H/J/\/�/� �/��/�/�/?�/4? "?D?�/�/�?�/j?�? �?�?�?O�?0Or?WO �? O�OO�O�O�O�O �O_JO/_nO�Ob_P_ �_t_�_�_�_�_"_o F_�_:o(o^oLo�opo �o�o�_�oo�o  6$ZH~�o�� n�j���2� � V��}��F������� ԏ
���.�p�U��� ���v���������П �H�-�l���`�N��� r��������4��D� ޯ8�&�\�J���n��� �˿
��������4� "�X�F�|Ͼ����l� ��������
�0��T� ��{ߺ�D߮ߜ����� �����,�n�S��� ��t��������4� �+������L���p� ���������0���$ 46H~l��� ���� 0 2Dz���j� ���/
/,/�� y/�R/�/�/�/�/�/ �/?Z/??~/?r?? �?�?�?�?�?�?2?O V?�?JO8OnO\O~O�O �O�O
O�O.O�O"__ F_4_j_X_z_�_�O�_ _�_�_�_ooBo0o fo�_�o�oVoxoRo�o �o�o>�oe�o .������� �X=�|�p�^��� ���������0��T� ޏH�6�l�Z���~��� ����,�Ɵ ��D� 2�h�V���Ο���|� �x����
�@�.�d� ����ʯT������п ���<�~�cϢ�,� �τϺϨ�������� V�;�z��n�\ߒ߀� �ߤ���������� ��4�j�X��|���� ���������0� f�T��������z��� ����,b�� ���R���� �j�a�:� ����� /B'/ f�Z/�j/�/~/�/ �/�//�/>/�/2? ? V?D?f?�?z?�?�/�? ?�?
O�?.OORO@O bO�O�?�O�?xO�O�O _�O*__N_�Ou_�_ >_`_:_�_�_�_o�_�&oh_Mo�_�Q�$S�ERV_MAILW  �U�`�rh�OUTPUT�h��P@vdRoV 20f  �`� (a\o�ovdS�AVE�l�iTOP�10 21�i d �_HZl~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�e�uYPscFZN_CFG 2e�c�T�a�e|�?GRP 23��q� ,B   A�Ơ�QD;� B�Ǡ�  B4�S�RB21�fHELL�4ev�`��o��/�>�%RSR>�?�Q���u��� ��ҿ������,��@P�;�t�_Ϙϩ���?�  �¼�P���Ϸͻ��P�L&�'�ސW��2�P�d��g��HK ;15�� ,ߡ� �ߥ���������@� ;�M�_���������������OMM �6��?��FTOV_ENB�d�au��OW_REG_�UI_�tbIMIO/FWDL*�7.�ɥ^��WAIT\�`ِ�����`���d��T�IM������V�A�`����_UNI�T[�*yLCy�T�RY��uv`ME�8���aw�rd ���9� ������<��X�Pڠ6p`?�  ���o+=�`VL�l�fM�ON_ALIAS� ?e.��`he Go������/ )/;/M/�q/�/�/�/ �/d/�/�/??%?�/ I?[?m??�?<?�?�? �?�?�?�?!O3OEOWO O{O�O�O�O�OnO�O �O__/_�OS_e_w_ �_�_F_�_�_�_�_�_ o+o=oOoaoo�o�o �o�o�oxo�o' 9�o]o��>� �����#�5�G� Y�k��������ŏ׏ ������1�C��g� y�����H���ӟ��� 	���-�?�Q�c�u� � ������ϯᯌ��� )�;��L�q������� R�˿ݿ��Ͼ�7� I�[�m��*ϣϵ��� ���ϖ��!�3�E��� i�{ߍߟ߱�\����� ������A�S�e�w� ��4���������� �+�=�O���s����� ����f�����' ��K]o��>� ����#5G Y}����l��$SMON_D�EFPROG �&����� &*SYSTEM*����RECALL ?�}� ( �}�/[/m//�/�/�/  I/�/�/�/?"?4?� �*copy mc�:diocfgs�v.io md:�=>192.16�8.56.1:17447?�?�?�?�*�5K2frs:or�derfil.d�at virt:�\temp\b<36372�?O#O5Ow }-�6*.d�?��=�?�O�O�O�&
x�yzrate 11 VOhOzO__/_�%�G�O�A�O�O�_Ƞ_�_�"8�?�8mpback�O}_o#on5o }/K3dbS@*�_�_�_�o�o�o�$3x�T:\To�`fo@�`o"4� 4�ea�o�o|e ��� �_�_co~o�!�3�Fo �jo��������oW i�o��/�Bӏ��x�������'tp?disc 0k����h�z���/��%t�pconn 0  ����������@�͓ S�e�w���,��� Z��������=�O�j� s���(ϻ�͏`�� 7ϔϦ�9�K�\�﯁� �$�6��J�����ϋ��߯�B_T_400  j�|���1�ğ���� �ߋ���B�T�f�x� 	��-�@��A������ ������������x�	 -@��A������� ������fx	 -@�R�ۿ���� ��̿g�{//0/ C��h����/�/�/ ��X/j/� �/?#?5? H��/�/�/�?�?�?� n?j?|?OO1OD��? �?�?�O�O�OBH���? dOvO__+_>P� t�_�_�_��i_��oo'o7l�$SN�PX_ASG 2�:���Va�� �@DP%y�7o~o  ?�Gf�PARAM ;�Ve`a �	*lkP>TDP>X�d�� ��I`O�FT_KB_CF�G  CS\eFcO�PIN_SIM + Vk�b+=�OYsI`RVNOR�DY_DO  ��eukrQSTP/_DSB~�b��>kSR <Vi� � & TELEO�e�{v>TW`�I`TOP_ON_�ERRxGb�PT�N VeP���D:�RING�_PRM'��rVC�NT_GP 2=tVe�ac`x 	����DP��я����BgV}D�RP 1>�i�`�Vq؏0�B�T� f�x���������ҟ� ����,�>�e�b�t� ��������ί��� +�(�:�L�^�p����� ����ʿ�� ��$� 6�H�Z�l�~ϐϷϴ� ��������� �2�D� V�}�zߌߞ߰����� ����
��C�@�R�d� v���������	� ��*�<�N�`�r��� ������������ &8J\n��� �����"4 [Xj|���� ���!//0/B/T/ f/x/�/�/�/�/�/�/ �/??,?>?P?b?t? �?�?�?�?�?�?�?O��PRG_COU�NT�f�P�)IENBe�+EMUC�dbO_UPD 1?�{T  
ODR�O �O�O�O�O__A_<_ N_`_�_�_�_�_�_�_ �_�_oo&o8oao\o no�o�o�o�o�o�o�o �o94FX�| �������� �0�Y�T�f�x����� ���������1�,� >�P�y�t��������� Ο��	���(�Q�L� ^�p����������ܯ � �)�$�6�H�q�l� ~�������ƿؿ����� �I�D�V�"L_I�NFO 1@�E��@��	 �yϽϨ����ɿ�z��>�3=�n߇�w~�� �@k�?���@i*,�]/H���r��
=q���  ?�` >�@��i� D��C�Ҭ�D�	�1��@�G���Y�p����-@YSDEBU)G:@�@�o�d�I��SP_PASS:E�B?��LOG �A���A  ro�i�v�  �A�o�UD1:\x��}���_MPC�ݐ�Ek�}�A&�� ��AK�SAV B���IA���*�i��1�SVB�TEM_TIME 1C��]�@ 0o��i��#�+��"���MEM�BK  �EA��������X�|�@� V�i��@��������h�9
�� ��@�as ���ϻ���nà@Rdv@�����
Le� //(/:/L/^/p/�/ �/�/�/�/�/�/ ??`$?6?H?Z?��SKV��[�EAj��?�?�?��:o�X]2���?i� �po��
:O. @R�O�O�O}N�o�� ��OBi��?�_&_8_,M2��Y_�_�_�_�_�_o�$ �_�_�o'o9oKo]o oo�o�o�o�o�o�o�o �o#5GYk_?�T1SVGUNS�PD�� '�����p2MODE_LIM D��Ҋt�2�p�qE�݉uA�BUI_DCS H}5���0�G� �D�D��|-�X�>���o*���� 
���e��i���r�i������uEDIT� I��xSCR/N J���rS�G K�.�(�0�߅SK_OPTI�ON��^����_D�I��ENB  ��E���BC2_G_RP 2L������&AMPC�ʓ�|B�CCF/�N���� 1����`�>� W�B�g���x�����կ ��������S�>� w�b���������Ͽ�� ���=�(�a�Lυ� ��Ň�϶�������v� �
�/�U�@�yߧ�� `�iМ��߰�����
� ��.��>�@�R��v� �����������*� �N�<�r�`������� ��������̀4 FX��|j��� ����B0 fTvx���� �/�,//</b/P/ �/t/�/�/�/�/�/�/ �/(??L?d?v?�? �?�?6?�?�?�?O O 6OHOZO(O~OlO�O�O �O�O�O�O�O __D_ 2_h_V_�_z_�_�_�_ �_�_
o�_.oo>o@o Ro�ovo�ob?�o�o�o �o<*Lr` �������� &��6�8�J���n��� ��ȏ���ڏ��"�� F�4�j�X���|����� ���֟��o$�6�T� f�x���������ү�� �����>�,�b�P� ��t��������ο� �(��L�:�\ς�p� �ϔ��ϸ������� � �H�6�l�"��ߖߴ� ����V������2� � V�h�z�H������ ��������
�@�.�d� R���v����������� ��*N<^` r������� &8�\Jl�� ������"// F/4/V/X/j/�/�/�/ �/�/�/?�/?B?0? f?T?�?x?�?�?�?�? �?O�?,O�DOVOtO �O�OO�O�O�O�O�O�_ V4P�$TBC�SG_GRP 2�O U� � �4Q 
 ?�  __q_[_�_ _�_�_�_�_�_o%k�8R?SQF\d��HTa?4Q	 H�A���#e>����>$a�\#eAT��A WR�o�h|djma�G�?Lfgr�bp�o�n�ffhfG��ͼb4P|j��o�*}@��Rhf�ff>�33pa#e<q!B�o+=xrRp�qrUy�rt~��H�y0 rIpTv�pBȺt~ 	xf	x(�;���f����N�`���ˏڋ�����	V3.00~WR	crxlڃ	*��3R~t2��HH��� \�.�n]�  cC.�X����8QJ2?SRF]�����CFG -T UPQ SPܚ+��r�ܟ1��1�W�e�	Pe� ��v�����ӯ����� ���Q�<�u�`��� ������Ϳ�޿�� ;�&�_�Jσ�nπϹ� ��������WRq@� 0�B���u�`߅߫ߖ� �ߺ������)�;�M� �q�\������4Q  _���O ���J�8� n�\������������� ����4"XFh j|������ .TBxf� �nO����// >/,/b/P/�/t/�/�/ �/�/�/�/�/?:?(? ^?p?�?�?N?�?�?�? �?�?�? O6O$OZOHO ~OlO�O�O�O�O�O�O �O __D_2_T_V_h_ �_�_�_�_�_�_
o�_ o@o�Xojo|o&o�o �o�o�o�o�o* N`r�B��� ����&��6�\� J���n�����ȏ��؏ ڏ�"��F�4�j�X� ��|���ğ���֟� ��0��@�B�T���x� ����ү䯎o���̯ ʯP�>�t�b������� �������Կ&�L� :�p�^ϔϦϸ��τ� ����� �"�H�6�l� Zߐ�~ߴߢ������� ���2� �V�D�z�h� ������������� 
�,�.�@�v����� ��\�������< *`N����x ���8J\ (������ ��/4/"/X/F/|/ j/�/�/�/�/�/�/�/ ??B?0?f?T?v?�? �?�?�?�?�?OO�� 2ODO�� O�OtO�O�O �O�O�O_�O(_:_L_ 
__�_p_�_�_�_�_ �_ o�_$oo4o6oHo ~olo�o�o�o�o�o�o �o D2hV� z�����
�� .��R�@�b���v��� &OXO֏菒����� N�<�r�`�������̟ ޟ🮟��$�&�8� n�������^�ȯ��� گ��� �"�4�j�X� ��|�����ֿĿ�� ��0��T�B�x�fψ� �Ϝ����������� >�P���h�zߌ�6߼� �����������:�(� ^�p���R�����8�� ���  &�*�� *�>�*��$�TBJOP_GR�P 2U����  ?�/��C*�	V�]��Wd������X  �*��� �,� � ���*�� @&�?��	 ߐA�����C��  DD�����>~v�>\? ���aG�:�o���;ߴAT������A�<��M�X����>��\)�?���8Q�|����L��>�0 ^&�;iG.���Ap< � F�A�ff�v��� ^):VM�.�� �S>o*�@��R�Cр	���������ff�:��6/�?�33�B   ��/�������>):�S���� �/�/@��H�%&/��/��=� <#��
*��v�;/��f�!?���4B�3 ?'?2	��2?hZ?D? R?�?�?�?F?�?�?�? �?OAOO�?`OzOdO�rO�O�O*�C�*����A��	V3.0}0{�crxl��*P��%�%c5Z F� JZ�H F6� F�^ F�� F��f F� G�� G5 G�<
 G^] G�� G���G��*�G�S G��; G��ERD�u�\E[� E�� F( F�-� FU` F�}  F�N F�� F�� F�ͺ F� F��V G� G�z Ga 9'ѷ�Q�LHefJQ4�o,b*�0c�1���OH�ED_TCH Xd�+X2S��&�&�d$�'X�o�o*�1F�T�ESTPARS c ��cV�HRpABLE 1Yd� N`*�����g)$j�g�h�h)�T1��g	�h
�h�hTHu*��h�h�h�%vRDI0n��GYk}��u	�O �#�-�?�Q�c�u�)r	S�l� �z6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ��I���m�Fwͩ�� ȏڏ쏘������x)r��NUM  ���n����2� Ep�)r_CF�G Z��I���@�V�IMEBF_T�TqD��e޶VE�R�����޳R {1[8{ 8�o�*�%�Q� ��د  9�K�]�oρϓϥ� �����������#�5� G�Y�k�}��ߡ߳��� ��������1���E� W�i�{�������� ������/�A�S�e� w���������������@+=O�_����@��`LIF7 \��D`�����DR�(FP
��!p�!p� d�� ��MI_CHA�N� � DB/GLVL��f�ETHERAD S?u��0`1��_}�ROUT6�!�j!��~SNMASKY|�j255.%�S///A/S�`OOLOFS_DIp��CORQCTRL ]8{��1o�-T�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OL�/6O%O�ZOcPE_DET�AI7�*PGL_�CONFIG �c������/c�ell/$CID?$/grp1^O�O �O�O
__|���G_ Y_k_}_�_�_0_�_�_ �_�_oo�_CoUogo yo�o�o,o>o�o�o�o 	-�oQcu� ��:����� )���_�q���������׮}N����%�@7�I�a�KOq�P��M� ����ʟܟ� �G�$� 6�H�Z�l�~������ Ưد������2�D� V�h�z������¿Կ ���
ϙ�.�@�R�d� vψϚ�)Ͼ������� �ߧ�<�N�`�r߄� ��%ߺ��������� &��J�\�n���� 3����������"��� F�X�j�|��������@��User �View �I}}�1234567890����+=�Ex �e����2 ��B������`r��3�Oas@����x4> //'/9/K/]/�~/x5��/�/�/�/�/?p/2?x6�/k?}?��?�?�?�?$?�?x7 Z?O1OCOUOgOyO�?�Ox8O�O�O�O	_�_-_�ON_TR �lCamera���O�_�_�_�_�_�_˂E�_o)o;n���Uogoyo�o�o�o�)  mV�	�_�o#5 GY o}���o�@�����F_�mV =�k�}�������ŏ l����X�1�C�U� g�y���2�D��"�ן �����1�؏U�g� y�ğ������ӯ��� ��D��k��E�W�i�{� ����F�ÿտ�2�� �/�A�S�e��nUY9 ������������	߰� -�?�Qߜ�u߇ߙ߫� ����v�D�If��-� ?�Q�c�u�ߙ��� �������)�;��� D��I����������� ����)t�M_@q���N�`�93 ��0B��S x�1�����(//�J	oU0�U/ g/y/�/�/�/V�/�/ �/�?-???Q?c?u? /./tPv[?�?�?�? OO(O�/LO^OpO�? �O�O�O�O�O�O�?oU �k�O:_L_^_p_�_�_ ;O�_�_�_'_ oo$o 6oHoZo_;%N��_�o �o�o�o�o �_$6 H�ol~���� moe��]�$�6�H� Z�l��������؏ ���� �2��e&� ɏ~�������Ɵ؟� ��� �k�D�V�h�z� ����E�e��5���� � �2�D��h�z��� ׯ��¿Կ���
ϱ�  ��9�K�]� oρϓϥϷ���������   ��5� G�Y�k�}ߏߡ߳��� ��������1�C�U� g�y���������� ��	��-�?�Q�c�u� ���������������);M_q� � 
��(  �>-�( 	 �� �����#3 5G}k����
� �Y�
// ./��R/d/v/�/�/�/ ����/�/�/A/?0? B?T?f?x?�/�?�?�? ?�?�?OO,O>O�? bOtO�O�?�O�O�O�O �O_KO]O:_L_^_�O �_�_�_�_�_�_#_ o o$ok_HoZolo~o�o �o�_�o�o�o1o  2DVh�o�o�� �	��
��.�@� �d�v��������Џ ���M�*�<�N��� r���������̟�%� ��&�m�J�\�n��� �����ȯگ�3�� "�4�F�X�j������� ����ֿ�����0� w���f�xϊ�ѿ���� �������O�,�>�P� ��t߆ߘߪ߼���� ����]�:�L�^�p�p����߻@ ����������� ���"frh:\t�pgl\robo�ts\crx!�1�0ia_l.xml��D�V�h�z�����`�������������� 0BTfx�� �������, >Pbt���� ����/(/:/L/ ^/p/�/�/�/�/�/�/ ��/?$?6?H?Z?l? ~?�?�?�?�?�?�/�? O O2ODOVOhOzO�O �O�O�O�O�?�O
__ ._@_R_d_v_�_�_�_ �_�_�O�_oo*o<o No`oro�o�o�o�o�ot�n �6� ���<< 	� ?��k!�o;i Oq������ ���%�S�9�k����o�����я����(��$TPGL_O�UTPUT f������� �&�8�J�\�n��� ������ȟڟ���� "�4�F�X�j�|�����в�į�p�ր23�45678901 �����1�C�K��� �r���������̿d��п��&�8�J��} T�|ώϠϲ���\�n� ����0�B�T���b� �ߜ߮�����j���� �,�>�P����߆�� �������x����(� :�L�^���l������� ����t���$6H Zlz���� ��� 2DVh  ������ �/./@/R/d/v// �/�/�/�/�/�/�/ۂ? $$��ί <7*?\?N?�?r?�?�? �?�?�?�?OO4O&O XOJO|OnO�O�O�O�O��O�O_�O0_"_T_} �an_�_�_�_�_�_�]�@�_o	z ( 	 V_Do2oho Vo�ozo�o�o�o�o�o 
�o.R@vd �������� �(�*�<�r�`���ܦ��  << I_ˏݏ������� :�L�֪��}���)��� ş�������k��C� ݟ/�y���e������ �������-�?��c� u�ӯ]�����W��� Ϳ��)χ���_�q�� yϧρϓ�����M�� %߿��[�5�Gߑߣ� ߫���s����!��� E�W��?���9��� ������i���A�S� ��w���c�u����/� ����=)s �����U�� �'9�!o	[ �����K�#/ 5/�Y/k/E/w/�/� /�/�/�/�/?�/? U?g?�/�?�?7?�?�?�?�?	OO��)WGL1.XML�_�PM�$TPOFF_LIM ���P����^FN_�SVf@  �T�xJP_MON Mg��zD�P�P�2ZISTRTCHOK h��xFk_�aBVTCOMPA�T�HQ|FVWVA/R i�M:X�D� �O R_�P��BbA_DEFP�ROG %�I�%TELEOP� Pi_VM_DIS�PLAYm@�N�RI�NST_MSK � �\ �ZIN�USER_�TLC�Kl�[QUICK�MEN:o�TSCR�EY`��Rtpsc�Tat`yi4xB�`_�iSTZxI�RACE_CFGW j�I:T�@�	[T
?��hHNL 2k�Z���aA[ gR-?Qcu����z�eITEM� 2l{ �%�$1234567�890 ��  =�<
�0�B�J�  !P�X�dP���[S ���"���X�
�|� ��W���r�֏����.� �0�B�\�f�����6� \�n�ҟ�������� >���"���.����� ίR����Ŀֿ:�� ^�p�9ϔ�Tϸ�xϊ� ��d���H��l� �>�Pߴ�\������� v� ������h�(�� �߰�4�L��ߦ��� ��@�R��v�6���Z� l���������*��� N��� ���������� ��X���J
 n���b�� ��"4F�/| </N/�Z/���// �/0/�/?f/?�/�/ e?�/�?�/�?�?�?,? �?P?b?t?�?�?DOjO |O�?�OOO(O�O�O ^O_0_�O<_�O�O�_ �O�__�_�_H_�_l_(~_Go�dS�bm�oLj��  �rLjq �a�o�Y
 �o��o�o�o{jUD1�:\|��^aR_�GRP 1n�{� 	 @�P Rd{N�r����~��p���q+�x�O�:�?�  j� |�f����������ҏ ����>�,�b�P���`t���������	e����\cSCB 2ohk U�R�d� v���������Я�Rl�UTORIAL �phk�o-�WgV_�CONFIG �qhm�a�o�o��<�O�UTPUT r<hi}�����ܿ � ��$�6�H�Z�l� ~ϐϢϴ�z�ɿ����  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������� �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/��/�/?? 0?B?T?f?x?�?�?�? �?�/�?�?OO,O>O PObOtO�O�O�O�O�? �O�O__(_:_L_^_ p_�_�_�_�_�_f�x� ǿoo,o>oPoboto �o�o�o�o�o�o�O (:L^p�� �����o ��$� 6�H�Z�l�~������� Ə؏��� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я�� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� ���������������X���# ��N�_r���� ���&8J ��n������ ��/"/4/F/X/i |/�/�/�/�/�/�/�/ ??0?B?T?e/x?�? �?�?�?�?�?�?OO ,O>OPOa?tO�O�O�O �O�O�O�O__(_:_ L_^_oO�_�_�_�_�_ �_�_ oo$o6oHoZo k_~o�o�o�o�o�o�o �o 2DVgoz �������
� �.�@�R�d�u���� ����Џ����*� <�N�`�q��������� ̟ޟ���&�8�J��\�k��$TX_S�CREEN 1s�% �}�k�����ӯ���	���Z��I�[�m� ������,�ٿ��� �!�3Ϫ�W�ο{ύ� �ϱ�����L���p�� /�A�S�e�w��� ߭� ���������~�+�� O�a�s���� ��� D�����'�9�K��� �������������R� ��v�#5GYk}�����$UALR�M_MSG ?����� �n�� �	:-^Qc ������ /��SEV  ��2&�ECFG �u����  }n�@�  Ab!�   B�n�
 /u����/�/�/�/ �/�/??%?7?I?W7~>!GRP 2vH+w 0n�	 /��?� I_BBL_NOTE wH*�T��l�u���w�T �2DE�FPRO� %� (%�Ow�	OBO -OfOQO�OuO�O�O�O��O�O_�O,_�<FK�EYDATA 1yx���0p W'n��?�_�_z_�_�_ưZ,(�_on�(�POINT  ]xonc NCEL@o�ko�PNDIREC�Tlono EXT �STEP�omTOUCHU�o�o�P�ORE INFO �o�o0B)fM� ����������>�P� ���/frh/gui�/whiteho?me.pngQ��������ŏ׏�h�pointz���/��A�S��  FRH�/FCGTP/wzcancel���������ʟܟk�i�i?ndirec����'�9�K�]�h�z�nex�������ϯ���h�touchup���/�A�S�e��}h�arwrg�� ����ÿտ�n��� (�:�L�^�p����Ϧ� ��������}��$�6� H�Z�l��ϐߢߴ��� �����ߋ� �2�D�V� h�z�	��������� ����.�@�R�d�v� ��_������������� �2DVhz� �����
� @Rdv��) ����//�</ N/`/r/�/�/%/�/�/ �/�/??&?�/J?\? n?�?�?�?3?�?�?�? �?O"O�?4OXOjO|O �O�O�OAO�O�O�O_ _0_�OT_f_x_�_�_ �_=_�_�_�_oo,o >o�_boto�o�o�o�o�W��k�b�����o}�o8J$v,6�{.��� ������/�� S�:�w���p�����я �ʏ��+��O�a� H���l�������ߟ� ��'�9�Ho]�o��� ������ɯX����� #�5�G�֯k�}����� ��ſT������1� C�U��yϋϝϯ��� ��b���	��-�?�Q� ��u߇ߙ߽߫����� p���)�;�M�_��� ���������l�� �%�7�I�[�m���� ����������z�! 3EWi����� ����П/A Sew~���� ��/�+/=/O/a/ s/�//�/�/�/�/�/ ?�/'?9?K?]?o?�? �?"?�?�?�?�?�?O �?5OGOYOkO}O�OO �O�O�O�O�O__�O C_U_g_y_�_�_,_�_ �_�_�_	oo�_?oQo couo�o�o�o:o�o�o �o)�oM_q ���6������%�7�9��>���b�t� ��^�������,��� �����3�E�,�i�P� ������ß������� ��A�S�:�w�^��� ����ѯ����ܯ�+� 
O�a�s�������� Ϳ߿���'�9�ȿ ]�oρϓϥϷ�F��� �����#�5���Y�k� }ߏߡ߳���T����� ��1�C���g�y�� �����P�����	�� -�?�Q���u������� ����^���); M��q����� �l%7I[ ������h �/!/3/E/W/i/@� �/�/�/�/�/�/�? ?/?A?S?e?w??�? �?�?�?�?�?�?O+O =OOOaOsOO�O�O�O �O�O�O_�O'_9_K_ ]_o_�__�_�_�_�_ �_�_�_#o5oGoYoko }o�oo�o�o�o�o�o �o1CUgy� �����	�� �?�Q�c�u�����(� ��Ϗ������;��M�_�q�������~ ����~ ���ҟ���Ο�*��,�[���f����� ��ٯ�������3�� W�i�P���t���ÿ�� �ο��/�A�(�e� Lωϛ�z/�������� ��(�=�O�a�s߅� �ߩ�8��������� '��K�]�o���� 4����������#�5� ��Y�k�}�������B� ������1��U gy����P� �	-?�cu ����L��/ /)/;/M/�q/�/�/ �/�/�/Z/�/??%? 7?I?�/m??�?�?�? �?�?���?O!O3OEO WO^?{O�O�O�O�O�O �OvO__/_A_S_e_ �O�_�_�_�_�_�_r_ oo+o=oOoaosoo �o�o�o�o�o�o�o '9K]o�o�� ������#�5� G�Y�k�}������ŏ ׏������1�C�U� g�y��������ӟ� ��	���-�?�Q�c�u� �������ϯ������0���0���B�T�f�>�����t�,��˿~�� ֿ�%��I�0�m�� fϣϊ����������� !�3��W�>�{�bߟ� �ߘ��߼�����?/� A�S�e�w���� ����������=�O� a�s�����&������� ����9K]o ���4���� #�GYk}� �0����// 1/�U/g/y/�/�/�/ >/�/�/�/	??-?�/ Q?c?u?�?�?�?�?L? �?�?OO)O;O�?_O qO�O�O�O�OHO�O�O __%_7_I_ �m__ �_�_�_�_�O�_�_o !o3oEoWo�_{o�o�o �o�o�odo�o/ AS�ow���� ��r��+�=�O� a����������͏ߏ n���'�9�K�]�o� ��������ɟ۟�|� �#�5�G�Y�k����� ����ůׯ������ 1�C�U�g�y������ ��ӿ������-�?ϠQ�c�uχ�^P��}�^P�����@���ͮ���
���,�� ;���_�F߃ߕ�|߹� �����������7�I� 0�m�T������� �����!��E�,�i� {�Z_������������ �/ASew� ������ +=Oas�� ����//�9/ K/]/o/�/�/"/�/�/ �/�/�/?�/5?G?Y? k?}?�?�?0?�?�?�? �?OO�?COUOgOyO �O�O,O�O�O�O�O	_ _-_�OQ_c_u_�_�_ �_:_�_�_�_oo)o �_Mo_oqo�o�o�o�o ���o�o%7>o [m����V ���!�3�E��i� {�������ÏR���� ��/�A�S��w��� ������џ`����� +�=�O�ޟs������� ��ͯ߯n���'�9� K�]�쯁�������ɿ ۿj����#�5�G�Y� k����ϡϳ������� x���1�C�U�g��� �ߝ߯����������`�����`���"�4�F��h�z�T�,f���^������ ���)��M�_�F��� j����������� ��7[B�x �����o!3 EWixߍ��� ����///A/S/ e/w//�/�/�/�/�/ �/�/?+?=?O?a?s? �??�?�?�?�?�?O �?'O9OKO]OoO�OO �O�O�O�O�O�O_�O 5_G_Y_k_}_�__�_ �_�_�_�_o�_1oCo Uogoyo�o�o,o�o�o �o�o	�o?Qc u��(���� ��)� M�_�q��� �����ˏݏ��� %�7�Ə[�m������ ��D�ٟ����!�3� W�i�{�������ï R������/�A�Я e�w���������N�� ����+�=�O�޿s� �ϗϩϻ���\���� �'�9�K���o߁ߓ� �߷�����j����#� 5�G�Y���}���� ����f�����1�C�hU�g�>�i��>������������������,�� ?&cu\��� ����)M 4q�j���� �/�%//I/[/:� /�/�/�/�/�/���/ ?!?3?E?W?i?�/�? �?�?�?�?�?v?OO /OAOSOeO�?�O�O�O �O�O�O�O�O_+_=_ O_a_s__�_�_�_�_ �_�_�_o'o9oKo]o oo�oo�o�o�o�o�o �o�o#5GYk} ������� �1�C�U�g�y���� ����ӏ���	���-� ?�Q�c�u�����p/�� ϟ�����;�M� _�q�������6�˯ݯ ���%���I�[�m� �����2�ǿٿ��� �!�3�¿W�i�{ύ� �ϱ�@��������� /߾�S�e�w߉ߛ߭� ��N�������+�=� ��a�s�����J� ������'�9�K��� o�����������X��� ��#5G��k}@����������������&�HZ4, F/�>/����� 	/�-/?/&/c/J/�/ �/�/�/�/�/�/�/? �/;?"?_?q?X?�?|? �?�?���?OO%O7O IOXmOO�O�O�O�O �OhO�O_!_3_E_W_ �O{_�_�_�_�_�_d_ �_oo/oAoSoeo�_ �o�o�o�o�o�oro +=Oa�o�� �������'� 9�K�]�o�������� ɏۏ�|��#�5�G� Y�k�}������şן ������1�C�U�g� y��������ӯ��� 	��?-�?�Q�c�u��� ������Ͽ���� ��;�M�_�qσϕ�$� ���������ߢ�7� I�[�m�ߑߣ�2��� �������!��E�W� i�{���.������� ����/���S�e�w� ������<������� +��Oas�� ��J��' 9�]o���� F���/#/5/G/��$UI_INU�SER  ����h!��  H/L/_M�ENHIST 1�yh%  �(u  �)/�SOFTPART�/GENLINK�?current�=menupag�e,1133,1 �/�/??�'�/�.71�/{?�?�?�?�y+E?�%edit�"?TELEOPj?O O'O�?D?V?2�/�O��O�O�O�(MO�/48,2�O
__._@_<�/�O,163i?�_@�_�_�_Q_c_uR2{_�o"o4oFo�O�_�!5�qO�o�o�o�o��� ��!�a�o�o!3EW �o|��� ��e���0�B� T��x���������ҏ �s���,�>�P�b� 񏆟������Ο��o� ��(�:�L�^�p��� ������ʯܯ��o� $�6�H�Z�l�~����� ��ƿؿ����� �2� D�V�h�z�	Ϟϰ��� ������
ߙ�.�@�R� d�v߈�߬߾����� ����*�<�N�`�r� ���%��������� ����J�\�n����� ������������" ��FXj|��/ ����0� Tfx���=� ��//,/�=/b/ t/�/�/�/�/K/�/�/ ??(?:?%��/p?�? �?�?�?�?�/�? OO $O6OHO�?lO~O�O�O �O�O�OgO�O_ _2_ D_V_�Oz_�_�_�_�_ �_c_�_
oo.o@oRo do�_�o�o�o�o�o�o qo*<N`K;��$UI_PAN�EDATA 1{�����q�  	�} � frh/cgt�p/flexde�v.stm?_w�idth=0&_�height=1�0�p�pice=T�P&_lines�=15&_col�umns=4�pf�ont=24&_�page=who�le�pmI6)  grim�9�  �p P�b�t���������� ��Ǐ��(�:�!�^� E�����{�����ܟ��՟�I6� � �   	 :�J�O�a�s��� ������ͯ@���� '�9�K���o���h��� ��ɿۿ¿���#�5� �Y�@�}Ϗ�vϳ�&��Ɠs�����)� ;�Mߠ�q�䯕ߧ߹� ������V��%��I� 0�m��f������ ������!��E�W��� �ύ�����������:� ~�/ASew� �����  =$asZ�~ ����d�v�'/9/ K/]/o/�/��/�/* �/�/�/?#?5?�/Y? @?}?�?v?�?�?�?�? �?O�?1OCO*OgONO �O�/�/�O�O�O	_ _-_�OQ_�/u_�_�_ �_�_�_6_�_o�_)o oMo_oFo�ojo�o�o �o�o�o�o%7�O �Om���� �^_�!�3�E�W�i� {������Ï����� ����A�S�:�w�^� ������џDV�� +�=�O�a�������
� ��ͯ߯���|�9�  �]�o�V���z���ɿ ���Կ�#�
�G�.�k�ޟ�}�|ϵ����������)��4ߧ� #�`�r߄ߖߨߺ�!� ���������8��\� C���y������������������$U�I_POSTYP�E  ��?� 	 �s��B�QUICKME/N  Q�`�v��D�RESTORE� 1|���  �*default���  INGLE~��PRIM���meditpa�ge,TELEOP,1Sew� ,������� /ASe���z ������/!/ �E/W/i/{/�/0/�/ �/�/�/�/�??*? �/e?w?�?�?�?P?�? �?�?OO+O�?OOaO sO�O�OB?�O�O�O:O __'_9_K_�Oo_�_ �_�_�_Z_�_�_�_o #o�O�_BoTo�_xo�o �o�o�o�o�o1 CU�oy�����{�SCRE��?���u1sc���u2�3�4��5�6�7�8���sTATM�� �����:�USER��p��rT�p�ksT���4��5��6���7��8��B�NDO_CFG }Q�X����B�PDE����None���v�_INFO �2~��)���0%�D���2�s�V��� ����͟ߟ��'� 9��]�o�R���z���OFFSET 	�Q�-���hs��p �����G�>�P�}� t���Я��׿ο�� ��C�:�L�^Ϩ����͘���
����av���WORK �!�����.�@ߢ�u�_UFRAM ����RTOL_A�BRT�����EN�B�ߣ�GRP 1������Cz  A������*�<�N�`�r��֐�U������MSK  ��)���N��%�!��%z����_EVN�����+�ׂ�3�«
 h��UEV��!t�d:\event?_user\�u�#C7z���jpF��n��SPs�x�spo�tweld��!�C6��������! ���G|'��5k Y�����> ���1�Ug ���/��	/^/ M/�/-/?/�/c/�/�/ �/�/$?�/H?�/:J��W�3�����8C?�?�? �?�?�?�? O+OOOOaO<O�O�O rO�O�O�O�O_�O'_ 9__]_o_J_�_�_�_��$VALD_C�PC 2�« ��_�_�  w��qd�R�*o_oqo��
hsNbd�j�`��i �da{�oav�_�ooo 3BoWi{�o�o�o �o��o�PA� 0�e�w������ ����(�=�L�a� s�
�������ʏ��� ��$�ޟH�:�o��� ������ڟ؟�����  �2�G�V�k�}����� ��¯ԯ�����.� �R�S�yϋϚ����� �����	��*�<�Q� `�u߇ߖϨϺ����� ����&�8�M�\�q� ���߶���n����� �"�4�F�[�j���� ������������! 0�B�Wf�{���� �������,> teT����� ��/+/:La/ p�/�/./���� �//'?6/H/?l/^? �?�?�/�/�/�/�/? #O�?D?V?kOz?�O�O �?�?�?�?�?_O1_ @ORO9_vOw_�_�_�O �O�O_�__-o<_N_ `_uo�_�o�o�_�_�_ �_o&o;Jo\oq �o����o�o�o�  �"7�FXj�� ���������!� 0�E�T�f�{������� ßҏ����
�,�A� P�b�����x�����Ο �����(�*�O�^� p���������R�ܯ�  ��Ϳ6�K�Z�l�&� ���Ϸ���ؿ���"�  �2�G���h�zϏߞ� ����������
��1� @�U�d�v�]�ߛ��� �������,��<�Q� `�r���������� ����&�;J�_n� ������������ �$F[j|� ������ 0E/Ti/x��/� �/�/�/�//,/.? P/e?t/�/�/�?�?�? �?�/??(?:?L?NO sO�?�?�O�?�O�OvO  OO$O6O�OZOo_~O �OJ_�O�_�_�_�O_� _F_D_V[�$VA�RS_CONFI�G ��Pxa�  FP�]S�\lCMR_�GRP 2�xk� ha	`�` � %1: SC�130EF2 *H�o�`]T�VU�P�h�`�5_Pa?��  A@%pp*`�NVn No9xC VXdv��a��<u�A�%p�q�_R���_R B���#�_Q'��H�� l�;���{�����؏Ï Տ�e��D�/�A�z��-�����ddIA_W�ORK �xe�ܐ�Pf,		�Qxe���G�P ����YǑRTSY�NCSET  �xi�xa-�WINU�RL ?=�`�����������ȯگ�SIONTMO�U9�]Sd� ���_CFG ��S۳�S۵P��` FR:�\��\DATA\�� �� M�C3�LOG@�  � UD13�EX�d�_Q' B@ ����x�e_ſ�x�ɿ�VW �� n6  ����VV��l�q  =���?�]T<��y�Y�TRAIN؎��N� 
gp?�CȞ��TK���b�xk (g����� _���������U�C� y�g߁ߋߝ߯����߮�_GE��xk�`_P�
�P�R���RE��xe*�`h�LEX�xl`1�-e�VMPHA�SE  xec��ecRTD_FILTER 2�xk �u�0��� �0�B�T�f�x����� VW�������� $�6HZl_iSHI�FTMENU 1��xk
 <�\%�������� ��=&sJ\ �������'/��	LIVE/�SNA�c%vs�fliv��9/���� 7�U�`\"menur/w//�/�/������]��MO���y��5`h`ZD�4�V�_Q<��0���$WAITDIN�END��a2p6OK  �i�<���?�S�?�9TIM�����<Gw?M�?*K��?
J�?
J�?�8RELE��:G6p3���r1_ACTO 9Hܑ��8_<� �ԙ��%�/:_af�BRDI�S�`�N�$XV�R��y��$Z�ABC�b1�S;S ,��j�I�2B_�ZmI1�@VSPT ��y��eG�
�*�/o�*!o7o�W�DCSCHG �ԛ(��P\g@��PIPL2�S?�i��o�o�o�ZMPC?F_G 1��ii��0'¯S;Ms�S�4�i��p'��g���e2��  ?}�Wν�s������I�~�ꞽ-M���C�=TH�}��)D�C�ҿ��D	I�1��҃ĝ<Ŧ��=�9H�w�������jc���ur��p�pG��t�p��p�x�H�p���}P���Z��~���Ï��y�1���@�G����Y�ڈE�ꄙ�҉�����*�@�N��x��vv�L�R���2���d���x�}�������@=���7�{"�Þ��B��DLW��I�&���B.g��L�?����=k�5�q�? �glp����o�_CYLINuD�� { Х� ,(  *=��N�G�:�w�^����� ��ѯ���7���� <�#�5�r��������� ��޿y�_����8�� ��nπ�㜻ã wQ �5�����S������(�ٻ�X�ז�r�A��SPHE_RE 2���ҿ ��"ϧ������P�c� >�P�̿t���ߪ�� ���'���]�o�L� ��p�W�i���������l���PZZ�F �6