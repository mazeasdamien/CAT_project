��   C��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN��/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER��q�C_GRP6�P L$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� )DEX� �5O n�8BUF�7TDP�HG�_@FO�SxAV��7R?EC_TRQX��MFLG�J5�� � � N IU�
@!(UF*����4OSV3EN_CG"��0_�!�AU�SCH2�SMP]L4PEXE���2�!_�SUR}A�`jAaW�@A@bVNE|Y]QnAVA?�UY�T7D�VWWnAF�[V�A�\�WTO�0oH
e7D�f�3
e�U
e�W QT�P�0IR	 DMM��A@  @ �$la�EREG_�OFS�aME�hA1SS1�A !la�RE-   �# �0�b{F�c{ĥd� M�d�b�c$�STD�hq�gFA � �h!q�g�"�f�"�c�/ la7   �$p`TIN�@��0SUL� �R}_@  $}�@ SW@�rO:}rR%	 dp~t�� �@JU� �s �/ FS4D6
 O� $�0PGF`~QC!$FIL�  �@�E�PmA�s�&�DIG4o@SCA��$�INTT?HRS_BI�AZ��SMAL%�CO�L��qATE_T=I�PROG�4U��s�!CMDAp FSOUTENV6�P $HR�Z_AXl�CU3VR2QLB܊�0���H������PNT_MV_AVR�C�S!pLkp�c$L`���fO�\��ST�:d�F�#STO v��FX�LECTEdDCp�Y{���FY��2t�Z{�ړFZc�!R�e��	�/ G#P��X $��_1IV����$!0�B"0�?0F�CCBwDDN=�CCIc�DUMMY23G ^�DEBU�A\!4PN�"TO�q9RP"�  Q09T6�� �;!��fB'UTTSP� ~@��q֥E40N ڡFS3ՁKQ1�r9T��I�NEW_UQI��VKP?U�p`��CCOORD�8\TCH���01P��mP��7 �l �!�3$�WEIGH���2 Us_�aF��T���WA{Q����NTER�Q��- ޵� �c��r�AS0�$JZA7STA�� �a��P� �,�26�36āW�!Ƨ ��ä"C*��Xw�Yw�Zw�_�CM��?��D��i�RSLy�u���~ɠ�Ǝ��ƚ�	"_Ϡ_�ҡT   �E0c"0VROU�NDCMVPERI}O��$F1PUU37F2D�'TM1� ̯S�_DcGA�MMc1b�TRX��UKt�K�K��C�L�`�&O00ADJ6�GA�UPDC0Rd"���E� QRED����FR_� _@W�۲��u�DL_1R��@�=�M_�5d�0n�#��}�"��}� �k�����������}�VLj�"����@A�7���`��L�P5A8@� 
D�A�����p"��y"��VIBƦ6�OV��DEH�� ���`,����*�� t� RTZ�MN1S�UfMN2YUFR Aq	��ShZA
`-G����OR�P�ҡA1L�ҤCJ��
HL��"�S8B�I$�L .$M�"P30+�Q �)k�}�S"PH�CD�GVz�GVv��GVړJDO°t]��S�$R��E���b�]�A�A�P)�DA��3$#VF�����1LVu��@IL�A���� # �� "�@fR!��$�DC+�����B #ПN�5OBOA@�vYԣW2�G'	�$�ԍ$�!#��E�K�`�+�eC?NPRGOV6��%�'P�t_TW,��"G:�3E�MNV�6�c04WT�cW�TR_L_SKIj�J�q�cN��GW6�
eR^<ENABF�Vq�V!� A$3SB}��xS�� �{P�tyR*�tX�yR QT$���2_Q���?p���ALARM�SER�QETOT~DFRZCHK1����62�9NC�4 N@�5L`N@�:vJ��vE
�22�;2�=NA9E�F'FIX2��BF�䦠�@I�dD���DON��t�95PSFW�0_wDF1"%BF2/_ vJ��|��4|�Pl��33=��5|�kH|�yJP�Z��U�23�;3�=8|�9E�SDIAu �6�RKq�B�VvEfvCM�3GA�@�@�� �R<iV1<d��sP�VQ0�U�Uf�S$��� ���FU�ED�S_HA�U�e�d�4GEF�k@�2�`�; �a��5!%�UzKq�#��X���s����Y��a�_FSI}W� � *�UX�RK��`H7p�_CHCK�!'�INS���w <B
U; �zH�NT���v�y �A`&| ��w�ΰP���8쑎���$����? ���2�=��=� '���SI�Oe�1� � XKC�IRT�U&@0�B�C�,S�V 2n�jp� X  �P������͊@͉	��<����F@ �߀|��B�  =�[�5�a�s����������ŕ=�d=�
ݐh ��������6�X�$� n�W�8�P�b�|���Ւ N�����̯⯨���� *�8�f��n�X����� ҿ����Ŀ���ڿ� �X�jτ�FϘϊ��� ��߲����L�B�p� ߔ�b߸߮�x���6����H��7�I�X��	MC: 56�78  Afs�dt1 78901234q����/  )y� ������.��q�Y�'Q���`� l#�5�B�~P1�+�|�o����� ����������0' 9Rx_�������DMM P����A U�W�(�FXj��POR �2	 [��[��Z1F���B?��S4D7 
!x�	/�'��,/>/��v}?��B�l �e�)***@/�/#!{/��/�C�pONFIoG n���_9�2[�� �$��/ّ��7  �z  D�3025Y��>��P0�e�C  C�3�h1�2DD�/B4�23N �#� 2�,�Ӳ?o��?�:�ד�=���As!�O <O3O��rO]OoO�O�O��O�O�O�O_�� :Z#S8_J_\_n_ �_�_�_�_�_�_�Y_ !ooEo0oioTo�oxo�o�o�I�� 3> [��`h�g A�e�g ��bBk!t�1C�`0�.t��=#�
��N�nk(EuK���QuLE@��eeu=�D��qu��;��=ʁu8I��u��/It$ �$�m5�@rI���uF��3�uBQOGO��x��t��+���E��.���Q���$�{��a�(4$�m��%�7�>�E���B�<~w����8E�=y��;�j��ar���х>��݅��?s ���B�H�g!s >���B A@��?E��qJ��b�@�sF���3Fs�"��E�~�b��vC���C�B��AB������j!AAo!,k!�Bpp#B6q���f!u�@u�@�s @p0@�u�:p7 3�	�	��l�c�u���`�.pݑ Bo C��?���g ݯ��`�?�33���a:�o-�?��a��c� ������������ڿ��?Ls�S�c~�8< ��0����B����� ̻p0%rk�a��8/x���
��<� >�-2��nπ�ߤ϶���e����߾�P��J������� �����V�A����@� ��)qݑ��)r��� �·������	��c�� �oI��+�y����O� a���ڑ��)rk v��l�1��_FCCOORD 32 `!�?����� ��r���
� =�d&�J| ���/��*/� ]//2/�/F/�/j/�/ �/�/�/#?�/�/J?? }?0?R?�?f?�?�?�? �?�?�?CO�?OjO,O �OPOrO�O�O�O�O�O __�Oc__8_�_L_ �_p_�_�_�_o�_�_ >o$oo�o6oXo�olo �o�o�o�o7�o ^D2�Vx�� ���$��W�
�<� ~�d�R�Ïv���ꏬ� �Џ�D��w�*�\� ����r�㟖���
�̟ =���d�&���J�|� ���������د*�� ]��2���F���j��� ޿Ŀ��#�ֿ��J�� }�0�RϤ�f��ϊϼ� ������C����j�,� ��P�r��߆��ߪ��� ����c��8��L� ��p���������� >�$����6�X���l� ��������7�� ^D2�Vx�� ���$�W
< ~dR�v��� /��D//w/*/\/ �/�/r/�/�/�/
? 3��$CC_FSI�W ����>1� K  6M81Y< w?�?�4