��   #��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	  /GR�P: $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2(��� RING��<�$]_d�REL�3� 1  	?���CLo:� � �AX~{  $PS_��TI���TIM�E �J� _C�MD��"FB�V|S �&CL_OV��� FRMZ�$DE�DX�$NA� {%�CURL�W���TCK�5�FMSV}�M_LIF	���;8G:w$�A9_0M:_��=�93x6�W� �"�PCCOYM��FB� M�0��MAL_�EC�I�PL!�"DTYkR_�"�5L#�1'ENDD��o/1 �5M�d �PL� W � � $STAL#TRGQ_M��0KN}FS� �HY�J� |G�I�JI�JI�E#3�AnCuB�A���$��ASS> ����	Q�����@V�ERSI� W  XKQ?IRTUAL_Q�S 1'X W���N �� �_w_�_�_�_�_�_�_ �_.ooRo=jQro`l��O����~����j���%���:�3���[ _o�o[o�l�o�o)&8�kkqrZ������d���<���=L��%�L�3?�M���@�m��� ����ȏڏ����"�04�F�X�� EU��p��{���T  2� �����*�<�N�`�r�����џ���� ү�����,�>�P� b�t���������ο� ���(�:�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z��������<������� � 2�D�V�h�z���������FP��(���� ��,P;M�q ������(��$&4 1b\��O�ڣL���LLay]N9��P�?�M���@�e`C���>B�(�>�A|;� e>��k�A�   �)��	/�� �\n��/l/�/�/��/�/�[}�j�[���/	?z� ��!�/9?�/]?H?�?�?u�%ΐ345?678901�?�4 �-�1���?��O
O@O ROǕ�0rO�O�$ZE�? �O2O�O�O�O_dO5_ G_�O�Oz_h_�_�_�_ �_*_�_N_`_�_�_.o doRo�o�_�_�oo&o �oro(N�ou ��o<����� �j;�����n� ����ȏ�0��T�f� 4���X�F�h���䏵� ǟ�|������B� T���{�Ο��Z�,��� �ү�^�p�A����� t�򯘿����ο$��� �Z���:�(�^�Lς� ��꿻�� Ϛ�l��� $��Hߞϰρ����� ��2��������d�5� G����z�h����� ��*���N�`����.� d�R����������&� ��r�(N��u ���<���� j;���n �����0/T�|2)P(/. �8��$PLCL_GR�P 1��� px5?�  r/�+|?�/x?�/ �/�/�/?�/?I?4? m?X?�?x?�/�?