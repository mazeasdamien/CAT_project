��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1RTU4QQ!Rx1R�� � $TIT91� ��� �Td��T0�ThP�T5�V6��V7�V8�V9�W0 �W�WOQ�U�WgQ�U�WU1�W1�W1�W1�W�2�R  �ASBoN_CF�!@$<!J� ; ;2�1�_CMNT�$�FLAGS]�C�HEK"$�b_O�PTJBL�(CE�LLSETUP o `@HO8@9 PR�1%�c#�aOREPR�hu0D+`�@��b{uHM9 �MN�B;1 UT�OBJ U��0 49DEVIMC�STI/@�� ��@b3�4pB�d�"V�AL�#ISP_UsNI�tp_DOcv<7�yFR_F�@|%�u13��A0s�C_�WA�t,q�zOFFu_T@N�DEL��Lw0dq�1�Vr?1^q�#S?�o`Qb"U�t#*�QTB�����MO� �E' � [M������REV�BI�L���!XI� v�R_  !D�`~��$NOc`�M�|����ɂ/ #ǆ� ԅ��ނ�@}Ded p E �RD_E��h�$�FSSB6�`KBoD_SE�uAG� G�2Q"_��2b�� V!�k5p`(��C�0�0q_ED� � G� t2�$!S�p&-D%$� �#�B9�ʀ_OK1��0] P_C� ʑ0t���U �`LACI�!��a�Y�� �qCOM9M� # $D
� ���@���J_\R BI�GALLOW�� (Ku2-B�@V�AR���!�AB ]`BqL�@� � ,Kțq���`S�p�@M_�O]˥��CC�FS_UT��0 @"�A�Cp'��+pXG�܂b�0 4� IMCM ��#S�p�9�H��i �_�"t� t��M�1 h$�IMPEE_F� s��s��� t�����D_�����D��F��L�_����0� T@L��L�D�I�s@G�� u�P�$Iȼ'����CFed X@GRU@��=Mb�NFLI�\��@UIRE�i42�� SWITn$`0_�N�`S 2CF�0M�� �#u�D���!��v`����`J�tV��[ E��.p��`�ʗELBOF � �շ�p`0���3����� F�2T��0A`�rq1J1��z _To!��p��gt���G� �r0WARNM�p#tC��v`�ç` � CORz-UrFLTR��/TRAT9 T%p� $ACCVq��� |��r$ORI�,_&�RT��S<����HG�0I���T�W��A�I'�T�rM�K�� �20p2�a1��HDR�2
��2�2J; S���U3��4��5��6��7��8��9KD׀
 ��2 @� TR�Q�$vf��'�1��<�_U<�G�_:�{COec  <� �P�b�t�53>B_�LL�EC��!~�MULTI�4�"u�Q;2�CHILD��;1���@T� "'�S�TY92	r��=��)�2�������ec# |r056$J ђ�a�`���uTO��:�E^	EXTt��p��2��22"�0����$`@D	�`&̒�p������ %�"��`%�ak�����s�`���&'�E�A�u��Mw�9 �% ���TR�� ' L@U#9 ���=At�$JOB�����P]`|IG��( dp������^'#`j�~ǝ�pOR�o) t$�FL��
RNG%Q@�TBA ΰ �v&r�*`1t(� �0 �x!�0�+P�p�%,/��*��͐U�Гq�!�;2J�_R��>�C<J�8&<J D`5CF9���0x"�@J��P_p�n7p+ \@RO"p�F�0��IT�s�0NOM��>Ҹ4s�2��J @U<PPgў�P8E,|Pn��0�P�9�͗ RA���l�?C��� �
$TͰtMKD3�0T��pU�`��΀+AHlr>�T1�JE�1\�J���PQ���\Q��hQCYNT|�P��PDBGD̰2�0-���PU6$$P0o�|�u�AX�����TAI�sBUFp,����A�1. ���l�F�`PI|�-@PvWMuXM�Y�@�V�FvWSIMQST}O�q$KEE�SPA��  ?B�B>C�B��A��/�`��MA�RG�u2�FAC<q�>�SLEW*1!@0����
۾ s�CW$c0'���pJB����qDECj�exk�eaV%1 Ħ��CHNR�MPs�#$G_@�gD�_�@s���1_FP�5�@TC�fFӓC�Й���qC���+�VK�*��"*�J�Rx���SEGFRf$`IOh!�0STN�gLIN>�csPVZ�z�Ц@�D2����r� 2��hr�r�2��3` +^?���եq �`��q|`�����t��|aSIZ#�!�� �T�_@%�I��qRS�*s��2y{�Ip{�pTpLF�@�`��gCRC����CCTр��Ipڈ�a���b��MIN��a1순���D<iC �C/���!u`c�OP4�n j�EVj����F��_!uF��N@����|a��=h?KNL�A�C2�AVSCA�@A��1�a��4�  cSF��$�;�Ir ��Q�&��05��	D -Oo%g��,,m�����ޟ��RC�6� n���sυ�Uz��R�0HANC���$LG��ɑDQ$ft�NDɖ��AR۰�N��aqg��ѫ�X�M�E��^�Y�[PS�RAg�X�AZ�П���rEOB�FCT��A��`��2t!Sh`0ADI��O��y�s"y�n!�� �����~#C�G3t!N��BMPmt@�Y�3�afAES$������W_;�BAS#X�YZWPR��*��m!��	M�U�87  ƀI@d���8\�p_C:T���#�- ��_L
 � 9 %���C�/�(zJ�KLB�$�3�D�<�5�FORC�b�w_AV;�MOM*�q�SaԫBP`Ր�yӐHBP�ɀE�F����A�YLOAD&$EAR�t&3�2�Xrpx�!!�� R_FD��_ : T`I�$Y3��E�&��Ct��[MS�PU
$(�kpD��9 �b�;��B�	EVId�
��!_IDX   $���B@X��X<&�SY5� �zR_HOPe�<>��ALARM��2W̭s�qR_�0= !hb Pnq�`M\qJ@O$PL`A&�M#�$�`��� 8�	��ҨV�]�0�$�U�PM�{�U��>�TITu�
%�![q�BsZ_;���? �B� pQk��6NO_HEADE^az��}ѯ ��`􂳃���dF�ق�t����@�@��>uCIRTR�`���ڈL��D�CB@4�R�J����[Q���1A�2>���OR�r���O����T`UN_OO�Ҁ$����T�����I�VaCnpO ?DBPXWOY���=B�$SKADR��DBT�TRL
��C��րfpbDs�L�~�DJj4 _�bDQ}��PL�q�wbWA���WcD��A��A=�2�U�MMY9��10L��0DB����D;v[QPR�� 
M8�Z���E O�Y1�$�a$8��L)F!/_c���0yGG/��9�PC�1�Hf/�2�PENE
A@Tf�I�/��,$��COR`"JH y@ �E$L�#F$#PR���+jp���nq�_D$�qPROSS]�
���R�r�` >u�$TRIG96�PAUS73ltETgURN72�MR:�eU 0Ł0EW$�~�`SIGNALA��QR$LA�З5�1�G$PD�H$PDİ�AI�0�A�C�4�C��DO�D�2�!��6GO_AWAY2MOZq�Z�W �DCS��CSCB�g�K Իa#���E+RI�0Nn�T�`$�����FCBPL�@QBGAGE���P��ED`|BD�wA[CD�OF�q�[F0�FoC��MPM�AB0XoC�$FRCIN��2Dk��@��O$NE�@�FD�L8�� L� �����=��Rw�_��P>� OVR10����lҠ�$ESC_|�`uDSBIO��p��pTe�E�VIB�� `s��Z��V��p�SSW��$�VL��:�Lk��X���ѣ�0bQ����USC�P��qA=�	Q��MP1%e@&S*`�(bt`'c5۳ESUd��-cWg&S Wg?cWd����Wd��Wd<.���AUTO$�Ya҃�ac�SB����-d���&SwB[��GB�f_$VOLT�g ���  �GAOD!��q���@:�ORQ�ҀKra�$DH_THE&0�Rgp� <qtnwALPHnt��o��w0 Vp]�$�.�Ra�[��s�5�`r�CQ�#BUD�S� F1M���sV
��;��L�b�tk���BRTHR��L��T`�Z���Vɖ��D)E  �1��2�⋅ ��������kѯ�a� �Tt0V�ꆸ������@̈Я�-�"�N~���sS2����INHB��ILTG0ɡ�T?� �3$�w��E��PqQxQ��TqPe��0Y�AF}�O�ນ��ڗ ��qPڳē����bPܙ���PL?���3���TMOU��ēS��� � ��s�/�S18���O��Aܙ��I����CDqIƑ˩o�STI��գ�O:ҋ�,0���AN��Qg�S��+r�#x$�����w�1_����PRA�P`�vC����MCN�eQe�����VER�S��r�oPIw�F�PåǲШ۷G.�DEN��G>�����F�2H�Ƿ�M�7�F��_�MN�D̠,���@�d�{ƭa����OB����U˱z���DI ���#���3�����A��w�Fx���3�O�N�5��Q��VAL��CR[�_SIZp��b�;Qn�REQ�R�b��]2b���CH q�΂�ڃ�Ռ�����:�n�S_U��X��wW�FLG���wU$CV�iMGP�QδFLXP�923R�u�L��EAL�P-�C	�F+rT��W��� �R��c���NDMS�7� ��K>S�P_M'0h�STWv������AL�P���Q����U���U�IAG@,�o��d�U�-�T"	A-`� ���A��� ��H`��Q`��6��Pq_D&��1s��.�P��F�>2�T�� ?7 1A>���#�#L��?`_=i @@>LD�pc�F�0�FRI�0 `Ѐ��1}Ѳ�IV\1�*�^1�U�P`��a��C�L!W��
`L=S&-c&&S�C.w��  L���!����d�Q$w!�҇��$w��p��
�P�5RSM��P���V0h � r�l�d^2AW�a_TRp�}�8@NS_PE�A����< ��$�SAVG�8�6G]%���CAR �`�!�$���"CRa���$ d�#qE�@��"STD���!Fpo��'QOF0��%��"RC���&RC۠�(F�2A�R#7����%, gMA�Q_�a��
QQ��al2��%u4Ib�r7I�R�9�wQ�7�8M/��!C:pR�  �p�2F<�SDN�a  � W2QM P $Mi��s$cA �$C�cm�9���4���AT�0CY_ �N LS!IG1@x'yB��y@@H2Y��NO����SDE�VI�@ O@�$�RBT:VSP0�3�CuT�DBY|�A�	W`3CHNDGD�AP H@GRP�HE iXL�U��VSЌFx2� DL1p aQ6ROp��FB�\]�FEN�@��S���ChAR d�@DyOd�PMCSb���P薇P�R��HOT�SWz42�DMpELE�1/e��C8`�RS T�@���r� hfl��`OL�GHA�F8k�Fs�� 
�D�A�@T � $M{DLUb 2S@�E���q�6�q	0�i�c�e�cJ��	uݢ�#�~5t+w�PTO���� �b���CSL�AVS� U  ��INP �	V�Њy�A_;�ENUAV; $R�PC_�q�2� 1bL�w�0 �tS{HO+� W ���A�a�q�2�r�v�u��v�sCF� X` ,f��r�OG gE��%D�h�lp�C�Iߣi�MAX��D�x AY?�W� �p�NTV	�D�VE\�0@�SKI��T�`Hg?Ň2�� JZs��! Cꆻ��f�_�SV/ �`XCLUt��H���ONL���'�Y�T��OT:eH�I_V,11 APPLY��HI4`;�U��_ML�� $�VRFY8�	�U�M{IOC_I���J �1/��߃O�@X�L�Sw"`@$DUM�MY4���ڑ�Cd L_TP���kC��^1CNFf���E ��@T�y� D_#UQa_��ݥ�YPCP��@=�� �����|��$����� Y �+�
0RT_;P��uNOCCb Z�r�TE���=�פr�DG�@[ D��P_BAe`Lkc�!��_���H�~T��E �\�pAb=cAR�GI�!$���`[SGNA] �8�`U��IGN�Տ�,�� ��V����>��ANNUN��&��˳�EU�J'�ATCH��J��Md�rA^ <@g�����&:c$Va����X�ᑴaEF] I��_ _ @@FͲ�ITb�	$TOT�i �C�O�c�rpEmM�@NI�a`tB���c���A>���D{AY@CLOAD�D�\�n���� �[EF7�XI�Ra���K���O%��a ��ADJ_R�!@b"��>�H2�"[�
 Hc�%��`a͠MPI��J��DHЏ�?�Ac �0��х�� ��Z��ϡ�Ui ��CTsRL� Yp d���TRA8 ?3IDLE_PW  �Ѡ��Q��V�GV_���`c� �o�;Q@e�� 1$��6`<cTAC-3��P�LQ�Z�Rz\ A-u:ɰSW;�A\����/J��`b�K�OH��(OPP; �#IR9O� �"BRK��#AB �O������@� _ ���F���`d͠x, j@S�RQDW��MS�P6X�'z��?IFECAL�� 10^tN��V���`��V�(0��CP
���N� Yb�0FL�A_#�OVL ��H�E���"SUPPO��ޑ\�L�p��R&2X�$Y-
Z-
W-
��/��0GR��XZ�q�$Y2�C	O�PJ�SA�X2R���*r�!��:��"trex0��0)�f `�@/CACHE��c؛�0�s0LAZ SU7FFI, C��lq\���6�~RM�SW�g 8�K�EYIMAG#TM�@S��n
2j�r|���ROCVIE���~�h �aBGLx����`�?� 	NaԚ��i��!`STπ!������������EMAI��`N��`A�@Z�FA�U� �j�"lq�a��U�4�u E�}�k< $dI#�US�� �IT'��BUF`��DN�B���SUBu$�DC�_���J"��"SAV �%�"k������';�r�P�$�UORD���UP_u �%��8OT�T��_B`��8@LM0l�F4��C7AX@Cv�b��Xu 	��#_G��
rpYN_���lT6���D�E��M��U��T��F��cavC�DI`BEDT)@IC��~�m�rI�G�!"c�&��l`��!��P���FZP n (�pSV� )d\�ρ����QA��o� �����>"$3C_R�IK��kB��hD{p�RfgE.(ADSPd~KBP�`�IIM�# �C�Aa�A��U�G��4�iCM! IP��KC��� �DTH� �S�B2*�T��CHS�3�CGBSC��� ��V�d�YVSP�#[T_DrcCONV�Grc[T� $�Fu F�ቐd�C�0�j1��SC5�e]CM�ER;dAFBCM�P;c@ETBc mp\FU DUi b��+�~�CD�I�%P702#@O���qWӏ�SQ��QǀSU���MSS�1ju�4`�T葡Aa��A�1r�� "�Й��4$Z!O@s���l�U6�&�2�eP���eCNc�l�x�l�l�iGROU�Wd)��S c�MN�k Nu�eNu�eNpR|b|�i��cH�pi��z
 �0CYC���s�w�c�6�zDEL�_D��RO�a���qVf���v{�O�2���1��t���:R�ua�.#� ��A	L� �1sˢI1¡��J0�PB��D  ERr^�T�Gbt ,!@���5��aGI1LcR1gs 
F ԠNO���1u���������P����Cڠ	�������1��J0�0vH *	�LU�1#J�Q� �V
�[�7Az���z�쑀z���z��z�Fz�7
w�8w�9w���y���U1��1��1��1��U1Ě1њ1ޚ1뚥2��2����2��2���2��2Ě2њ2�ޚ2�3��3��3T����3��3��3ĚU3њ3ޚ3�4��&�bXTF��1w6�.(��0�f�0�U�0ŷ�e���FDR5�xTU VE��?1���,SR��RE�F����OVM~C)�A2�T7ROV2�DT� R�MXa�IN2���Q�N2�INDp�r�
���0�0�0Gu1��[�G`��{�D_�[�RIVx�P�b�GEAR~AKIOr�K"N�0��y�p�5`@�a�Z_MCM� ������UR�Ryǀ��!?g ��p?n�.��?n�ER�vѐ=a�!�P��zI:�PXqB�RI0%�`�#�ETUP2_ 3{ ���#TDPR�%TBp������I ��wBAC�2| T��"�4)�:%	`^B��]p�IFI��� 1Mc���.�PT��!�FLUI�} 1� ��K UR�c!����B�1SPx E�EM�P�p�2$��S^��?x��Jق0
3V�RT���0x$SH�O��Lq�6 ASS�cP=1��PӴBG_ ��������FORC3"f�d[~)"FUY�1�2�\�2�1�h� p�� |��NAV�a)�������S!"�c?$VISI��#�SCM4SE����:0jE�V�O��$��X�M���$��I���@�FMR2>��� �5` �r�@�� �2�PI�9 F�"�_���?LIMIT_1�d�C_LM������D�GCLF����DY&�LD����5����$�ĸ�M�Fc�D!u	? T�FS0Ed�� P��QC�0�$EX_QhQ1Pi0�P�aQ3�5�s�GoQ��� ���6�RSW�%ON�PXÏEBUG��'�GiRBp�@U�SBK)q�O1L� ��P�OY 
)��P��M���OXta`SM��E��"�a���`_E � �0�� �T�ERMZ%�c%��O�RI�1_ �c'�KSMepO��_ �c&h�`�`�(��)UP>� �� -��F�b���q#� ���yG�*� ELTO��p�0�PFIrc�1Y���P�$�$�$UFR�$��1L0Le� OTY7�PT4q��k3NST�pPA�T�q4PTHJ��a`EG`*C�p1ART� !5� y2$2�REL�:)ASHF�TR1�1�8_��R(�Pc�& � $�'@��� ��s�1 @I��0�U�R G�PA�YLO�@�qDYN_k���.b�1|��'PERV��RA��H�� g7�p�2�J�E-�J��RC���ASYM�FLTR�1WJ*7����E�ӱ1�I��aUT�pbA�5�F��5P�PlC�Q1FOR�pM�I!����W��/&�0F0�c�9H��Ed� �m2N�,��5`OC1!?�$OP����c������bRE��PR.3�1a�F��3e��R�5e�X�1(�e$PWR��_����@R_�S�4��et$3�UD��$�R72 ����$H'�!^�`ADDR�fHL!�G�2�a�a�aT��R���U�� H��SSC����e-��e���eƪ�SEE��HS{CD��� $����P_�_ B!rP􍀌�� �HTT�P_��HU�� (��OBJ��b(��$�fLEx3Tt��� � ���ะ_��T?#�rS�P��z�sKRN�LgHIT܇ 5��P���P�r������PL��PSS<�ҴJ�QUERY_FL�A 1�qB_WEBwSOC���HW��1U���`6PIN'CPU���Oh��q�����d���d���� ��IHMI_ED^� T �RH�;?$��FAV� d�~ŁR�IOLN
◓ 8��R�@�$SLiR$INoPUT_($
`���P�� ـS�LA� �����5�1��C��B��I�O6pF_AS7��$L%�}w%�A��\b.1�����T@HYķ����E�h�wUOP4� `y� ґ�f�¤�������`PCC
`����#��>mQIP_ME��7� Xy�IP�`�U�_NET�9����Rĳs�)��DSaP(�Op=��BG`�p����A��� lp�:CTAjB�pAF T�I�-U��Y ޥ�0PmSݦBUY IDI��rF ��P�� ��� �y0�,�����Ҥ�NQ�Y R���IRCA�i� ך ěy0�CY�`EA�����񘼀�CC����R�0�A�7Q�DAY_���NTVA����$��5 ����SCAd@��CL���� ������8�Y��2e�o�N_��PCP�q��ⱶ�� ,�N����
�xr���x:p�N� 2�����(ᵁ����xr۠�LABy1��Y ��U�NIR��Ë ITqY듭��e��s��#�5���R_U{RL���$AL0 �EN��ҭ� ;�T��T_U��ABKsY_z��2DISԐ��AR�Jg�����P�$���E��g�R���З A�/���J����FLs��7 Ȁ|���
�UJR� ���F{0G��E7��J7 O^ R$J8I�7�H�R�d�7��E�8{��H�APHIQ�S��DeJ7J8�B��L_KE*� � �K��LM�[� � <X�X�Rl�u���WATCH_VA��o@D�tvOFIELc��cy.L��4� � o1Vx@���-�CT[�9�m��_C�LGH���� $��LG_SIZ�t�z�2y�,p�y�FD��Ix��� +!��w�\ ����v��S ���2��p��������\ ���A�0_gCAM]3NzU
RFQ�\vv�d(u�"B��2�p����I��+ �\ ���v�RS���0 } �ZIPDUƣ�p�LN=��ސ �p�z6���f�>sDr�PLMCDAUi�EAFp���TuGqH�R��|�BOO�a?�� C��I��IT+���`��RE���SCR� �s���DI��SF0�`RGIO"$D�����TH("�t|�S�s{�W$�|�X��JGM^'MgNCH;�|�FN��ba&K�'uЅ)UF�(�1@�(FWD�(HL.�)STP�*V�(%�X�(��(RS9HIP�+��C[T�# R��&p:'^9U=q�$9'�H%�C𜓚"Gw)�0PO �7�*��#W}$���)�EX��TUI�%I ���Ï���rCO#C�� *�$S��	�)��B@�NOFAcNA|��Q
�AI|�8�t:��EDCS��c��C�c�BO�HO�GSȅ��B�HS�H(IGN�����!O���D�DEV<7LL�����-��Ц(�;�T�$��2�p�����*�#A���(�`뀸{�Y��POS1�U2��U3�Qˑ�2�@�Ш# ��{�PtD�� ��&q)��0�d��V+STӐR�YU�B@~ ` �$E.fC.k�p<p=fPf5�Sh��Щ LRТ�  ��x�c�p��<�Fp�dxY�@!�_ ������Kq&���c�{MC7� ����CLDPӐ��TR�QLI#ѽ�ytFAL��,r�5s8�D�5wS�LD5ut5uO�RG��91HrCRESERV���t���t��c�� �� 	u95t5u��PITp��	xq�t�vRCLMC�������qF�M��k�������$DEBUGMAS��ް��?%U8$T@��Ee�g���pFRQՔ�� � j�HRS�_RU7��a��A<��k5FREQ� ��$/@x�OVER���n��V#�P�!EFI �%�a��g�8ǒ���t� \R�ԁ�d�$U�P��?��p�PS�P��	�߃C��͢a��U�\�l�?(P�/PMwISC� d@��QRQ��	��TB�  � Ȗ0A՘A�X����ؗ�EXC�ESj�A4<���M���\��������c�_:��SC�P '� H��̔_��Ƙ�ǰ]����MK�HԳK�J� m�B_^K�FLIC�dB��QUIREG3MO���O˫3�<�L�`MGմ �`��T�t���Y�MNDU��]��>��k�G�D|f��INAUT����RSM>�a��@N��r]3-��a5�PS�TL\�� 4X�L�OC�VRI%��UEXɶANGuBu��q�ODA����������MFO�����Y�b@�e4�2k�S�UP�eQ�FX��I�GG� � � �p�c���cQ6�dD� %�b|�!`��!`��|�0�3w�ZWa�TI��p�;� M��[�� tV��MD��I�)��@���HݰM��GDIA�����W,!P�wQ�1�D�)��qO���]�� 0�CU��VP��pu���O!_V��ѻ �`��S�X�5����B��P��0N���P���KES2���-$B8� ����ND2�����2_TX�dXTcRA�C?�/��M�|q�`�Pv��XҰ��Pt SBq`�USWCS��T��	����PULS��A�NS�ޔ��R��JOI�N��H��~`j�=���b��b�����P=�`�$��b$���TA��@��S���S�HS�E��SCF�aPJ��R��{PLQ� ��LO��н.���^� ��8��������0�RR2���� 1��eA�q Kd$��Iΐ+�G�A�2+/� ΍PRIN�<$R SW0"�a/�wABC�D_J%�¡���_J3�
��1SPܠeЛ�P���3��р`��B�J/���r�qO8QyIF��CSKP"z�{�{�J���Q�L2LBҰ_A1Z�r�~ELQ��OCMPೕ�T����RT�����1�+���P1��>@�Z�SMG0��=�;JG�`SCL�͵OSPH_�@��%�VЛ� RTER0`  �< A_�@G1�"�A�@c��\$D�I�
"23UDgF  ǀ~ LW�(7VELqIN�b)@� _BL�@u��$G �q�$�'�'�%`<�� �ECHZR/�TSAY_`� ���E}`B<����5�B���1:}`_�� �)5D2d%�A4I��N9t&R�DH�A���ÀP�$V `�#>A$���Ͳ�$Q�R}ӆ��H �$BELvᵆ<!_ACCE�!c��7</��0IRC_] ���pNTT��S$PS�rL� d�/E s��F{�@F
��9�gGCgG36B���_��Q�2�@�A���1_MGăDD�A]"ͲFW�`���3�EC�2��HDE�KPPAByN>G��SPEE�B �Q%_pB�QY�Y��1>1$USE_��,`]Pk�CTReTYP��0�q P�YN��A e�V)хQM����ķ��@O� YA�TINCo�ڱ�B�DՒ�WG֑ENC����u�.Ax�2Ӕ+@INPOQ�aI6Be��$NT�#>�%NT23_�"�2�IcLO� �2_`��I �_�if� _�k�? �`� ej�C400fMOS�I�A���ОA䃔�P?ERCH  �c��B" �g��c��lb=������oUu@�@	A6B(uLeT	~�1epT�ljgv�fTRK@%�AY��"sY��q6B��u�s۰�]��RU�McOMq�ՒY�MP�^��C�s�CJR���DUF �BS_BC?KLSH_C6B)� ���f���St�H��RR�|�QDCLALM-dp���pm0��CHK|���GLRTY����d��Y��)Üd_UM]�ԉC��A!��=PLMT� _L �0��9��E�.�  ��#E)�#H� =��Q�3po�xPC�axHpW�頿EׅCMCE�\�@�GCN_,ND�LΖ�SF�1�iVoR���g<!��6B���CATގSH)�,�D fY��f��7A���f܀PAބ�R_P݅�s_ �v���s,����JG�T]����Y�����TORQU`aP��c�yPOU��0�b��P%�_W�u�t���1D��3C��3C�I*K�IY�I�3F�6������@VC�00RQ�t��1���@ӿ��ȳJRK�����Up�DB M��UpMC� DL�1BrGRV�J�Cĭ3Cĳ3$�H_p��"�j@q�COS~��~�LN���µ�� �0�����u����̓�b�Z���f$�MY���؊���>�THE{T0reNK23�3�hҧ3��CBm�CB�3C! AS� ��u�0�ѭ3��m�SB�3��Nx�GTS$=QC������������$DU��Kw�B�%(�
�%Qq_��sq��x�{�K���b(��\�A�`Չ��p�{�{�LP!H~�g�Aeg�Sµ�� ������g������֊��V��V��0��V���V��V��V��V*	�V�V%�H��������G�����H��H���H	�H�H%�OJ��O��OV	��O��UO��O��O��O	�O�O�Fg���	������SPBAL�ANCE_-�LmE��H_`�SP!1��A��A��PFULCElTl��.:{1��UTO_�����T1T2��22N���29`�!�qnPL�=B�3�qTXpOv |
A4�INSEG�2��aREV��`aD3IF�uS91�8't"1�6`OB.!t�M���w2�9`��,�LC�HWARRCBAB�� ��#�`-ФQ 5
�X�qPR��&��2�� 
�""��1e7ROB͠CR6B5���  �C�1_���T � x $WEIGH�PFrp$��?3àI�Q�g`IFYQ�@LAGĒRq�S�R �RBI�Lx5OD�p�`V2S�T�0V2P!t�W0P�01�&1/0�30
�Px�2�QA  2řd^[6DEBUg3L_@z�2�MMY9&E� Nz�Drp$D�_A�a$�0��O� �  �DO_:@A.1� <B0�6��m�Q�B�2�0N�-cdH_p`�P �2O��� �� %"��T`"a��T/!�4�)@TICKh3| TE11@%�C ��@N͠�XC͠R?��Q�"�E��"�E8@PROMP��SE~� $I�R��Q��R;pZRMCAI)��Q�R4U_r0C2S; �q�PR8�7COD�3FU�Pd6ID_[�vU R!�G_SUFFu� �l3�Q;Q�BD�O�G �E�0�FGR r3�"�T�C�T�"�U�"��Uׁ�T8D�0�B0Hnb _FI�19*c7ORD�1 50�2�36V�+b�Q1@$�ZDT}U���1;E��4 *:!L_N�AmA�@�b�EDEF_I�h�b�F�d�E�2��F�4�F�c�E�e�FISP��PAKp�Ds�C�d��44בi��2�D�"�It�3D�O|#OBLOCKEz���S�O�O�Gq�R�PUM�U�b�T�c�T�e�T !r�R�s�U�c�T�d�R �6�q�S� ���U�b��U�c�S�Z��X�@P@` t�@qe�)@W�xt���ss0�TE��<D�( l1LOOMB_��ɇ0V2wVIS;�ITYV2�A��O�3A_FR1I��a SIq�BQR�@��@�3�3
V2W��W�4����9_e��QEAS^3�R@ϡ��_�[p:R�4��5�6_3ORMU�LA_Iz���T�HR^2H�Gtg��30f��<8�5COEFF_O�A	 ��A���GR�^3Sg0BC�AnO/C$��]3a�_:�1GRP� ?� � $�p�YBX�@TM~w���u��B�s��bCER, T�ttsd�0�  �L�L�TSpS~�_SV Nt�ߐ���0�����0� ��SETUsMEA*P�P���W0�1+b/0� � h��  @ڐo� l�o�cqz��b�@cqq`tP�G��R�� Q\p*q[p��>�c �NPREC>at��5@MSK_$|��� PB11_USER�e"�{ ���VEL���{ 0��$Ō!I]`��MT�ACFG��� � �@@ O�"NO�RE-0l@o�V�SIb.1�d��6�"UXK��fP!��DE�� �$KEY_�3>�$JOG�� SV������!��}��SW�"�a\aS�ՐT�|�GI���| ^�� 4 h��'d2�!XYZc���3z� �_ERR#�C� 8Ԡ�AfPV��d��1����$BU�F��X��_M_�M�OR|�� HB0CUd�lA�!��GQ\aB�<,"!a$� ��9�a����_�?��G~�� � $cSIՐ���VO��<T� OBJE_���ADJU)B��EL�AY���%�DR�O�U.`=ղВQ0b=��T���0���;BDIR���; I�"�0DYNW�#���T���"R���@�0�"��OPWORK����,%@SYSBUy�SOP��ޑ�U�; P�pN�<��PA�t�>�"��OP�PUd!0�`!�Ľl�IMAGw��B0y�2IM�Õ�I�Ne�d��RGOVCRD��-��o�Pq����0��J�Os���"L�pBa���o�PMC�_Ee`���1Ny M� A�21�2�S�L_��� � $OVSL�ǫ�?qD�`��2�" -�_�� k�P��k�Pu���2�C� �`�Ź�^��_ZER�D��$G�� :82=���� @*����%Oh`RI��� 
 JP8+T�=!/��L��ح�T� �0A�TUS��TRC_T���sB��}f�s�9s�1Re`��� !DFAm����L���"`��0a� ޱ��XEw {�����C0�vUP��+p	qPX�P�j�43 ���PG\���$SUBe�%�qe9JMPWAIT ,z}%LO��F�A�RCVFBQ�@x"�!qR�� �x"ACC� �R&�B�'IGNR�_PL9DBTB2�0Pqy!BWbP�$2w�Uy@�%IGT�P=I��TNLN�&2�R��rL�NP��P�EED \HADCOW�06�w��E[pq4jO!�`SPDV!� LbAz�`�07�3UNIr��02"!R��LYZ`� �o��PH_PK���e�RETRI�E9{�q����0'PFI"�� �G`�0D� 2�g�DBG�LV�#LOGSIYZ��EqKT�!U��2VDD�#$0_T�G��MՐCݱ��|@eMR�vC}�3�CHECK�0��H�PO�V!�2k�I��LE(!���PArpT�2K�W���@P2V!� h $ARIBiR� c��a/�O�P8�ӐATT��2�IF|@z�Aq�4S�3UX���T�PsLI2V!� $g����ITCHx"[�W� �AS9�wSL�LBV!�� �$BA�DYs��BCAM!���Y9�P#J5��Q��R6�V�Q_KNOW�Cb���U��AD�XV��0D��+iPAYLOAt��Ic_��Rg�Rg�ZOcL�q��PLC{L_�� !7���b�QB��d���fF��iC֠�js��d�IB�hRؠ�g�ҢdB��2��J��q_J�a#���AND��Ĳ.t��b�a�q�PL0AL_ �P�0�Ш�QրC��DNcEά��J3CpWv� =TPPDCK����|��P�_ALPHgs��sBE��gy|��K�1�� � ����HoD_1Oj2ydDP�AR�*��x;�&���TIA4U�u5U�6��MOM��@a���n���{�Y�B� �ADa���n���{�PUB��R��҅n�҅�{��2�Wp��W � � PMsbT�� �2xQ���� e$PI��81�@�TgJ��niJ�IV�Id�Ir��[��3!��>!��r�Ӫ�U3HIG�SU3�%�4 얎4�%� ���"�����!
��!�%SAMP ���^��_��%�P4s ю���[ 	� ��3 ���0���&���@����^��Sp��H&0	�IN�SpB�����뤕"��6��6�V�GAMM�SyI�� #ETْ��;�D�tA�;
$ZpIBR!62]IT�$HIِ_��H����˶E��ظAҾ���LWͽ�
���@7���rЖ,0�qC�%�CHK��" �~I_A�����Rr �Rqܥ�Ǚ��ԥ��ɾWs �$�x �1���I7RC�H_DA� RN{��#�LE��ǒ!�,��x���90MSWsFL�$�SCR((G100��R@��3]B ��ç��a����َ0���PI3A9�MET�HO����%��AX�H�XX0԰62ESRI��^�3��R�0$u	��pF{�_���I?ⲣ1�L�L�_�a�OOP����wᜲ���APP:���F����@{���أRT�V�OBp�0T����;��� 1�I��� ���r���RA�@MG�A1B&�SV-��;P�CURg�;��GRO[0S_SaA�Q��Y�#NO�pC!"�tY��Zo lox�������!b����&�DO�1A���A�� ��Х��A���A"�WXS�c sTM)��� � ��YL(H�qܧ��SrZ� ]B�o��0��ĵq�_�C1��M_W����g���c�M@� �`Vq�$pԐx1o�3"�PMJ�,��C �'A� 9�!Wi:�$�LWQ|ai �tg�tg�tg{t� ��N`���S��SpX�0O�sRqZ��P� �*�� ���M�� ������������X���X ��@�qPL�q_~R� |�q#(Y����& n��&{�Y�Z��'�&t���Q���4�#0��qP�}`�$PQ�PMO�N_QUc� �{ 8�@QCOU��n%PQTH��HO�n^0HYS:PES�RF^0UEI0O��@O|T�  �0PGõz�RUN_TO�q:�0ْ.�� PE`�5C��A<�IND}E�ROGRA�nP� 2g�NE_NO�4�5IT��0�0�INFO�1� ІQ�:A�ȇOI�B� (��SLE�QݖFAѕF@�6eOySy�T� 4�@�ENAB��0PT�ION.S%0ERV�E���G��� zCGC]F�A� @R0J$�Rq�2���R�H�O�G "�EDITN�1� �v�K�jޓʱE�NU0W�*XAUTu�-UCO�PY�ِN\����M�ѱNXP\[q�PRU�T9� _RN�@OUC�$G�2�T�p��$$CL`?0[��&���a�a� �P�S�@�X��PXK�QIGRTU��_�PA� _WRK 2 e��@ 0 � �5�QMoYh\Jo|m |l	�`�m�oa�`��o�o�f�e�l}�aI�[ct'`BS�*� �1�Y� <7����� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P��b�t���������srC�C��LMT?0����s  dѴIN�ڿ�дPRE_EXE��)�Ƅ0jP���za'`DV��S��@e)�%s�elect_macro����kϤ�qt�IOCNVVB�� 5��P��USňw����0V 14kP $$p��a�|�`?���߰>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ ���$�ѰLARMRE?COV ^������LMDG ��Ь�LM_�IF ��d�  YST-04�0 Operat�ion mode AUTO S��ed P) )�t.(L:6)�� ����)�;�M�_�q�~�, 
 ����#�>TELEO�P ǘLINE Y6ǑقPA��DǙ�JOINT 10�0 %�����$8���@�$�@���ATAǒ0ǐ3���������  clear䀪���ί���NGTOL  >@� 	 A\����ѰPPINFO7 �� f�L�p^�p����  �� ����k���ۿſ��� ��5��Y�C�iϏ�%���ٯ��������� �'�9�K�]�o߁ߓ����PPLICAT�ION ?t���|��Handling�Toolǖ 
�V9.40P/1}7\�
883ǀ�����F0�	�54�9��������7D�F5�О�ǓNon}e��FRA��� ؒ��,�_A�CTIVE1�  ��� �  ��ڀM�OD��������CHGAPONL��� �OUPLE�D 1	��� �>�B�T�f���CUR�EQ 1
��  UTp�p�p�	�� ������l��������������i3l�;p���^�H��A�t
HTTHKY�FXv |��*<N `������� �//&/8/J/\/�/ �/�/�/�/�/�/�/�/ ?"?4?F?X?�?|?�? �?�?�?�?�?�?OO 0OBOTO�OxO�O�O�O �O�O�O�O__,_>_ P_�_t_�_�_�_�_�_ �_�_oo(o:oLo�o po�o�o�o�o�o�o�o  $6H�l~ ��������  �2�D���h�z����� ��ԏ���
��.� @���d�v���������Ƃ�TO�����DO?_CLEAN���E�NM  �� p�������ɯۯ�v�DSPDRYRLL���HI��o�@�� G�Y�k�}�������ſ�׿����ϻ�MA�X��,�����=�X�,���9����PLU�GG,�-�9���PRUC��Bm�q�6��(ϗ�O����SEGF�K���� �m� �G�Y�k�}ߏ�����LAP$�7ޡ���� ��+�=�O�a�s������ �TOTA�L_ƈ� �USENU$�1� �������RGDISPM+MC�d�C�O��@@�1�O"�D���-�_STRIN�G 1��
��M��S��
~��_ITEM1��  n���������  $6HZl~ ��������I/O SI�GNAL��T�ryout Mo{de��InpN�Simulate�d��Out`�OVERR!� �= 100��I?n cyclT���Prog Ab�orj��JSt�atus��	Heartbeat���MH Faul<��Aler�! /!/3/E/W/i/{/�/�/�/ (���(� ���/??&?8?J?\? n?�?�?�?�?�?�?�?��?O"O4OFO�/WORИ�~A�/XO�O�O �O�O�O __$_6_H_ Z_l_~_�_�_�_�_�_�_�^PO���"` �KoEoWoio{o�o�o �o�o�o�o�o/�ASew��bDEV%n�p9o��� �#�5�G�Y�k�}��� ����ŏ׏�����|1�C�PALT�- j��OD�������ȟڟ ����"�4�F�X�j��|�������į֯X�GRIB�������6� H�Z�l�~�������ƿ ؿ���� �2�D�V�h�z�����R�-��&� ���������"�4�F� X�j�|ߎߠ߲�������������PREGn�W���0�~��� ����������� �2� D�V�h�z���������~$�$ARG_~@�D ?	����� � 	$$	[]�$:	���SBN_CONF�IG�XW�qRCII_SAVE  $zm���TCELLSE�TUP 
%�  OME_IO�$$%MOV_qH� ��REP���#��UTOBAC�K� 	t�FRA:\D� �.D�z '`��D�w� �s � 25/1�1/29 20:_26:16D�;�D���#//h�� C/j/|/�/�/�/�/D��X/�/??(?:?L? �/p?�?�?�?�?�?�? g? OO$O6OHOZO�? ~O�O�O�O�O�O�O��ׁ  c_F_\�ATBCKCTL.TM�)_;_M___\q_8INIm���j~CMESSA�G� �Qz �[ODGE_D� �j�X�O�p�_@PAUS�6` !� ,� 	�; ��v�>b����|_?�����?�ܾ0<�,		2aNijoTo �oxo�o�o�o�o�o�o B,Nxd`?TSK  mwxz�9UPDT�P�Wd�p�VXWZD_ENB�Tf
�v�STA�U�u��X�ISX UNT 2��vwy � 	 �ݟ���� �"���� �R� �0Q�D�R���k��5��U=��Z��<��Im������R�4E� [��L � ����w�X �9d����U�����4�MET��2�@��y PQ�B�lA�eA���B4M�B
6��B�w�>���>�@�? ��x?��?���v@q5�S�CRDCFG 1�Y �������%�7�I�pD�Q�	ܟ���� ��ϯ��Z��~�;� M�_�q�������6���FGR9��p�_ԳPkNA� 	FnѶ_ED�P1���� 
 �%-PEDT-¿ R�v���E�<�GE�
D�;9/�>���/  ����2��� ��B� ����{�����j�����3��#� �G� Y���G�ߠ�6�����a4�W������Z݀���Z�l������5 K��ߘ��Y�t���&�8���\���6��d ��Y�@����(��7�S0wY�@w��f���8����{�IZ��C/��2/���9{/��//LZݤ/?V/h/�/�/��CR���?�? Tn?�? ?2?�?V?԰~!�NO_DEL��ҲGE_UNUS�E޿дIGALL�OW 1� �  (*SY�STEM*��	�$SERV_GR�[�@`REG�Eq$�C���@NUM�J<�C�MPMU?@���LAYK���PMPAL�P>UCYC10 N3^�P!^YSULSU`_�M5Ra�CLo_��TBOXOR���CUR_�P�M�PMCNVV�P10I^�PT4D�LI�p�_�I	*P�ROGRA�DPG_MI!^Ko]`�AL+ejoTe]`B��o�N$FLUI_RESU9W�o�O��o�dMR�N�@�< �?�;M_q�� �������%� 7�I�[�m�������� Ǐُ����!�3�E��W�2BLAL_OU�T �K���W?D_ABOR:PcO���ITR_RTN�  �$�빸�N�ONSTO��� lHCCFS_U?TIL �̷�CC_AUXAX�IS 3$� �h}�j�|�����ƽCE_RIA_I`@��נ��F?CFG $�/�z#��_LIM�B�2+� �� �� 	��B\���$j� 
Ԡ��)�Z��%�/�����[������ ���!������L��(
5�����P}A�`GP 1H�����A�S�e�w�j6�CC� C7��UJ��]��p�����_�� C������U���������é�U̩�ձ�ߩ���������;���PC�k�����������*��������ɱ���������� D_� D!�!е!�!� ��&?��HE@ONFqIpC�G_P�P;1H� +EH� �ߟ߱����������C�KPAUS�Q1H�ף IR�S� H�A��e������ ��������E�+�i� {�a���A?Iץ��MؐNFO 1���� ��3��$:Ң �D/q�  D1>��4  ´J\�O� � ���LLECT_�!0�����EN+`㕸ʒ���NDE��#�/�12�34567890��"�A��/ҵHw��#)j��<i{ ��;��/��/ `/+/=/O/�/s/�/�/ �/�/�/�/8???'? �?K?]?o?�?�?�?�?�O�?��$� ���IO &��A▒O�O�Ol�O`GTR�2'DM�(��^�?�NN�(�oM Z��_MOR)q3)H��7ىU3� �Y�_�_�_�_�_�[bRT�kQ*H�,S�?<�<Ѡ<cz�KFd���%P,��;ϒo �o�o˿�o�oœh�U�A	@E�oA� �sja�P�DB.���4c?pmidbg3�L�Рs:��>uqpz|��v  ��>x��}.��}�l`��|�<�mgP���t��~f������>@ud1:�?���XqDEF -���zC)*�cO�b?uf.txtJ��|�K�[`�/DM��>����R�A��MC&iR20_{RCd���hS21����G�A�CzA�d4�EI��jA��	C-]��G/X"B�h�\F]�H�j��D��GF�1�J��iF���I؂�L���YHe4�JN��N��mJ���MSo��A����f23DLD(�	>z�!� 2��}�k�yc
�@x9�&) C��e Da I��E���  E�%q�F�� E�p�u�F�P� E��fF�3H ��G�M��Ъ5�>�33���?�xn9�q@��Q5����RpA�?aA=L��<#�QU�@,�Cϒ����RSMOFST� +i�����P_�T1Ɠ4DMA �=ք�MODE 5dm�@��	Q�i�;��%��?����<�M>�{�Ͷ�TESTc�)2i�`�R�6�O�DK�|AB�An� 8���\�n�CdB�j��Cu @p������p:d�QS ����(������4�IJ7>���>B8m�5$�RT_c�P�ROG %j%�d�1�h@NUSE�R��x�KEY_T�BL  e������	
��� !"#$%&'�()*+,-./�(:;<=>?@�ABCc�GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������>��͓���������������������������������耇���������������������9�4A8�LCK��F�<y��STAT��2�=X�_ALM������_AUTO_D�O�E�FDRw 3:i�2h&q�[~�� B�UOSYST-3�22 Auto �status c�heck tim?e out ������$TELE�O8��� ���)qA�ʜ@��������?��ڛMsB��õ�?*?���?Mf=���o�TR���-���D.��B���C����B�N�*p�4m�N4�J5HjC5H��>���BJ��d�BF��pZ��[~�bbt�����5/�M*F�B��GA+$����@R��J��}BQ�H�����������2>��@ǿ@���&��CBxHCK?H<B��6>T�bt��/��u�U S�H?Z?l?��$7?�? :�� mϸ?�?p���? �?OO�?,OfOxO�M 6?�O�O�O~?�O	_�? *_$_BOD_6_p_~_T_ �_�_�_�_�Oo)o;o �OLoqo_�o�o�_�o �o�o�o�o�oFX o��No���o ����@�N�$� b�x�����n���� ��A��b�\�z�|� n�������ʟ���(� ֏O�a�s������T� ʯį��֯���� 2�H�~���>���ɿۿ ���ϼ�2�,�J�L� >�xφ�\Ϛϰ����� ���1�C��T�y�$� �ߔ߲ϴߦ������� ��N�`�߇��� V߼��������� �H�V�,�j������� v�����$I�� jd���v��� ��0��Wi{ &��\���� �/&/�:/P/�/�/ F�/�/�/��/?� :?4?R/T?F?�?�?d? �?�?�? O�/'O9OKO �/\O�O,?�O�O�?�O �O�O�O�O
_ _V_h_ O�_�_�_^O�_�_�O 
oo"_$ooPo^o4o ro�o�o�o~_�o	 �_,Q�_rl�o� ~�����&�8� �o_�q���.����d ڏԏ��� �.�� B�X�����N�ǟٟ� ����!�̏B�<�Z�\� N�����l�������� ��/�A�S���d���4� ����¯Ŀ�����Կ �(�^�p���ϩϻ� f����Ϝ���*�,� �X�f�<�zߐ����� �����#���4�Y�� z�t�ߔ������� ����.�@���g�y��� 6����l��������� ��(6J`�� V������)�� JDbdV��t ���/�7/I/[/ l/�/<�/�/��/ �/�/?�/?0?f?x? &/�?�?�?n/�?�?�/ OO2?4O&O`OnODO �O�O�O�O�?__+_ �?<_a_O�_|_�O�_ �_�_�_�_�_ o6oHo �Ooo�o�o>_�o�ot_ �o�oo�o0> Rh��^o��� �o�1��oR�L�jl� ^�����|���Џ�� �?�Q�c��t���D� ����ҏԟƟ ��� "�8�n���.�����˯ v�ܯ���"��:�<� .�h�v�L�����ֿ� ���!�3�ޯD�i�� �τϢ��ϖ����ϴ� ���>�P���w߉ߛ� FϬ���|�����
�� ��8�F��Z�p��� f���������9��� Z�T�r�t�f������� ���� ��GYk �|�L������ ��*@v� 6���~�	/� */$/BD/6/p/~/T/ �/�/�/�/�?)?;? �L?q?/�?�?�/�? �?�?�?�?�?OFOXO ?O�O�ON?�O�O�? �O�OO__@_N_$_ b_x_�_�_nO�_�_o �OoAo�Obo\oz_|o no�o�o�o�o�o( �_Oaso��To ���o����� 2�H�~���>��ɏۏ ����2�,�J�L� >�x���\�������� ���1�C��T�y�$� ������������į ��N�`�������� V���ῌ������ �H�V�,�jπ϶��� v����߾�$�I��� j�d߂τ�v߰߾ߔ� �����0���W�i�{� &ߌ��\��������� ���&���:�P����� F������������ :4R�TF��d ��� ��'9K ��\�,���� ����
/ /V/h/ �/�/�/^�/�/� 
??"/$??P?^?4? r?�?�?�?~/�?	OO �/,OQO�/rOlO�?�O ~O�O�O�O�O�O&_8_ �?__q_�_.O�_�_dO �_�_�O�_�_ o.oo�BoXo�otc�$CR�_FDR_CFG� ;re��Q
UD1:��W�P�aJ�d  ��`�\�bHIST �3<rf  �` � ?�R�@tAtB�bUC�PCpDtEtUItg�Ppot�w�_��bINDT�_EN6p�T��q�bT1?_DO  �U�u�sT2��wVAR� 2=�gp �hq  �m��m��R�n�44�n4�m[��RZ��`STOP��rT�RL_DELET�Np�t ��_SCREEN re~�rkcsc�r�Uw�MMENU �1>��  <�\%�_��T�� R��S/�U���e�w�ğ ������џ�	�B�� +�x�O�a��������� ��ͯ߯,���b�9� K�q�������࿷�ɿ ����%�^�5�Gϔ� k�}��ϡϳ������ ��H��1�~�U�gߍ� �ߝ߯�������2�	� �A�z�Q�c���� �������.���d� ;�M���q�������������YӃ_MAN�UAL{��rZCDƳa?�y�rG +���R�f"
�^"
?|(��PdT�GRP 2@�y��B� � s���� �$DBCO�pRIG���v��G_ERRLOG' A��Q�I�[m �NUM�LIM�s��u
��PXWORK 1B�8����//�}DBTB_�� C%����S"� �aDB_A�WAY��QGC;P �r=�ןm"G_AL�F�_��Yz����p�vk  �1D� , 
���/"�/%?/(_Mؘpqw,@�=5ON�TIM����t��_6�)
�0�'MOTNENFpF�;�RECORD 2�J� �-?�SG�O��1�?"x"!O 3OEOWO�8_O�O�?�O O�O�O�O�O�O(_�O L_�Op_�_�_�_A_�_ 9_�_]_o$o6oHo�_ lo�_�o�_�o�o�o�o Yo}o2�oVhz ��o��C�
� �.��R��K���� ����Џ?��ߏ�*� ����+�b�t�㏘��� ��Ο=�O�����:� %���p�ߟ񟦯��O� ǯ�]������H�Z� ��������#�5�����ϩ�i"TOLEoRENCK4Bȿ"� L��� CSS�_CCSCB 2%K�\0"?" {ϰϟ���7��
�� ��@�R�d�3߈ߚ�"�x���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg0y��� ���d���R�LL]��La�m1T#2 7C�C��F\�^ A�C�pC�ɴ�#�0� 	� A���B<���?�  �$�0���\0袰�0��B��`#s�K/]/(o/�ϓ/�/�/�s/�/�/�K�K8�Lg��Ҡ\�1� 1�3�OȦ��/��/T`?;�@��O? �?�?�?Ȏ0AF��?{F�A OO�7�1 ���9M	AB
AZO dBAE�9$O�O�O�Oi:�P��`�@0�DzJCA� @��
X-.
[h=��	 M?�>O�ڴ�q_@�_�_�_:W�A<o :[<ǲ/o�/�_�+oPoboto�eAC�HC�V�WB$�Dz�cD�`�a=/�o�o o�oW�a.+!��2=t,y�J?�.s�s �js�w�yj���@����Q�Qs�@ `��$�����A���� Bމ�o��'�9��_ ]�o�N���r���ɟ۟ _�B�ʄ��YZ>`�+�ۘBό�B�e@���@B뻷��@�Z�l�~���� `_м¯���
���̯ 9�,�]�o��� �H��� ��ٿ뿊��ƿ3�E� W�iϬ���$ϱ�����  Ϟ����/�A�S߶� w�V�h߭ߌ��S������_�f	��H� ?�Q�~�u����� �������D��-� g�q������������� 
@7Icmp��߾�  � ����)M@q dv������ �//I/P�m/�v/ �/�/�/�/�/�/�/? 3?*?<?i?`?r?�?^/ �?�?�?�?�?O/O&O 8OJO\O�O�O�O�O�O��O�O�g	  VQ�P�s �]PC4p*p�p6U6P\C9:p/p�� ]V^P*M]�6P�:P�>P�VVJ_�^P�bP�fP��Vr]v���p Q
@k���_oo�id1Q&oNo ;o_co�o<ˏUUA   �o�k1Q@�  �o�k�b������P�p �� 1��6��1C���C�cPfL���?#�c>�{�e��`�cP�@@�dX��r�`B�cP>�sv�qC��p����b��t<�o?�PH�)S�B�t`q�q�p�r�`B����eIC�&�Q�4( ��oz�UU*�� ����9�Y=��@@����4Q��-RBQ�[��K$�7��BQ��Y�b��`ځ` � ?�p���U�[?����}t��$����$DCSS_CL�LB2 2M���p�P�^?�NSTCY 2N����  �������ʟ؟� ��� �2�D�Z�h�z� ������¯ԯ��SA��DEVICE 2%O��!�$��4& V�h�������˿¿Կ ���
�7�.�[�R�π�ϣϵ�����4(A�HNDGD P���*�Cz�A�LS 2Q��_�Q�c�u���ߙ߽߫���?�PA?RAM RP���1�`�&�RBT 2}T�� 8�P	<C�'pÀ�pi�l��s@"�R��(qI�ʹX��0�pB CW  ��B\x�N���Z����%��)� ��X�j��p����zq��I���B �(s,�F� �p�V��q���b��B ��4&c �S�e� l�4+����H1~ޡ���D�C��$Z��b���A�,� 4�u@�X�@��^@w����]B���B��cP%��C4��C3:^C4��nЬ ��p8�-�B{B���A���� l���C�C3��JC4jC3���yn+�3 Dff 2�A PB W4+@:�]o�W �����/�/ P/'/9/K/]/o/�/�/ �/�/?�/�/�/?#? 5?�?Y?k?�?�?�o�? �?O�?6O!OZOlOWO �O�Es�?�?�?�O�O _�O�OL_#_5_G_Y_ k_}_�_�_�_ o�_�_ �_oo1o~oUogo�o �o�o�o�owO D /Aze����O �o�o
��o��R�)� ;���_�q��������� �ݏ�<��%�r�I� [�m��������ǟٟ &�8��\�G���k��� ����گů����� F��/�A�S�e�w�Ŀ ������ѿ����� +�x�O�aϮυϗϩ� ������,���b�t� ﯘ߃߼ߧ������ ���:��C�U߂�Y� k����������� 6���l�C�U�g�y� ���������� ��	 -?Q���� ���@+d vQ������ ��*///%/r/I/ [/�//�/�/�/�/�/ &?�/?\?3?E?�?i? {?�?�?U�?�?"O4O OXOCO|OgO�O{� �?�O�?�O�O0___ f_=_O_a_s_�_�_�_ �_�_o�_oo'o9o Ko�ooo�o�o�o�o�o �O:%^I�������H�$D�CSS_SLAV�E U����	���z_�4D  	��A�R_MENU V	� �j�|�������ď�BY�� ��~�?�SHOW 2W>	� � �b�a G�Q�X�v��������� П֏���� @�:� d�a�s���������� ߯��*�$�N�K�]� o�������̯ɿۿ� ��8�5�G�Y�k�}� �϶�����������"� �1�C�U�g�yߠϝ� ���������	��-� ?�Q�c��s����� ��������)�;�M� t�������������� ��%7Ip�m ���������� !3ZWi�� �J����// DA/S/e/��/��/ �/�/�/�/?./+?=? O?v/p?�/�?�?�?�? �?�??O'O9O`?ZO �?�O�O�O�O�O�OO �O_#_JOD_nOk_}_ �_�_�_�_�O�_�_o 4_.oX_Uogoyo�o�o �o�_�o�o�ooBo ?Qcu���o:����CFG MX)�3�3q5p��FRA:\�!�L+�%04d.WCSV|	p}�� �qA g�CHo�zv�	����3q�����́܏� �|��4��JP�����qp1� �R�C_OUT Y���C��_�C_FSI ?~i� .� ������͟����� >�9�K�]��������� ίɯۯ���#�5� ^�Y�k�}�������ſ �����6�1�C�U� ~�yϋϝ��������� �	��-�V�Q�c�u� �ߙ߽߫�������� .�)�;�M�v�q��� ����������%� N�I�[�m��������� ��������&!3E ni{����� ��FASe �������� //+/=/f/a/s/�/ �/�/�/�/�/�/?? >?9?K?]?�?�?�?�? �?�?�?�?OO#O5O ^OYOkO}O�O�O�O�O �O�O�O_6_1_C_U_ ~_y_�_�_�_�_�_�_ o	oo-oVoQocouo �o�o�o�o�o�o�o .);Mvq�� �������%� N�I�[�m��������� ޏُ���&�!�3�E� n�i�{�������ß՟ ������F�A�S�e� ��������֯ѯ��� ��+�=�f�a�s��� ������Ϳ����� >�9�K�]φρϓϥ� ����������#�5� ^�Y�k�}ߦߡ߳��� �������6�1�C�U� ~�y����������� �	��-�V�Q�c�u� �������������� .);Mvq�� ����% NI[m���� ����&/!/3/E/ n/i/{/�/�/�/�/�/��/�/3�$DCS�_C_FSO ?����71 P ? ?T?}?x?�?�?�?�? �?�?OOO,OUOPO bOtO�O�O�O�O�O�O �O_-_(_:_L_u_p_ �_�_�_�_�_�_o o o$oMoHoZolo�o�o �o�o�o�o�o�o%  2Dmhz��� ����
��E�@� R�d���������ՏЏ ����*�<�e�`� r���������̟��� ��=�8�J�\�����|��?C_RPI4>F?�������3?��&�o����� >SLү@d������%� 7�`�[�m�Ϩϣϵ� ���������8�3�E� W߀�{ߍߟ������� �����/�X�S�e� w����������� �0�+�=�O�x�s��� ���������� 'PK]o��� �����(#5 Gpk}����� Q���/6/1/C/U/ ~/y/�/�/�/�/�/�/ ?	??-?V?Q?c?u? �?�?�?�?�?�?�?O .O)O;OMOvOqO�O�O �O�O�O�O___%_ N_I_[_m_�_�_�_�_ �_�_�_�_&o!o3oEo noio{o�o�o�o�o�o �o�oFASe�������>�N�OCODE Z�U��?�P�RE_CHK �\U��pA �p?�< ��pU�x]�o�U� 	 <Q� �������ۏ�Ǐ� #����Y�k�E����� {�şן��ß���� C�U�/�y�����s��� ӯm���	���?�� +�u���a�������ɿ �Ϳ߿)�;��_�q� K�}ϧϝ������ω� ��%����[�m�Gߑ� ��}߯��߳����!� ��E�W�1�c��g�y� ������������A� S�-�w���c������� ������+=a sM_����� �'�]o	 ������/ #/�G/Y/3/e/�/i/ {/�/�/�/�/?�/? C?9Ky?�?%?�?�? �?�?�?	O�?-O?OO KOuOOOaO�O�O�O�O �O�O�O)_____q_ K_�_�_a?�_�_�_�_ o%o�_Io[o5oGo�o �o}o�o�o�o�o�o �oEW1{�g� ��_����/�A� �M�w�Q�c������� ���Ϗ�+���a� s�M���������ߟ� ��'���3�]�7�I� �����ɯۯ���� ���G�Y�3�}���i� ��ſ��������1� C���+�yϋ�eϯ��� ����������-�?�� c�u�Oߙ߫߅ߗ��� �����)��M�_�U� G���A�������� �����I�[�5���� k������������� 3EQ{q�� �]����/A ewQ���� ���/+//7/a/ ;/M/�/�/�/�/�/� �/?'??K?]?7?�? �?m??�?�?�?�?O �?5OGO!O3O}O�OiO �O�O�O�O�O�/�O1_ C_�Og_y_S_�_�_�_ �_�_�_�_o-oo9o co=oOo�o�o�o�o�o �o�o__M_�o k�o����� ���I�#�5���� k���Ǐ��ӏ��׏� 3�E��i�{�5c��� ß�����ӟ�/�	� �e�w�Q�������ѯ 㯽�ϯ�+��O�a� ;��������Ϳ߿y� ���!�K�%�7ρ� ��mϷ��ϣ������� ��5�G�!�k�}�W߉� �ߩ������ߕ��1� ��g�y�S���� ��������-��Q� c�=�o���s������� ������M_9 ��o���� �7I#mY k������!/ 3/)/i/{//�/�/ �/�/�/�/�/?/?	? S?e???q?�?u?�?�? �?�?OO�?%OOOE/ W/�O�O1O�O�O�O�O __�O9_K_%_W_�_ [_m_�_�_�_�_�_�_ o5oo!oko}oWo�o �omO�o�o�o�o1 UgAS��� ���	����Q� c�=�����s���Ϗ�o ������;�M�'�Y� ��]�o���˟���� ۟�7��#�m��Y� �����������!� 3�ͯ?�i�C�U����� ��տ�������	� S�e�?ωϛ�uϧ����Ͻ������$�DCS_SGN �]	�E��-����01-D�EC-25 13�:03 ��2�9-NOVV�20�:27_�x�x�� [}�t��q��т�xҚك�JѨ��EƼÞ� �ۈǖ�  1�HO�W ^	�� x�/�VE�RSION �=�V4.5.�2��EFLOGI�C 1_���  	�����C���R�%�PROG_E_NB  ��:��{�s�ULSE  �X��%�_AC�CLIM������d��WRSTgJNT��E��-�EMO|�zя�$���INIT `2�����OPT_S�L ?		�	�
 	R575��V]�74b�6c�7c�50��1���C��|�@�TO  L��� �V�DEXҞ�dE�x�PA�TH A=�A�\k}��HCP�_CLNTID y?�:� D���ռ��IAG_G�RP 2e	�����z�	 �@�  
ff�?aG���BG�  2��/�8�[I@c�ς!��7@�z�@^��@
�!���mp2m15 �89012345�67���� � ?��?��=q?��
?���R?�Q�?ѯ�?�����?(�?�z����x�@�  A_�A�p !7A�8�8_�B4�� ��L�x�
�@����@��\@~��R@xQ�@q���@j�H@c��
@\��@U�@Mp��//�'$�; �O)H���@Ct >d 9���@4�/\)@)�� #t {@��/�/�/�/�/P'�?���?����_ ?}p�?u?n{?s ;?\�Q�? ?�2?D?V?h8�
=?�����0w5�z��H?p�h��?^�R�?�?�?�?��?h8��t0����@�?��0� ;@&O8OJO\OnOP' �$_�_Y_k_�O?_ �_�_�_�_�_s_�_�_ 1oCo!ogoyoo�o���Bj"� �2{1�@"?���f�t0�d"�5!�
u4V��u"�B3t�A>u��U?@[q��@`,�=q�=b���=�E1>�J��>�n�>��H�"<�o �z�s��q��� �x�C��@<(�Uz� �4�� ����A@x�?*�o��m*� P�b���tn���2����Ώ�����i>J���&�bN2�"�'�G�N��o@�@v�奈0����@f�fr!l ��33����(��"C��� ƒI�CH��)C.dB؃�"8"����' ���"~�A?�&"K���,�pf�B��@�p��������p���������ƥx�D/  ��1����������3��N�T���
�C+ �o#����� ȿ���׿����?,��<�o��CT_C�ONFIG f���|�e�gY��STBF_TTS��
�������}���1�MAU�������MSW_C5F��g�  # �ڿOCVIEW��h!�-���s߅� �ߩ߻��ߟ�a���� �,�>�P���t��� �����]�����(� :�L�^���������� ����k� $6H Z��~����� �y 2DVh �������v�KRC�i���!� ��/S/B/w/f/�/�/��/��SBL_FA?ULT j*6�>�!GPMSK���'���TDIAG ik��-�������UD1: 6�78901234A5I2��=1�Ǥ�P\� �?�?�?�?�?�?�?O O'O9OKO]OoO�O�O �Od696���r
t?�O>|�TRECP"?4:
B44_[7��s?p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�O��O�O�o7�UMP__OPTIO=��.F�aTR����)u�PME��Y_T�EMP  ÈW�3BC�gp�B�QtUNI����gq��YN_BRK �lL�7�EDITO�R�a�a@�r_
PE�NT 1m) � ,&TEL�EO[p���&?SET_WCp,�|�l�pPSNAP^P|X�?�MTPG�p W�i��/��IĦ��ʏ ���=�$�a�H��� ��~�����ߟ�؟� ��9� �2�o�V���z� ��ɯ���ԯ�#�
��G�DɴpMGDI_�STAzuV�gq�uN�C_INFO 1yn!��b���X�`��������n�1o!ۇ ��o����
�d�oU�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫� �� u����
��*�B� *�P�b�t����� ��������(�:�L� ^�p���������2��� ����9�CUg y������� 	-?Qcu� �������// 1;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�?� �?�?�?O)/OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_ �_�_�_�?�?�_�_o �_3O=oOoaoso�o�o �o�o�o�o�o' 9K]o����_ �_����+o5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y��������ӟ��� 	�#�-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ����7� I�[�m�ϑϣϵ��� �������!�3�E�W� i�{ߍߟ߹������� ���%�/�A�S�e�w� ������������ �+�=�O�a�s����� �����������' 9K]o���� ����#5G Yk}�	���� ��/1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?��?�?�?�?/O )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�?�_�_ �_�_O�_!o3oEoWo io{o�o�o�o�o�o�o �o/ASew ��_�_����o �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o������� ɟ۟���#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߝ��� �����������%�7� I�[�m������� �������!�3�E�W� i�{��߇��������� �/ASew ������� +=Oas���� ������//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/?#?5?G? Y?k?���?�?�?�? ��?OO1OCOUOgO yO�O�O�O�O�O�O�O 	__-_?_Q_c_u_�? �_�_�_�_�?�_oo )o;oMo_oqo�o�o�o �o�o�o�o%7 I[m�_u��� �_���!�3�E�W� i�{�������ÏՏ� ����/�A�S�e� �������u����� �+�=�O�a�s����� ����ͯ߯���'� 9�K�]�w��������� ɿ�����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� ���ߝ߯���ۿ���� 	��-�?�Q�c�u�� ������������ )�;�M�_�y߃����� ��������%7 I[m���� ���!3EW q�c�������� �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?i{�?�? �?�?��?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ �?s?}_�_�_�_�?�_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	-?Qk_u� ���_����� )�;�M�_�q������� ��ˏݏ���%�7� I�cQ��������� ٟ����!�3�E�W� i�{�������ïկ������/�A�[� ��$ENETMOD�E 1p����  k��k�f�����j�OATCFG q��/��Ѵ���C���DATA �1rw�Ӱ���*	�*��'�9�K�D]�l�dlύ�e� �ϻ���������'� �ϳ�]�o߁ߓߥ߷� 1���U����#�5�G� Y����ߏ������� ����u��1�C�U�g� y������)������� 	-����cu������j�RPO_ST_LO��t�[
׶#5Gi�RROR_PR� �%w�%L�XTABLE  w��ȟ����RSEV_NUM ��  ����  �_AUTO_?ENB  ����X_NO5! u�w���"  *U�x �x �x �x �+ +w �/�/�/Q$F�LTR=/O&HIS�#]�J+_ALMw 1vw� �[x,e�+�/Q?c? u?�?�?�?�/_"W   w�v!���:�j�TCP_VER� !w�!x�?$�EXT� _REQ��&�H)BCSIZ\KO=DSTKhIf%��?BTOL  �]Dz�"�A= =D_BWD�0�@��&�A���CDI�A �wķ���]�KS�TEP�O�Oj�PO�P_DO�Oh�FD�R_GRP 1xw��!d 	�?�_���yPs�Y�Q'��M"����l��T� �����VyS�_�]yPA�8��B5�A��
�A1)l@?���A��
�T�A��@՚�o@�d�bqn�@ oGo�_Wo}oho�o�o��om?�L%@&���?��?o�"�n
 L��*v b�`]@8> J@!�4:�o^I���Y@`�t@S33�u�]@�q�g��yPF@ ��|yP�G�  @�Fg��fC�8RL��]?��`i��~6�X�����875t���5���5`+�����/OFEATU�RE y���@���Hand�lingTool� �]Eng�lish Dictionary��4D St��ar�d��Analo�g I/O>�G�g�le Shift�Z�uto Sof�tware Up�date�mat�ic Backu�p���groun?d Edit ���CameraU�F�Y�CnrRndI�m���ommon� calib U�I��nˑ�Mo�nitor$�tr~�Reliabn���DHCP �[�a�ta Acqui�s3�\�iagno�s��R�v�ispl�ayΑLicen�sZ�`�ocume�nt Viewe�?�^�ual Ch�eck Safe�ty��hanc�ed���s�F�rܐ�xt. D7IO /�fi��@�wend�Err>�QL��\�4�s[�rP��K� �@
�FCTN_ Menu��vZ����TP In��f�acĵ�GigE�־�Đp Mas_k Exc�g=��HT԰Proxy� Sv��igh�-Spe�Ski��� Ť�O�mmun�ic��onsV�u�r����q�V�ײconnect 2���ncrְstruH!��ʴ�eۡ��J���X�KAREL C�md. L�ua����Run-Ti�<�Env�Ȟ�el� +��s��S/W��ƥ���r�Boo�k(System�)
�MACROs�,M�/Offse�u�p�HO���o�u�M�R8�4���Mech/Stop+�t����"p�im�q���x�R�쪐��odo�wit#ch�ӟ�.��4�OptmF��,�f�il䬳�g��p�ulti-T�Γ�PCM fun��¼�o��������Re�gie�rq���ri�ݠF���S�Num� Sel��/�:� Adjua�*�W�q�h�tatu��ߪ��RDM Rob�ot�scove�'���ea��<�Freq Anlyq�'Rem��O�n5���>��ServoO�!�~�SNPX b-�vv�SN԰Cliܡ<?r�Libr&�_��� ��q +oJ�t��ssag��X�@a ����	�@/Iս>�MILIB��?P Firm����P��AccŐ͛T�PTXk��eln���������or�quo�imulah=��|u(�Pa&���ĐX�B�&+�ev�.���ri��T�USB port- �iPf�aݠ&?R EVNT� nexcept�`����%5��VC�rl�c���V���"h�%q�+SR SCN��/SGE�/�%UI~	�Web Pl�� >��A43��ۡ���ZDT Applxj�
�{1EOAT�౔�&0?�7Gri�d�񾡬=�?iR��".5� F���/גR�X-10iA/L��?Alarm C�ause/��ed�(�All Smo�oth5���C�sc�ii+�V�Load�䠌JUpl�@w�t�oS ��rity�AvoidM(�sb7�t�@�ycn�`����_�CS+����. c��XJo ���-T3_H�.RX���U���Xcolla3bo����RA�:�.9D��in���gNRTHI
�On��e Hel����ֿ������1trU�R?OS Eth$��A@������;,�G �B�,|HUpV�%�fW�t ԰�_iRS��ݐ�64MB D�RAM�o�cFROp���L8F FlD������2M �A:�op�m�ԕex@V�
�sh��q��wce�u��p,��|tyn�sA�
��%�r����J��^�.v� P)Q/sbS�`�p��O�N��mai���U���R�q�T�1�^FC+Ԍ%̋F�s9�ˌk̋��Ty-p߽FC%�hױV�:N Sp�ForްK��Ԭ�lu!����cp�OPG j�֡�RJ:�[L`Sup"}�0�֐f��crFP��3lu� ��al�����r��i�
q�4�@а�uest,IMPLE ׀6*�|HZ���c0�BTe�a(�|���$rtu8���V�9HMI�¤���UIFc�pono2D�BC�:�L�y� p���������ʿܿ	�  ��?�6�H�u�l�~� �Ϣϴ��������� ;�2�D�q�h�zߧߞ� ���������
�7�.� @�m�d�v����� �������3�*�<�i� `�r������������� ��/&8e\n �������� +"4aXj�� ������'// 0/]/T/f/�/�/�/�/ �/�/�/�/#??,?Y? P?b?�?�?�?�?�?�? �?�?OO(OUOLO^O �O�O�O�O�O�O�O�O __$_Q_H_Z_�_~_ �_�_�_�_�_�_oo  oMoDoVo�ozo�o�o �o�o�o�o
I @Rv���� �����E�<�N� {�r�������Տ̏ޏ ���A�8�J�w�n� ������џȟڟ��� �=�4�F�s�j�|��� ��ͯį֯����9� 0�B�o�f�x�����ɿ ��ҿ�����5�,�>� k�b�tφϘ��ϼ��� �����1�(�:�g�^� p߂ߔ��߸�������  �-�$�6�c�Z�l�~� ������������)�  �2�_�V�h�z����� ����������%. [Rdv���� ���!*WN `r������ �//&/S/J/\/n/ �/�/�/�/�/�/�/? ?"?O?F?X?j?|?�? �?�?�?�?�?OOO KOBOTOfOxO�O�O�O �O�O�O___G_>_ P_b_t_�_�_�_�_�_ �_oooCo:oLo^o po�o�o�o�o�o�o	  ?6HZl� �������� ;�2�D�V�h������� ˏԏ���
�7�.� @�R�d�������ǟ�� П�����3�*�<�N� `�������ï��̯�� ��/�&�8�J�\��� ��������ȿ����� +�"�4�F�Xυ�|ώ� �ϲ���������'�� 0�B�T߁�xߊ߷߮� ��������#��,�>� P�}�t������� ������(�:�L�y� p��������������� $6Hul~�����  H552�v�21R78{50J614�ATUP'545z'6VCAMwCRIbUIF'�28cNRE5�2VR63SC�HLIC�DO�CV�CSU8�69'02EIOuC�4R69V�ESET?UJ7�UR68MAS�KPRXY{7.OCO#(3?�+ &3j&J6%5u3�H�(LCHR&�OPLG?0�&M�HCRS&S�'MC�S>0.'552MgDSW+7u'OPu'GMPRv&��(0&7PCMzR0q7+ �2� �'51J51��80JPRS"'6�9j&FRDbFR�EQMCN9=3&SNBA��'/SHLBFM1G��82&HTC>T�MIL�TPA��TPTXcFEL�F� �8J�95�TUTv'9�5j&UEV"&UE�CR&UFRbVCuC
XO�&VIPnFwCSC�FCSG���IWEB>HTT>R6��H;�RVCGiWIGQWI�PGS�VRCnFD�Gu'H7�7R66�J5'R�8R5U1
(6�(2�(5VR�J8�86�L=Ih% �84g662wR64NVD"&�R6�'R84�g7�9�(4�S5i'J[76j&D0�gF x�RTSFCR�gC;RXv&CLIZ8I�CMS�Sp>STuYnG6)7CTO>���7�NNj&O�RS�&C &FCBn�FCF�7CH>wFCR"&FCI�VKFC�'J�PO7GBf�M�8OLaxENDvS&LU�&CPR�7ULWS�xC�STx�TE�gS60F�VR�IN�7IH aF�я�����+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi{ ������� /ASew�� �����//+/ =/O/a/s/�/�/�/�/ �/�/�/??'?9?K? ]?o?�?�?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_ �_�_�_�_�_�_	oo -o?oQocouo�o�o�o �o�o�o�o); M_q����� ����%�7�I�[� m��������Ǐُ��  H5�52��21�R�78�50�J6{14�ATUP7��5457�6�VC�AM�CRI��U�IF7�28��NR�E�52v�R63��SCH�LIC�ƚDOCV�CS]U�8697�0F��EIOCǛ4�R{69v�ESETW�vu�J7u�R68��MASK�PRXuY��7�OCO���3W����6�3�J�65�536�H$�L{CHƪOPLGW��0�MHCRǪS���MCSV�0��5=5F�MDSW���;OP��MPR��㐺6�06�PCM��R�0E˓�F���6�51�f�51��0f�PR�S��69�FRDކ�FREQ�MC�N�936�SNByAכ%�SHLB��ME��ּ26�HT=CV�TMIL�6��TPAV�TPTXF��ELړ�6�8%��#��J95��TU�T��95�UEVUECƪUFR���VCCf�O��V�IP��CSC��C�SGƚ$�I�WE�BV�HTTV�R6�՜��S���CG��I�G��IPGS'�RmC��DG��H7�˗R66f�5�u�R���R51f�6�2��5v�#�J׼��6B��LU�5�s�v�4���66F�R64�N�VD��R6��R8�4�79�4��S�5�J76�D0�uFRTS&�C�R�CRX��CL9I&�e�CMSV�s�V�STY��6�C�TOV�#�V�75�NN�ORS����6�wFCBV�FCF�˻CHV�FCR��F[CIF�FC��J#�j�G
M��OL��ENDǪLU��C�PR��Lu�S�C�$�StTE�S6�0�FVRV�IN��IH���m??�? �?�?�?�?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_e_w_�_�_�_�_�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9K]o� �������� #�5�G�Y�k�}����� ��ŏ׏�����1� C�U�g�y��������� ӟ���	��-�?�Q� c�u���������ϯ� ���)�;�M�_�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�e�w������� ������+�=�O�a� s��������������� '9K]o� ������� #5GYk}�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a��s���������͏ߏ��STD�LANG��� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ�ܰ���RBT
�OPTN������'�9� K�]�o�����������DPN	��� )�;�M�_�q������� ��������%7 I[m���� ����!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O �O�O�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o	-?Qcu �������� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ �����/�A�S�e� w���������ѿ��� ��+�=�O�a�sυ� �ϩϻ��������� '�9�K�]�o߁ߓߥ� �����������#�5� G�Y�k�}������ ��������1�C�U� g�y����������������	-?Qc��f�������99��$FEA�T_ADD ?	����  	�#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ���������DEMO y~   � L�B�T߁�xߊ߷߮� ����������G�>� P�}�t������� ������C�:�L�y� p��������������� ?6Hul~ ������ ;2Dqhz�� ���� /
/7/./ @/m/d/v/�/�/�/�/ �/�/�/?3?*?<?i? `?r?�?�?�?�?�?�? �?O/O&O8OeO\OnO �O�O�O�O�O�O�O�O +_"_4_a_X_j_�_�_ �_�_�_�_�_�_'oo 0o]oTofo�o�o�o�o �o�o�o�o#,Y Pb������ ����(�U�L�^� ����������ʏ�� ��$�Q�H�Z���~� ������Ɵ�����  �M�D�V���z����� ��¯ܯ��
��I� @�R��v��������� ؿ����E�<�N� {�rτϱϨϺ����� ���A�8�J�w�n� �߭ߤ߶�������� �=�4�F�s�j�|�� �����������9� 0�B�o�f�x������� ��������5,> kbt����� ��1(:g^ p�������  /-/$/6/c/Z/l/�/ �/�/�/�/�/�/�/)?  ?2?_?V?h?�?�?�? �?�?�?�?�?%OO.O [OROdO�O�O�O�O�O �O�O�O!__*_W_N_ `_�_�_�_�_�_�_�_ �_oo&oSoJo\o�o �o�o�o�o�o�o�o "OFX�|� �������� K�B�T���x������� ۏҏ����G�>� P�}�t�������ןΟ �����C�:�L�y� p�������ӯʯܯ	�  ��?�6�H�u�l�~� ����Ͽƿؿ���� ;�2�D�q�h�zϔϞ� ���������
�7�.� @�m�d�vߐߚ��߾� �������3�*�<�i� `�r���������� ���/�&�8�e�\�n� ���������������� +"4aXj�� ������' 0]Tf���� ����#//,/Y/ P/b/|/�/�/�/�/�/ �/�/??(?U?L?^? x?�?�?�?�?�?�?�? OO$OQOHOZOtO~O �O�O�O�O�O�O__  _M_D_V_p_z_�_�_ �_�_�_�_o
ooIo @oRolovo�o�o�o�o �o�oE<N hr������ ���A�8�J�d�n� ������яȏڏ��� �=�4�F�`�j����� ��͟ğ֟����9� 0�B�\�f�������ɯ ��ү�����5�,�>� X�b�������ſ��ο ����1�(�:�T�^� �ςϔ��ϸ�������  �-�$�6�P�Z߇�~� �߽ߴ���������)�  �2�L�V��z��� ����������%��.� H�R��v��������� ������!*DN {r������ �&@Jwn �������/ /"/</F/s/j/|/�/ �/�/�/�/�/??? 8?B?o?f?x?�?�?�? �?�?�?OOO4O>O kObOtO�O�O�O�O�O��O__0]  'XF_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o�o "4FXj|�� �������0� B�T�f�x��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰπ��������
��.�  /�)�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ���(:L ^p������ � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?V?h?z?�? �?�?�?�?�?�?
OO .O@OROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo\o no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x����� ����ҏ�����,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� ������&�8�J�\� n��������������� ��"4FXj| ������� 0BTfx�� �����//,/ >/P/b/t/�/�/�/�/ �/�/�/??(?:?L? ^?p?�?�?�?�?�?�? �? OO$O6OHOZOlO ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_ �_�_�_�_�_�_
oo .o@oRodovo�o�o�o �o�o�o�o*< N`r����� ����&�8�J�\� n���������ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T�f�x����� ����ү�����,� >�P�b�t��������� ο����(�:�L� ^�pςϔϦϸ����Ϡ�� ��$�4�8� +�N�`�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�o�o �o�o�o&8J \n������ ���"�4�F�X�j� |�������ď֏��� ��0�B�T�f�x��� ������ҟ����� ,�>�P�b�t������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��� �2�D�V�h�z� �ߞ߰���������
� �.�@�R�d�v��� �����������*� <�N�`�r��������� ������&8J \n������ ��"4FXj |������� //0/B/T/f/x/�/ �/�/�/�/�/�/?? ,?>?P?b?t?�?�?�? �?�?�?�?OO(O:O LO^OpO�O�O�O�O�O��O�O __$_6Y�$�FEAT_DEM�OIN  ;T��fP�<PNTINWDEX[[jQ�NP�ILECOMP �z����Q�iRIU�PSET�UP2 {�U��R�  N ��Q�S_AP2BC�K 1|�Y G �)7Xok%�_8o<P�P&oco9U�_ �oo�oBo�o�oxo �o1C�og�o�� ,�P����� ?��L�u����(��� Ϗ^�󏂏�)���M� ܏q������6�˟Z� ؟���%���I�[�� ������D�ٯh��� ���3�¯W��d��� ���@�տ�v�Ϛ� /�A�пe����ϛ�*� ��N���r���ߨ�=� ��a�s�ߗ�&߻��� \��߀��'��K��� o���|��4���X��� ���#���G�Y���}� �����B���f������1�Y�PP�_ }2�P*.VR8���*�������l PC���FR6:�2�V�TzPz��w�]PG���*#.Fo/��	��:,�^/�STM@i/�/ /�-M/�/�H�/?�'?�/8�/g?�GIFq?�?��%�?D?V?�?�JPG�?O�%O�?�?oOF�
JSyO�O��5C��OMO%
Java?Script�O�?�CS�O&_�&_�O �%Cascad�ing Styl�e Sheets�R_��
ARGNA�ME.DT�_��� \�_S_�A�T�_�_}�PDISP*�_���To�_�QLaZo�oCLLB.Z�Iwo2o$ :\�a\��o�i�AColl�abo�o�o
TP�EINS.XML��_:\![o�QC�ustom To�olbarbiPASSWORDQo~��FRS:\��dB`Passwo�rd Config���/��(�e� �������N��r�� ���=�̏a������ &���J���񟀟��� 9�K�ڟo�������4� ɯX��|���#���G� ֯@�}����0�ſ׿ f������1���U�� y��ϯ�>���b��� 	ߘ�-߼�Q�c��χ� ߽߫�L���p��� ��;���_���X��$� ��H�����~����7� I���m���� �2��� V���z���!��E�� i{
�.��d ����S�w p�<�`�/ �+/�O/a/��// �/8/J/�/n/?�/�/ 9?�/]?�/�?�?"?�? F?�?�?|?O�?5O�? �?kO�?�OO�O�OTO �OxO__�OC_�Og_ y__�_,_�_P_b_�_ �_o�_oQo�_uoo �o�o:o�o^o�o�o )�oM�o�o�� 6��l��%�7� �[����� ���D� ُh�z����3�,� i��������ßR���v������$FI�LE_DGBCK� 1|������ <� �)
SUMM?ARY.DG!�͜OMD:U���ِ�Diag Su�mmary����
CONSLOG���n���ٯ���Co�nsole lo�g���	TPACCN�t�%\������TP Acco�untin;����FR6:IPKD?MP.ZIPͿј�
�ϥ���Exc?eption"�ӻ���MEMCHEC�K��������-�M�emory Da�ta����6n =)��RIPE�~ϸ��%ߴ�%�� �Packet L<:���L�$�c���STAT��߭�� %A�St�atus��^�	F�TP����	���/�mment T�BD2�^� >I)�ETHERNE�w�
�d�u�﨡E�thernJ�1�figuraAϩ��?DCSVRF&����7����� ve�rify all�:����4��DIFF/��'���;�Q�diff��r�d�>��CHG01�������A����it�2���270���f�x3���I� �p�VT�RNDIAG.LASu&8����O Ope��L� ���nostic�����)VDEV�DAT�������Vis�De�vice�+IM�G��,/>/�/:��i$Imagu/+�UP ES/�/�FRS:\?Z=���Updates� ListZ?���� FLEXEVEAN��/�/�?���1 UIF EvM��M���-vZ)�CRSENSPK�/˞�\!O����CR_TAOR_P�EAKbOͩPSRBWLD.CM�O�͜E2�O\?.�PS�_ROBOWEL<S���:GIG��@_��?d_��GigE��(O��N�@�)}UQHADOW__�D_V_�_��Sha�dow Chansge����.dt�R?RCMERR�_�_��_oo��4`CFG� Erroro t�ailo MA��k�CMSGLIBgoNo`o�o|R�e���z0ic�o�a�)�`ZD0_O�osn��ZD�Pad��l �RNOTI��Rd���Notific����,�AG��P�ӟt� ��������Ώ]��� ��(���L�^�폂�� ����G�ܟk� ���� 6�şZ��~������ C�د�y����2�D� ӯh��������¿Q� �u�
�ϫ�@�Ͽd� v�Ϛ�)Ͼ���_��� ��ߧ�%�N���r�� �ߨ�7���[����� &��J�\��߀��� 3����i����"�4� ��X���|������A� ����w���0��= f�����O� s�>�bt �'�K��� /�:/L/�p/��/ �/5/�/Y/�/ ?�/$? �/H?�/U?~??�?1? �?�?g?�?�? O2O�? VO�?zO�OO�O?O�O cO�O
_�O._�OR_d_ �O�__�_�_M_�_q_ oo�_<o�_`o�_mo �o%o�oIo�o�oo �o8J�on�o�� 3�W�{�"�� F��j�|����/�ď�֏e������0��$�FILE_FRS�PRT  ��������?�MDONLY� 1|S�� �
 �)MD:�_VDAEXTP.ZZZ1�⏹�ț�6%NO �Back fil�e ���S�6P �����>��K�t��� ��'���ί]�򯁯� (���L�ۯp������ 5�ʿY�׿ Ϗ�$ϳ� H�Z��~�Ϣϴ�C� ��g���ߝ�2���V� ��cߌ�߰�?����� u�
��.�@���d�������C�VISBC�Kq�[���*.V�D����S�FR:�\��ION\DA�TA\��v�S��Vision VD���Y�k���� y��B�����x��� 1C��g���, �P����? �Pu�(�� ^��/��M/� q/�/>/�/6/�/Z/�/ ?�/%?�/I?[?�/?�?�?2?D?�?9�LU�I_CONFIG7 }S����;� $ �3v�{ S�;OMO_OqO�O�O�I#@|x�?�O�O�O_ _%\�OH_Z_l_~_�_ '_�_�_�_�_�_o�_ 2oDoVohozo�o#o�o �o�o�o�o
�o.@ Rdv���� ����*�<�N�`� r��������̏ޏ�� ���&�8�J�\�n��� �����ȟڟ쟃��� "�4�F�X�j������ ��į֯����0� B�T�f����������� ҿ�{���,�>�P� b����ϘϪϼ����� w���(�:�L�^��� �ߔߦ߸�����s� � �$�6�H���Y�~�� �����]������ � 2�D���h�z������� ��Y�����
.@ ��dv����U ��*<�` r����Q�� //&/8/�\/n/�/ �/�/;/�/�/�/�/? "?�/F?X?j?|?�?�? 7?�?�?�?�?OO�? BOTOfOxO�O�O3O�O �O�O�O__�O>_P_ b_t_�_�_/_�_�_�_ �_oo�_:oLo^opo��o�o$h  x��o�c�$FLUI�_DATA ~�����a�(a�dRESU_LT 3�ep� �T�/�wizard/g�uided/st�eps/Expert�o=Oas���������z��Continu�e with Gpance�:�L� ^�p���������ʏ܏,� � �b-�a�e>�0 �0`���c�a?��ps ���������ҟ��� ��,�>�P��0ow� ��������ѯ���� �+�=�O�a�?�1�C�zU�e�cllbs� ֿ�����0�B�T� f�xϊϜ�[������� ����,�>�P�b�t� �ߘߪ�i�{��ߟ�]�e�rip(pſ-� ?�Q�c�u����� ��������)�;�M� _�q����������������������`��e�#pTimeUS/DST	��� ����!3E~�Enabl(� y��������	//-/?/Q/�b��)�/M_q24 |�/�/??)?;?M? _?q?�?�?Tf�?�? �?OO%O7OIO[OmO O�O�Ob/t/�/�/Z��"qRegion �O5_G_Y_k_}_�_�_�_�_�_�_�America!�#o5o GoYoko}o�o�o�o�o�o�o��Ay�O�O3��O_qEditor�o����������+�=� � T�ouch Pan�el rs (re�commenp�) K�������Ə؏��� � �2�D�|�%���I[qaccesoܟ� ��$�6��H�Z�l�~�����C�onnect t�o Network��֯�����0��B�T�f�x�����x�B�@��}����,!���s Introduct!_4�F�X�j�|� �Ϡϲ��������� �0�B�T�f�xߊߜ�`����������  ɿ��"�i�{�� ������������� /�A� �e�w������� ��������+="�H�3��+� O�����  2DVhz�K�� ����
//./@/ R/d/v/�/�/Yk} �/�??*?<?N?`? r?�?�?�?�?�?�?� �?O&O8OJO\OnO�O �O�O�O�O�O�O�/_ �/1_�/X_j_|_�_�_ �_�_�_�_�_oo0o BoS_foxo�o�o�o�o �o�o�o,>�O _!_�E_���� ���(�:�L�^�p� ����So��ʏ܏� � �$�6�H�Z�l�~��� O��s՟���� � 2�D�V�h�z������� ¯ԯ毥�
��.�@� R�d�v���������п ⿡��ş'�9���`� rτϖϨϺ������� ��&�8���\�n߀� �ߤ߶���������� "�4��=��a��M� ������������0� B�T�f�x���I߮��� ������,>P bt�E��i�� ��(:L^p �������� / /$/6/H/Z/l/~/�/ �/�/�/�/���� /?�V?h?z?�?�?�? �?�?�?�?
OO.O� ROdOvO�O�O�O�O�O �O�O__*_<_�/? ?�_C?�_�_�_�_�_ oo&o8oJo\ono�o ?O�o�o�o�o�o�o "4FXj|�M_ __q_��_���0� B�T�f�x��������� ҏ�o���,�>�P� b�t���������Ο�� ���%��L�^�p� ��������ʯܯ� � �$�6�G�Z�l�~��� ����ƿؿ���� � 2��S��w�9��ϰ� ��������
��.�@� R�d�v߈�G��߾��� ������*�<�N�`� r��Cϥ�g���ύ� ��&�8�J�\�n��� �������������� "4FXj|�� ��������- ��Tfx���� ���//,/��P/ b/t/�/�/�/�/�/�/ �/??(?�1U? ?A�?�?�?�?�? O O$O6OHOZOlO~O=/ �O�O�O�O�O�O_ _ 2_D_V_h_z_9?�?]? �_�_�?�_
oo.o@o Rodovo�o�o�o�o�o �O�o*<N` r������_�_ �_�_#��_J�\�n��� ������ȏڏ���� "��oF�X�j�|����� ��ğ֟�����0� ���u�7������� ү�����,�>�P� b�t�3�������ο� ���(�:�L�^�p� ��A�S�e��ω��� � �$�6�H�Z�l�~ߐ� �ߴ��߅������ � 2�D�V�h�z���� �����������@� R�d�v����������� ����*;�N` r������� &��G	�k-� �������/ "/4/F/X/j/|/;�/ �/�/�/�/�/??0? B?T?f?x?7�?[�? �?�?OO,O>OPO bOtO�O�O�O�O�O�/ �O__(_:_L_^_p_ �_�_�_�_�_�?�_�? o!o�OHoZolo~o�o �o�o�o�o�o�o  �ODVhz��� ����
���_%o �_I�s�5o������Џ ����*�<�N�`� r�1������̟ޟ� ��&�8�J�\�n�-� w�Q���ů������ "�4�F�X�j�|����� ��Ŀ�������0� B�T�f�xϊϜϮ��� ��������ٯ>�P� b�t߆ߘߪ߼����� ����տ:�L�^�p� ����������� � �$������i�+ߐ� ������������  2DVh'��� ����
.@ Rdv5�G�Y��}� ��//*/</N/`/ r/�/�/�/�/y�/�/ ??&?8?J?\?n?�? �?�?�?�?��?�O �4OFOXOjO|O�O�O �O�O�O�O�O__/O B_T_f_x_�_�_�_�_ �_�_�_oo�?;o�? _o!O�o�o�o�o�o�o �o(:L^p /_������ � �$�6�H�Z�l�+o�� Oo��sou����� � 2�D�V�h�z������� ����
��.�@� R�d�v���������}� ߯����ٟ<�N�`� r���������̿޿� ��ӟ8�J�\�nπ� �Ϥ϶���������� ϯ��=�g�)��ߠ� ������������0� B�T�f�%ϊ����� ��������,�>�P� b�!�k�Eߏ���{��� ��(:L^p ����w���  $6HZl~� ��s�������/�� 2/D/V/h/z/�/�/�/ �/�/�/�/
?�.?@? R?d?v?�?�?�?�?�? �?�?OO���]O /�O�O�O�O�O�O�O __&_8_J_\_?�_ �_�_�_�_�_�_�_o "o4oFoXojo)O;OMO �oqO�o�o�o0 BTfx���m_ �����,�>�P� b�t���������{oݏ �o��o(�:�L�^�p� ��������ʟܟ� � �#�6�H�Z�l�~��� ����Ưد����͏ /��S��z������� ¿Կ���
��.�@� R�d�#��ϚϬϾ��� ������*�<�N�`� ���C���g�i����� ��&�8�J�\�n�� ����u�������� "�4�F�X�j�|����� ��q�������	��0 BTfx���� �����,>P bt������ �/����1/[/ �/�/�/�/�/�/�/ ? ?$?6?H?Z?~?�? �?�?�?�?�?�?O O 2ODOVO/_/9/�O�O o/�O�O�O
__._@_ R_d_v_�_�_�_k?�_ �_�_oo*o<oNo`o ro�o�o�ogOyO�O�O �o�O&8J\n� ��������_ "�4�F�X�j�|����� ��ď֏�����o�o �oQ�x��������� ҟ�����,�>�P� �t���������ί� ���(�:�L�^�� /�A���e�ʿܿ� � �$�6�H�Z�l�~ϐ� ��a���������� � 2�D�V�h�zߌߞ߰� o��ߓ��߷��.�@� R�d�v������� ������*�<�N�`� r��������������� ��#��G	�n� ������� "4FX�|�� �����//0/ B/T/u/7�/[]/ �/�/�/??,?>?P? b?t?�?�?�?i�?�? �?OO(O:OLO^OpO �O�O�Oe/�O�/�O�O �?$_6_H_Z_l_~_�_ �_�_�_�_�_�_�? o 2oDoVohozo�o�o�o �o�o�o�o�O_�O% O_v����� ����*�<�N�o r���������̏ޏ�� ��&�8�J�	S- w���cȟڟ���� "�4�F�X�j�|����� _�į֯�����0� B�T�f�x�����[�m� ���󿵟�,�>�P� b�tφϘϪϼ����� �ϱ��(�:�L�^�p� �ߔߦ߸������� � ��ѿ�E��l�~�� ������������ � 2�D��h�z������� ��������
.@ R�#�5�Y�� ��*<N` r��U����� //&/8/J/\/n/�/ �/�/c�/��/�? "?4?F?X?j?|?�?�? �?�?�?�?�??O0O BOTOfOxO�O�O�O�O �O�O�O�/_�/;_�/ b_t_�_�_�_�_�_�_ �_oo(o:oLoOpo �o�o�o�o�o�o�o  $6H_i+_� O_Q����� � 2�D�V�h�z�����]o ԏ���
��.�@� R�d�v�����Y��} ߟ񟵏�*�<�N�`� r���������̯ޯ� ���&�8�J�\�n��� ������ȿڿ쿫��� ϟ�C��j�|ώϠ� ������������0� B��f�xߊߜ߮��� ��������,�>��� G�!�k��Wϼ����� ����(�:�L�^�p� ����S߸�������  $6HZl~� O�a�s�����  2DVhz��� �����
//./@/ R/d/v/�/�/�/�/�/ �/�/���9?�`? r?�?�?�?�?�?�?�? OO&O8O�\OnO�O �O�O�O�O�O�O�O_ "_4_F_??)?�_M? �_�_�_�_�_oo0o BoTofoxo�oIO�o�o �o�o�o,>P bt��W_�{_� �_��(�:�L�^�p� ��������ʏ܏�� �$�6�H�Z�l�~��� ����Ɵ؟꟩�� /��V�h�z������� ¯ԯ���
��.�@� ��d�v���������п �����*�<���]� ���C�EϺ������� ��&�8�J�\�n߀� ��Q������������ "�4�F�X�j�|��M� ��q��������0� B�T�f�x��������� ������,>P bt������ ������7��^p ������� / /$/6/��Z/l/~/�/ �/�/�/�/�/�/? ? 2?�;_?�?K�? �?�?�?�?
OO.O@O ROdOvO�OG/�O�O�O �O�O__*_<_N_`_ r_�_C?U?g?y?�_�? oo&o8oJo\ono�o �o�o�o�o�o�O�o "4FXj|�� �����_�_�_-� �_T�f�x��������� ҏ�����,��oP� b�t���������Ο�� ���(�:���� �A�����ʯܯ� � �$�6�H�Z�l�~�=� ����ƿؿ���� � 2�D�V�h�zό�K��� o��ϓ���
��.�@� R�d�v߈ߚ߬߾��� ������*�<�N�`� r���������� ����#���J�\�n��� �������������� "4��Xj|�� �����0 ��Q�u7�9�� ���//,/>/P/ b/t/�/E�/�/�/�/ �/??(?:?L?^?p? �?A�?e�?�?�/ O O$O6OHOZOlO~O�O �O�O�O�O�/�O_ _ 2_D_V_h_z_�_�_�_ �_�_�?�?�?o+o�? Rodovo�o�o�o�o�o �o�o*�ON` r������� ��&��_/o	oS�}� ?o����ȏڏ���� "�4�F�X�j�|�;�� ��ğ֟�����0� B�T�f�x�7�I�[�m� ϯ������,�>�P� b�t���������ο�� ���(�:�L�^�p� �ϔϦϸ����ϛ��� ��!��H�Z�l�~ߐ� �ߴ���������� � ߿D�V�h�z���� ��������
��.��� ���s�5ߚ������� ����*<N` r1������ &8J\n� ?��c������/ "/4/F/X/j/|/�/�/ �/�/�/��/??0? B?T?f?x?�?�?�?�? �?��?�O�>OPO bOtO�O�O�O�O�O�O �O__(_�/L_^_p_ �_�_�_�_�_�_�_ o o$o�?EoOio+O-o �o�o�o�o�o�o  2DVhz9_�� ����
��.�@� R�d�v�5o��Yo��͏ ����*�<�N�`� r���������̟�� ��&�8�J�\�n��� ������ȯ��я���� ��F�X�j�|����� ��Ŀֿ�����ݟ B�T�f�xϊϜϮ��� ��������ٯ#��� G�q�3��ߪ߼����� ����(�:�L�^�p� /ϔ��������� � �$�6�H�Z�l�+�=� O�a���������  2DVhz��� �����
.@ Rdv����� ������/��</N/`/ r/�/�/�/�/�/�/�/ ??�8?J?\?n?�? �?�?�?�?�?�?�?O "O��/gO)/�O�O �O�O�O�O�O__0_ B_T_f_%?w_�_�_�_ �_�_�_oo,o>oPo boto3O�oWO�o{O�o �o(:L^p ������o� � �$�6�H�Z�l�~��� ����Ə�o珩o��o 2�D�V�h�z������� ԟ���
���@� R�d�v���������Я �����׏9���]� �!�������̿޿� ��&�8�J�\�n�-� �Ϥ϶���������� "�4�F�X�j�)���M� ���߅�������0� B�T�f�x������ �������,�>�P� b�t���������{��� ������:L^p �������  ��6HZl~� ������/�� ��;/e/'�/�/�/ �/�/�/�/
??.?@? R?d?#�?�?�?�?�? �?�?OO*O<ONO`O /1/C/U/�Oy/�O�O __&_8_J_\_n_�_ �_�_�_u?�_�_�_o "o4oFoXojo|o�o�o �o�o�O�O�O	�O0 BTfx���� �����_,�>�P� b�t���������Ώ�� ����o�o�o[� ��������ʟܟ� � �$�6�H�Z��k��� ����Ưد���� � 2�D�V�h�'���K��� o�Կ���
��.�@� R�d�vψϚϬϾ�Ͽ ������*�<�N�`� r߄ߖߨߺ�y��ߝ� ����&�8�J�\�n�� ������������� ��4�F�X�j�|����� ������������- ��Q����� ���,>P b!������� �//(/:/L/^/ /A�/�/y�/�/ ? ?$?6?H?Z?l?~?�? �?�?s�?�?�?O O 2ODOVOhOzO�O�O�O o/�/�/�O_�/._@_ R_d_v_�_�_�_�_�_ �_�_o�?*o<oNo`o ro�o�o�o�o�o�o�o �O_�O/Y_� �������� "�4�F�X�o|����� ��ď֏�����0� B�T�%7I��m ҟ�����,�>�P� b�t�������i�ί� ���(�:�L�^�p� ��������w������� ��$�6�H�Z�l�~ϐ� �ϴ��������ϻ� � 2�D�V�h�zߌߞ߰� ��������
�ɿۿ� O��v������� ������*�<�N�� _��������������� &8J\�} ?�c����� "4FXj|�� �����//0/ B/T/f/x/�/�/�/m �/��/�?,?>?P? b?t?�?�?�?�?�?�? �?O�(O:OLO^OpO �O�O�O�O�O�O�O _ �/!_�/E_?	_~_�_ �_�_�_�_�_�_o o 2oDoVoOzo�o�o�o �o�o�o�o
.@ R_s5_��mo� ����*�<�N�`� r�������gȍޏ�� ��&�8�J�\�n��� ����c��џ��� "�4�F�X�j�|����� ��į֯������0� B�T�f�x��������� ҿ�������ٟ#�M� �tφϘϪϼ����� ����(�:�L��p� �ߔߦ߸������� � �$�6�H���+�=� ��a���������� � 2�D�V�h�z�����]� ��������
.@ Rdv���k�}�������$FMR�2_GRP 1���� ��C4  B�.��	 ��9K^6F@ a@��6G�  �Fg?�fC�8R�y�?�  ��66��X���875�t��5���5�`+�yA�  �/+BH�w-%@'S339%�5[/l-6@6!�/xl/�/ �/�/�/?�/&??J?�5?G?�?k?�?��_�CFG �T�K�?�? OO�9NO� 
F0�FA K@�<RM_C�HKTYP  ���$&� RO=Ma@_MINg@��W���@�R X�SSB�3�� 7�O���C�O�O�5TP_D�EF_OW  ��$WIRCO�Mf@_�$GENOVRD_DO�F���E]TH��D �dbUdKT_ENB�7_ KPRAVC���G�@ �@Y�O�_�?oyo�&oI* �QOU*�NAIRI<�@��oGo��o�o�o��C�p3@��O:��B��+sL�i�O�PSM�T��Y(�@
t��$HOSTC�219��@�5� MC��R{����  27.�00�1�  e �]�o�������K�ď�֏��������	a�nonymous@!�O�a�s����� �4��������D� !�3�E�W�i������� ��ï柀�.���/� A�S���课�П��� �Ŀ����+�r�O� a�sυϗϺ����� ����'�n������� �ϓ�ڿ���������� F�#�5�G�Y�k���� �����������B�T� f�C�z�g��ߋ����� �������	-P� ����u����� �(�:�<)p�M_ q�������� /$ZlI/[/m// �/����//�/D !?3?E?W?/?�?�? �?�?�/�?./OO/O AOSO�/�/�/�/�?�O ?�O�O__+_r?O_ a_s_�_�_�O�?O�_��_oo'o�t�qEN�T 1�hk P�!�_no  �p \o�o�o�o�o�o�o �o�o:_"�F �j�����%� �I��m�0���T�f� Ǐ��돮��ҏ3��� ,�i�X���P���t�՟ ��៼�
�/��S�� w�:���^���������ฯ�ܯ=� �QU�ICC0J�&�!�192.168.O1.10c�X�1��v�8��\�2�ƿؿ�9�!ROUTER:��!��a��?PCJOG��e�_!* ��0��~U�CAMPRT��ƶ�!�����RT�S���x� !S�oftware �Operator? PanelU߇����7kNAME �!Kj!ROBO�����S_CFG �1�Ki ��Auto-s�tarted�DFTP�Oa�O�_ ���O����������E_ �.�@�R�u�c�	��� ��������cN:�L�^� ;r���R���� ����%H� [m���jO|O �O�O4!/hE/W/i/ {/�/T�/�/�/�/�/ /�//?A?S?e?w?�? ����??�?</O +O=OOO?sO�O�O�O �O�?`O�O__'_9_ K_�?�?�?�?�O�_�? �_�_�_o#o�OGoYo ko}o�o�_4o�o�o�o �of_x_�_g�o ��_�����o� �-�?�Q�tu���� ����Ϗ�(:L^ `�2��q��������� ��ݟ���%�H�ʟ [�m�����������  �ί4�!�h�E�W�i� {���T���ÿտ�
� Ϟ�/�A�S�e�w�����_ERR ���ڇϗ�PDUSI�Z  �^6�����>��WRD �?(����  �guest ���+�=�O�a����SCD_GROUoP 3�(� ,��"�IFT��$P�A��OMP��� ��_SH��ED��� $C��COM���TTP_AUT�H 1��� <�!iPenda�nm�x�#�+!K?AREL:*x����KC�������VISION SET��(����?�-�W�R���v������������������G�C�TRL ����a�
��F�FF9E3���FRS:DEFA�ULT�FA�NUC Web ?Server�
t dG����/� �2DV��WR_C�ONFIG �.��������IDL_CPU_kPC� �B����� BH�MIN�����GNR_I�O������ȰHM�I_EDIT =���
 ($/C/ ��2/k/V/�/z/�/�/ �/�/�/?�/1??U? @?y?d?�?�?./�?�? �?�?OO?OQO<OuO `O�O�O�O�O�O�O�O�__;_�NPT_�SIM_DO��*NSTAL_S7CRN� �\UQ�TPMODNTOqL�Wl[�RTYbXp�qV�K�ENB�W��ӭOLNK 1�����o%o7o�Io[omoo�RMAS�TE��Y%OSLAVE �����eRAMCACH�E�o�ROM�O_CcFG�o�S�cUO'���bCMT_OPp�  "��5sYCL�o�u� _ASG 19����
 �o� ������"�4��F�X�j�|����kwrN�UM����
�bI�P�o�gRTRY_�CN@uQ_UP)D��a��� �bp�b��n��M��а�P}T?��k ��._������ɟ۟� �S���)�;�M�_�q�  �������˯ݯ�~� �%�7�I�[�m���� ����ǿٿ�����!� 3�E�W�i�{�
ϟϱ� �������ψϚ�/�A� S�e�w߉�߭߿��� ������+�=�O�a� s���&�������� ����9�K�]�o��� ��"����������� ����GYk}�� 0����� CUgy��,> ���	//-/�Q/ c/u/�/�/�/:/�/�/ �/??)?�/�/_?q? �?�?�?�?H?�?�?O O%O7O�?[OmOO�O �O�ODOVO�O�O_!_ 3_E_�Oi_{_�_�_�_ �_R_�_�_oo/oAo �_�_wo�o�o�o�o�o `o�o+=O�o s�����\n ��'�9�K�]�����������ɏۏi�c�_�MEMBERS �2�:� �  $:� ����v���1���R�CA_ACC 2��� �  [��bw�f�l�6"���W  l�l���6 М������J�����a�BUF00�1 2�n�= ��u0  u0���,�:�I��V�e�r��������������������R���������U)��7��F��S���b��pul�u ������Ҥ�ҤӴҤy��������U��(�5�UD�Q�a�n�}|�� H Q�-����J�*J�����GJ�TJ�dJ�q�J�A���J��J���J��J��J��J��JJ����ߙ2� ���������x!��)�t@ �0� �9��A��I��Q� �Y��a��i��q� �y������� ���¡��©��±� �¹�������ɠʡС �ء�������� ���������� ��!��)��1�� 9��A��I��P�R� X�U�a�U�i�UҲ�x� Uҁ�U҉�Uґ�U�J� ��Uҩ�Uұ�Uҹ�U� ��U�ɰU�ѰU�ٰ���ߙ3������ ���!�/��1�?� �A�O��Q�_��a� o��q��⁢�Ö� ���Ö⡢�ÖⱢ�� ������l�У����� ��������l��� ��'��)�7��9� G��I�W�^��`�o� ^��x���^򉲗�^� S䠳��^򱲿�^������^�Ѳ������C�FG 2�n� Q4��l�l�<l��47��HIS�钜n� ��� 2025-12�-�l� 6�4�����h �  7 p + �xl�;s�1O4 �l�7 ��o9 ���b��(7[~�qq1�-3�  � # &f � ' "7�� + P
X
`
� �  ��   $ } �  8 @�	��{�9, ��~��!  8�$�d�q4[}�RM29}	�R/d/v/��/�/�/�/�-( �%  ��-��R  *gl��,B��=/*?<?N?`? r?�?�?�?�?�??? OO&O8OJO\OnO�O �O�O�?�?�O�O�O_ "_4_F_X_j_|_�O�O �_�_�_�_�_oo0o BoTo�O��[m
7d_o�o�o�o�+ _� %g>� "�"	�b  3"!"�o;TM_8 cm8� �����c��b�|�b� +  X� U � X|c	,: �J"0  }Q�1 
 R T"��: b(:�q %/7/m��������ǏPُ��(5�c��2!R ,�� 1� \�_ �_I�[�m�������� ǟٟ럑_4�!�3�E� W�i�{�������ï�� �Я��/�A�S�e� w�����ү������ ��+�=�O�a�s�ao N�Ѐo�o
3���ϐ�����:q� Bq� Dqe�	e�I^� J��e�r�H`r�v
qm�� ���ߧ�ҵ�ҽ�҈� ��� ?�G(O� 2_�q���"J� .q Z�  ��J�\�������@��������*T�[� 6�� �澿пr����� ����������K� ]�J\n���� ���#5"4F Xj|����� �//0/B/T/f/�x/�/�/��_I_C�FG 2��� �H
Cycle� Time�B�usy�Idl��"�min�+�1Up�&��Read�'DCow8?F� 1�#�Count�	N'um �"����<�p>�qaPROG��"�������)/softpa�rt/genli�nk?curre�nt=menup�age,1133,�gOO&O8O<b5�leSDT_ISO_LC  ����p��/J23_DS/P_EN>�vK0~�@INC ��M|s�@A   ?&p�=���<#�
<�A�I:�o&��N`_t�O<_�GOB�0�C�C"�1�FVQG_�GROUP 1�vvK1r<�P�Cy�_D_?x�?�_pQ�_o.o@o�_ dovo�o�ow,_NY�G_IN_AUT�O �MPOSRE�^_pVKANJI_�MASK v�HqR�ELMON ��˔?��y_ox������.6r�3��7ĲC���u�o�DKCwL_L�`NUM(���EYLOGGING ����Q�E�0�LANGUAGE� ��~���DEFAULT� ����LG�!���:2�?�3��80VЬ��'�� _ � 
��ћ���GOUF ;��
~��(UT1:%�� � �-�?�Q�h� u���������ϟ����(g4�8i�N_DISP ��O�8�_�_��LOCT3OL����Dz<�A��A��GBOOK ���d�1
�
�۠������#�5��G�Y�i���3{�W�	��쉞QQJ¿Կ1���_BUFF ;2�vK ��Ё25
�ڢVB&�7� Collaborativ�=�O� �ώϠϲ��������� '��0�]�T�fߓߊ�����DCS � �9�B�Ax���Rh�%��-�?�Q���IO 2��� ���Q��������� ����*�<�N�b�r� ���������������&:e�ER_ITMsNd�o��� ����#5G Yk}�����p����hSEV�`��MdTYPsN��c/u/�/
-�aRS�T5���SCRN__FL 2�s��0����/??1?C?U?�g?�/TPK�sOR">��NGNAM�D���~�N�UPS_AC�R� �4DIGI��8+)U_LOA�D[PG %�:%�T_NOVIC�Et?��MAXUA�LRM2��a���2�E
ZB�1_P�5�`� ��y�Z@CY���˭�O+���ۡ�D|PPw 2�˫ �Uf	R/_
_C_._g_y_ \_�_�_�_�_�_�_�_ oo?oQo4ouo`o�o |o�o�o�o�o�o) M8qTf�� �����%��I� ,�>��j�����Ǐُ �����!���W�B� {�f�������՟���� ܟ�/��S�>�w��� l�����ѯ��Ư�� +��O�a�D���p����RHDBGDEF ���E�ѱO��_L?DXDISA�0�;�c�MEMO_AP޻0E ?�;
 ױ��3�E�W�i��{ύϟϱ�Z@FRQ_CFG ��Gm۳A ��@�����<��d%�� ���t���B��K���*i�/k� **:tҔ�g�y�� ���߱��������� �J�Es�J d������,(H���[� ����@�'�Q�v�]� ���������������*NPJISC 31��9Z� ���� ��ܿ�����	Z�l_MSTR ��#-,SCD 1�"͠{��� �����//A/ ,/e/P/�/t/�/�/�/ �/�/?�/+??O?:? L?�?p?�?�?�?�?�? �?O'OOKO6OoOZO �O~O�O�O�O�O�O_ �O5_ _Y_D_i_�_z_ �_�_�_�_�_�_o
o oUo@oyodo�o�o�o �o�o�o�o?*�cN�MK���;љ$MLT�ARM���N��r ��հ��>İMETPU��zr���CNDSP?_ADCOL%�ٰ�0�CMNTF� �9�FNb�f�7�FS�TLI��x�4 �;ڎ�s����9�_POSCF��q��PRPMe��STvD�1�; 4�#�
v��qv����� r��������̟ޟ � ��V�8�J���n����¯�������9�SI�NG_CHK  }��$MODA����t�{�~2�DE�V 	�	M�C:f�HSIZE���zp�2�TASK� %�%$12�3456789 �ӿ�0�TRIG ;1�; lĵ��2ϻ�!�bϻ�YP蠱��H�1�EM_�INF 1�N��`)AT&F�V0E0g���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ��2�ԁH6�^���Rφ��A��߶�q��������  ��5������ߏ�B� ������������1� C�*�g��,��P�b� t������R�?�� �u0������ ���������M q ���Z���/ �%/��[/ 2 �/�/h�//�/�/� 3?�/W?>?{?�?@/�? d/v/�/�/O�//OAO x?eO?�ODO�O�O�O|�O_�NITORÀ�G ?z�   	EXEC1~s�&R2,X3,X4,X5�,X��.V7,X8,X9~s'R�2�T+R�T7R �TCR�TOR�T[R�TgR��TsR�TR�T�R�S2��X2�X2�X2�X2��X2�X2�X2�X2��X2h3�X3�X3�7R2�R_GRP_�SV 1��� a(��o.���_D�B����cION_DB�<��@�zq  ��$��$��Y�1t �&zp'>w�Zp��Zp�Y��@N Kp"ZKp#>{��p�Y�-ud1������8�PG_JOG� �ʏ�{
�2��`:�o�=���?����@0�B��~\�n���������H�?��C�@�pŏ׏���  ������qL_NAM�E !ĵ8���!Defaul�t Person�ality (from FD)qp�0�RMK_ENOgNLY�_�R2�a� 1�L�XL��8�gpl d����şן���� �1�C�U�g�y����� ����ӯ���	���� 
�<�N�`�r�������p��̿޿� :� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w���������������+��<�Se w�������x��A�a��AB�Bw��Pf ������/!/ 3/E/W/i/{/�/�/�/ ���/�/??/?A? S?e?w?�?�?�?�?�? �?�?�/�/+O=OOOaO sO�O�O�O�O�O�O�O __'_9_&O�S^Q��x_�]�rd�d �_�^�_�_�W��_[�op.ooRog Fh qogoyo�o�o�o�o�o�E`�p"|��Fe	�`[oUgy8qK�A�\����s� A� ��y@h�Q�Q��"����Tk\$�_�  ��P�P�E�xC�  � I�@oa�<o��p��������ߏ
f�Q*������0��PCr� �� 3r �.� @oD�  A�?�G��-�?.I�.@I��A����  ;��	lY�	 ��X  ������� �, � �����̀�K�o�����]�K��K]�/K	�.��w�r_x	��̀@
�)��b�1�����I��Y�����T;f�Y�{S���3�	���I�>J���;Î?v�>��=@�O����E�΂ѯ�עZ���wp��u�� kD!�3��7p�g  �  ��9�͏W���	'�� � u�I� �  ��u���:�È��È�=��ͱ�E�@��ǰ�3��\�3��E�&���N�pC�  'Y�&�Z�i�b�1@f�i�n�C���¢I�C����b	��r�� p����B�p�Ŕq���}ر�.DzƏ<ߛ�`�K߸pߖ߁��������А #4P����.z��d�  �Pؠ?��ff�_��	�� !2p>�P��8.f�t�>L���U���(.��P��������
����� x��;e��m��KZ;�=�g;�4�<<a����%�G��3�|���p?fff?ذ�?&S���@=0e�?��q�+�r N�Z���I���G���7� ��(�����!E0 iT����+��F�p���#�� D��w��� ����//=/(/ a/L/�/p/��/�p� 6�/Z#?�/ ?Y?k? }?��?�?>?�?�?�? �?�?1O�����KD�y�^KCO�OO�O��ɃذO�O�O�Oai����J��}�DD1���.�D��@�AmQa���9N,ȴA;��^@��T@|j�@$�?�V��>�z�ý���=#�
>\�)?��
=�G}�-]�{=����,��C+�ןBp���P��6���C98R����?N@��(���5-]G�p��Gsb�F�}��G�>.E�V�D�Kn����I�� F�W��E��'E����D��;n����I��`E����G��cE�vmD���-_�oQ_ �o�o�o �o$H 3X~i���� �����D�/�h� S���w��������я 
���.��R�=�v�a� s�����П����ߟ� �(�N�9�r�]����� ����ޯɯۯ���8� #�\�G���k������� ڿſ���"��F�1� C�|�gϠϋ��ϯ����������P(�Q343�] �����Q�	�x9�Oߵ53~�mm��aҀ5Q�߫�a�Ǔ����ߵ1��������1��U�C�(y�g��%P�P���!�/��'���
���.������4�;�t� _��������������� :%��/�/d������� �7%[I�m���027� � B�S@J@�CH#PzS@�0@ZO/1/@C/U/g/y/�-�#���/�/�/�/�/�3?��3�� @�35�0�0�!3��5
 ?f?x?�?�? �?�?�?�?�?OO,Op>OPO�Z@1 �������c/�$MR�_CABLE 2�ƕ� ��TT��&�ڰO���O �)�@���C_���_ O_u_7_I__�_�_�_ �_�_o�_�_oKoqo 3oEo{o�o�o�o�o�o �o�o�oGm/�K!�"���O�����ذ�$�6����*Y�** �COM� ȖI����~D�f�#%�% 234567O8901���� ��HÏ��� � !� ��!
���M�not sent� b��W���TESTFECS�ALGR  egD�*!d[�41�
k�������$pB����������� 9U�D1:\main�tenances�.xmlğ�  �C:�DEF�AULT�,�BGR�P 2�z�  嬓 ;��%  ��%!1st cl�eaning o�f cont. �v�ilatio�n 56��ڧ�!0�����+B��*�`����+��"%���mech��cal� check1�  �k�0u�|��ԯ����Ϳ߿��@���rollerS�e�w�ū��m���ϣϵ�@�Bas�ic quarterly�*�<�ƪ,\�)�;�M�_�q�8�cMJ��ߓ "8��!� ���ߕ ��� ��+�=��C�g��ߋ�ʦ�߹���������@�Overghau�ߔ��?�C x� I�P����@}���������� $n� ������)l�ASe w������ � +=O�s� ������/R �9/�(/��/�/�/ �/�//�/�/N/#?r/ G?Y?k?}?�?�/�?? ?�?8?OO1OCOUO �?yO�?�?�O�?�O�O �O	__jO?_�O�Ou_ �O�_�_�_�_�_0_o T_f_;o�__oqo�o�o �o�_�oo,oPo% 7I[m�o��o�o ����!�3�� W��������ÏՏ �6����l����e� w���������џ�2� �V�+�=�O�a�s� �����ͯ���� '�9���]�������� ��ɿۿ���N�#�r� ��YϨ�}Ϗϡϳ��� ���8�J��n�C�U� g�yߋ��ϯ������ 4�	��-�?�Q��u� �����ߞ�������� �f�;�������� ���������P��� t�I[m���� ��:!3E W�{��� � ��//lA/�� w/��/�/�/�/�/X*�"	 X�/?.?@?�)B a/o?m/o%w? �?�?}?�?�?OO�? �?OOaOsO1OCO�O�O �O�O�O__'_�O�O ]_o_�_?_Q_�_�_�_��_�_�\ Џ!?�  @�!  M?HoZolo�&4o�o�oܽo�(*�o** F�@ �Q�V�` o'9�o]o�����/^&�o� ����/�A�S�e� ��#�����я��� ��+�q�����7��� ����k�͟ߟ��I� [���K�]�o���C������ɯ��o$�!��$MR_HIST� 2��U#�� �
 \7"$ 23�45678901P3�;���b2�90/ ����[���./���� ǿٿF�X�j�!�3ρ� ����{��ϟ����� B���f�x�/ߜ�S��� �߉��߭��,���P��t��=��$�S�KCFMAP  ]�U&��b�
�� ����ON?REL  �$#�������EXCFE�NB�
����&�F�NC-��JOGO/VLIM�d#�v���KEY�y���_PAN������RUNi�y����SFSPDTY�PM����SIGN|��T1MOTk�����_CE_G�RP 1��U ��+�0�ow�#d� �����& �6\�7y� m���/�4/F/ -/j/!/t/�/�/�/{/��/�/�/?�+��QZ_EDIT
�����TCOM_CFG 1���0�}?�?��? 
^1SI 	�N����?�?��!�?$O����?XO~78T_ARC_*��X�T_MN_oMODE
�U:�_SPL{O;�UA�P_CPL�O<�N�OCHECK ?��� ��  _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo���NO_WAITc_L	S7> NTf1�����%��qa_7ERRH2��������?o�o�o�o��POGj�@O�cӦm�|�g?n��<���?���t��|a~�bPARAM�b]����t^��8
�.�@� =  n�]�o�w�Q������� ����Ϗ�)��7��[�m� �����ODRDSP�C8��OFFSET_C�ARI0�OǖDIS�ԟœS_A�@AR�K
T9OPEN_FILE��1T6��0OPTION_�IO����K�M_P�RG %��%$�*����'�WO�-�Ns�ǥ� ��5�9���	 �������>d���RG�_DSBL  �����jN���RI_ENTTO���C�����A ��U^�@IM_DS����r��V��LCT �{mP2ڢ�3̹���d��%���_PEqX�@���RAT�G� d8��̐UP� װ�:����`S�e�Kωϗ��$�r�2G�L�XLwȚ�l� ��������'�9�K� ]�o߁ߓߥ߷����߀�����#�5�G���2 ��v�������������e�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?�q1�~?�?�?�?�? �?�?�?O O2ODO�yA�a�tn?~M��~O�O�P�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�O�Oo $o6oHoZolo~o�o�o �o�o�o�o�o �_ oVhz���� ���
��.�@�R�0d�QOES������
B�d�ӏ�ʏ� �������Y�D�}�0��r���������ԟ ڟ���p���=�M��q�	`��������c�:�o�¯ԯ�����A�  P�k�C�C�ڰ"ڰ����O��/  ���-���~)�C�  �t� k���g�����Կ��ѿ�
�5���_:�ĳ�OU����/��/��H��n�� o� ^�\�� @D�  p�?��v�\�?:px�:qC�4r�p�(��  ;��	l��	 ��X  ������� �,? � ��������Hʪ�����H���Hw�_zH�����8�B���B�  �Xѐ�`�o�*��3�	���t�>u���fC{�����:pB\�
��Ѵ9:qK�t�� ����$����*��� DP��^��b�g  �  �h������)�	'� � ���I� � � ��'�=��q�����t�@��@��!�b��^;b�t��U�(�N��r�  '���E�C�И�t�C��И��ߗ���jA�@!�����%�B�� ���,���H:qDz �k�ߏz���w�����А 4P��D�:uz:���	f�~�?�ff'�&8� ]�mb�8:p��>L��H���$�(:p�P���	������:� �x�;e�m"��KZ;�=g;�?4�<<���E/�Tv��b���?offf?�?&� �)�@=0�%?��%_9��}!��$� x��/v��/f'��W,? ?P?;?t?_?�?�?�? �?�?�?O�?(OOLO �/�/�/EO�OAO�O�O �O�O_�O_H_3_l_ W_�_{_�_�_1��_A� ��eO+o�ORooOo�o �o�oK/�o�omo�o@*'`+�,�zt���CL�H��}?�����
������u����#D1�/n�t��p�qޜ�@I�h~,���A;�^@���T@|j@$��?�V�n�z��ý��=#��
>\)?���
=�G�����{=��,���C+��Bp�����6��C98R���?}p���(��5���G�p�Gsb��F�}�G�>�.E�VD�K�L����I��� F�W�E���'E���D���;L����I���`E�G���cE�vmD���\�՟��ҟ���/� �S�>�w�b������� ѯ�������=�(� :�s�^���������߿ ʿ�� �9�$�]�H� ��lϥϐϢ������� ��#��G�2�W�}�h� �ߌ��߰�������� 
�C�.�g�R��v�� �������	���-�� Q�<�u�`�r������� ������'M�=(�34�]O!����8h~�%3�~�m����5qQ������<�!���  �`N�r��	eP@"P��Q�_/V�/9/$/]/H)����c/j/�/�/�/�/�/ �/�/!??E?0?i?T?�"&�_�_�?�?�8� �?�?O�?OBO0OfO TO�OxO�O�O�O�Oy2f?_  B��p,yp$QCHR�z�p@�N_`_r_�_�_�_�]c�O�_�_oo�+o?�Bc� @*d4�QqJc�D
 2o �o�o�o�o�o�o %7I[m��oa� �����c/��$PARAM_MENU ? ��  �DEFPU�LSE��	WAITTMOUT�{�RCV� �SHELL_WR�K.$CUR_S�TYL�p"�OsPT8Q8�PTBM��G�C�R_DECSN�p��������� �����-�(�:�L��u�p��������qSS�REL_ID  ���̕USE�_PROG %��z%���͓CCR��pޒ��s1�_HO�ST !�z!6�s�+�T�=���V��h���˯*�_TI�ME�rޖF��pGDEBUGܐ�{͓�GINP_FLM3SK��#�TR2�#�WPGAP� ��_�b�CH1�"�TYPE�|�P����� ���0�Y�T�f�x� �ϜϮ���������� 1�,�>�P�y�t߆ߘ� �߼�����	���(��Q�L�^�p��%�WO�RD ?	�{
 �	PR�p#�MAI��q"SU�d���TE��p#��	91���COLn%��!���L�� !���F�d�TRA�CECTL 1�v �q �_� �#��|��_�DT Q� ���z�D � _� K`�� c`��_`���������� 1CUgy� ������	 -?Qcu��� ����//)/;/ M/_/q/�/�/�/�/�/ �/�/??%?7?I?[? m??�?�?�?�?�?�? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�[��_�_�_�W��� oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�.�oP�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
.@Rdv ������� *<N`r�� �����//&/ 8/J/\/n/Dϒ/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6 HZl~���� ���� �2�D�V��h�z����������$�PGTRACEL�EN  ��  ������Ά_UP �/����������΁_CFG7 ���烸�
���*�:�D�O�|��O�  �O���DEFSPD ���������΀H_CONFI�G ���� U����dĔ�݂ ��ǑP^�a�㑶���΀IN�T�RL ��=�8l^���PE��೗���*�ÑO�΀WLID���	T��LLB 1ⳙ� ��BӐB94��O� 䘼�����Q� << ��?���� ���M�3�U���i��� ������ӿ��	�7�T�Ϣk�b�tϡ������������S�GRoP 1爬����@A!���4I����A �Cu��C�OCj+VF�/��Ȕa�0zي�ÑÐ�t��ޯs���´�ӿߨ�B������������A�S�&�B34��_������j ���������	�B� -���Q���M�������  Dz����.��� ��&L7p[� �������6!Zh)w
�V7.10bet�a1*�Ɛ@��*�@�) @��+A Ē?���
?fff>�����B33A��Q�0�B(���A���AK�� h����//'/9/P�p*�W�ӑ��n/�/�%���R�fh����*� ��P2�LR��/�/�/ �/�/H?�Ĕ�I�u�&:���?��x?�?`A���P!\3 Bu�3B��?�5BH�3[4���o��4��[45��/B\3x3Dx��?YO�?aOkO}O�< <�R@��O�C�O�O�O��O�DA�X�KNOW_M  Z�%�X��SV 賚 ڒ]��_�_�_?�_@�_�_o����W�M+�]鳛 ��	@�?3#���_�o��\A��
]bV4�@u��u��e�oX�l,�X�MR+��Jm�T3?��W�1C{�O�ADBANFWD�L_V�ST+�1 15����P4C�� �[��i/���� �?�1�C���g�y��� �����ӏ�*�	�� `�?�Q�c��w2�|Va�up�<ʟ���pA3��Ɵ؟Ꟃw4��+�=��w5Z�l�~����w6����ѯ㯂wA7 ��$�6��w8S��e�w����wMAmp������OVLD  ��yo߄r�PARNUM  ��{+þ�?υqSC-H�� �
��X�8��{s��UPDX�)�����Ϧ�_CMP_0@`���p|P'yuԿER_CHK����yqbb3��.�RqSpp?Q_MOm��_}ߥ�_RES+_G�p쩻
�e� ����0�#�T�G�x�k� }��������������׳��������� :�Y�^���Y�y����� �Ӭ������������� ��R�6UZ��॰u����V 1��FvpVa@k��p��THR_IN�Rp��(byudM�ASS Z)M�NGMON_QUEUE �u�yvup\!��N�U�Z�NW��END8��߶EXE�����BE���OP�TIO��ۚPR�OGRAM %�z%��~ϘT�ASK_I��.O?CFG �z+ϼn/� DATACc�֪+�0�A+ 2 �??/?0A?S?]51 s?�? �?�?�?�6p1�?�?�?�O"O,F�!INFO
Cc��-��bdlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_@�_�_�_�/A@FD��,c 	��!��K_�!��)fN!fENB���0m��Pf2YokhG��!2�0k X,�		d�=���&�o���e�a$�pd���i�i�g_EDIT ��/%7�����*SYSTE�M*upV9.40�107 cr7/2�3/2021 �A��Pw��P�RGADJ_p ? h $X[�p_ $Y�xZ�x�W�xқtZқtSP�EED_�p�p$�NEXT_CYC;LE�p���q�{FG�p ��p�ALGO_V ��pNYQ_FRE�Q�WIN_TYuP�q)�SIZ1�O�LAP�r!�[���M+����qCRE�ATED�r�IF�Y�r@!NAM�p�%h�_GJ�STA�TU��J�DEBU�G�rMAILTI:����EVEU���LAST�����tE�LEM� � ?$ENAB�rN��EASI򁼁AX;IS�p$P߄������qROT_R9A" �rMAX ��qjE��LC�AB
�y��C D_LVՁ`�BAS��`�1�{�r��_� ��$x����RM� RB�;�D�IS����X_SP8o�΁�� �t�P�� | 	� �2 \�AN�� �;������Ӓ�� �0�P�AYLO��3�V�_DOU�qS���p�t�PREF� ( $GRID��E
���R���Y:� ��OTOƀ�q�  �p��!��p��k�OXY�� � $L��_�PO|�נVa�S�RV��)���DI?RECT_1� �U2(�3(�4(�5(��6(�7(�8�  W�PF��A�� �$VALu�G�ROUP����qF��� !���@!�������R#AN泲���R��/���TOTA��F���PW�I=!%�REGEN#�8���@����/���ڶnTz�����#�_S����8��(�V[�'���4���G#RE��w���H��D�܅���V_H��DAuY3�V��S_Y��Œ;�SUMMAR���2 $CONFIG_SEȃ8���ʅ_RUN�m��C�С�$CMPR:��P�DEV���_�I�ZP�*��q���ENHANCE*�	�
���1�N��INT��qM)b��q�2K����OVmRo�PGu�IX��;���OVCT�����>v�
 4 ����|a˟��PSLG"�>� \ �;��?�1���SƁϕc�U�����Ò��4�U�q]�Tp�G (`�-��rJ<��O� CK�IL_M�J���VN�+��TQ�n{�N5���C�U�LȀD�V(�C6�P�_�຀@�MW�V1VV�V1d�2s�2d�U3s�3d�4s�4d� �'�	�������p	�{IN	VIB1qp�1� 2!pq/,3* 3,4 4,�p ?��;��A���N��������PL��TO�Rr3�	��[�S{AV��d�MC_FOLD ?	$SL�����M,�I��L�� �pL�b��KE�EP_HNADD�	!Ke�UCCOMc�k��
�lOP���pl\��lREM�k���΢���U��enkHPW� K�SBM��ŠCOLLAB|�Ӱn��n��+�IT�O���$NOL�FCALX� �DON�r����� ,��FL|���$SYN�y,M�C=����U_P_DLY�qs"�DELA� ����Y�(�AD��$TA�BTP_R�#��QSKIPj% ����OR� �6�� P_��� �)�� �p7��%9��%9A�$: N�$:[�$:h�$:u�$:t��$:9�q�RA��� X�����M}B�NFLIC]���0"�U!�o���NO�_H� �\�< _S�WITCHk�RA_PARAMG�O ��p��U���WJ��:Cӣ�NGRLT� OO�U���p��X�<A��T_Ja1�F�rAPS�WEI{GH]�J4CH��aDOR��aD��OO��)�2�_FJװ���saA�AV��C�HOB.�L.�l�J2�0�q$��EX��T$�'QIT ��'Q�pG'Q-�G���RDC�m" �# ��<��
R]��
xH���RGEA��84��U�FLG`g�̉H��ER	�SP9C6R�rUM_'P��2TH2No��@Q� 1 @E�D����  D� �وIi�2_P��25cS�ᰁ+�L10_CI��p
f� �pk����U ՖD��zaxT�p�Q(�;a��c��޲+��i���e��` P>`DESIGRb$�VL1:i1Gf�c�g;10�_DS��D��Xp
`FPOS11�q l�pr��xL1C/#AT�B��9U
WusIND��}��mqCp�mq`B	�HO[ME�r >u2GrM_q����!
@s3Gr��� �P�$�`!@s4GrG��Y�k�}�������?t5Grď֏�����W �?t6GrA�@S�e�w�������7Gr��П������w8Gr;�M�_�q���䕯6�S �q    �@sM��P6��<K@��! T`M�L�M�IO��m�I��:2�OK _OPy���� »Q�2�pWEG" 7�x EQA�E � #s%Ȳ$wDSBo�GNA�b�� C�P2�BS2;32S�$ �iP��9xc�ICE<@%�cPE`2� @IT���P�OPB7 1�FLOW�TRa@2���U$�CUN��`�AU�XT��2Ѷ�ERFSAC3İUU�^`�``SCH��% t�<_9�EЎA$�FREEFROM�Ц�A�PX q�UcPD"YbA�PT.�FpEEX0����!��FA%bҬ��RV��aG� &  �C�E�" 1�AL"�  �+�jc'��D��  2& �S�\PcP(
  �$�7P�%�R�2� ��T��`AXU���DSP ���@�W���:`$��RANP�%�@����K���_MIR�����MT��AP���P"�qD�QSYz�������QPG7�BRKH����ƅ AXI�  ^��i���1 <����BSOC����N��DUMMY1�6�1$SV�D�E��I�FSPD_�OVR79� DL����OR��֠N"`b��F_����@OV��;SF�RUN��"1F0�����UF"@G�;TOd�LCH�"�%RECOV��9@�@W�`&�ӂH��:`�_0�  @�RT�INVE��8AOF�S��CK�KbFWD�������1B��TeR�a�B �FD�� ��1= B1pBL@� �6� A1L�V�� Kb����#��@+<�AM:��0��j���_M@ ~�@h���T�$X`x ��T$H�BK���F��A�8����PPA�
���	������DVC_DB�3@pA�A"��X1`�X3`��Se@�`�0��qUꣳ�h�CABPP 
R�S #��c�B�@|���GUBCPU�"��S�P�`R��11�)ARŲ�!$HW_CGpl�11� F&�A1Ԡ@8p�$U�NITr�l e A�TTRIr@y"��C3YC5B�CA���FLTR_2_FAI������2bP���CHK_��SCT6��F_e'F_o,�"Ɓ*FS�Jj"CH�A�Q�'91Is�82RSD����1����_Tg�`� i�E)M�NPMf�T&2 �8p&2- �6DIA�GpERAILAC4NTBMw�LO@�Q���7��PS��� X� ��PRBSZ`J�`BC4&�	���FUN5s��RI�N�PZaߠ�07Dh�RAH@���`� `C�@��`C�Q�CBLCURuH�DA�K�!�H�HDAp�aA�H�C�ELD������C��jA�1�CTIBUu��8p$CE_RIYA�QJ�AF P��>S�`DUT2�0C���};OI0D�F_LC�H���k�L�MLF�aHRDYYO���RG�@HZ0���ߠ�@�UMULS�E�P�'3iB$�J��J����FA�N_ALM�dbW{RNeHARD�$�ƽ�P��k@2aN�dr�J�_}�AUJ �R+4�TO_SBR��~b�Іje 6?A��cMPINF��p{!�d�A�cREG榣NV��ɣZ�D��N�FLW%6r$M@�@� ��f� �0 h6'uCM4NF�!�ON	 e!e#�(b*r3F�3	�	 ���q�)5�$�$Y��r��u�_��p*o$ �/�EG������qAR��i����2�3�u�@<�AXE��ROB��RED&��WR��c�_���CSY`��q� ?�SI��WRI���vE ST�հ�ӭ d���Eg!D���t8��^a��B����9�3� OTOr�a����ARY��`ǂ�1�����FIE�~��$LINK�Q�GTH��T_4������30����XYZ���!*�O�FF�����ˀB��,Bl���e���m�FI� ��C@I�4��,B��_J$�F�@����S`����3-!�$1�w0���R��CL��,�DU���3�P.�3TUR`XS.��Ձ�bXX�� ݗFL��d���pL�0���3y4���� 1)�%K��M�5�5%8B'��ORQ�6�� fC㘴��0B�O;�D��,������a�OV	E��rM�����s2� �s2��r1���0���0�g /�AN=!�2�DQ �q���q�}R�*���6����s��V���ER��jA	�2E��.�C��A���0��XE�20Ӈ�A��AAX��F� �A�N!�SŴ1_��Q _Ɇ�^ʬ�^ʴ�^��0 ^ʙ�^ʷ�^�1&�^� �P[ɒPkɒP{ɒP�� �P�ɒP�ɒP�ɒP�ɀ�P�����ɪ �R>�D7EBU=#$8ADc0�2����
�AB�7�����V� <" 
 ��i�q��-!��%��� ���׬��״����1�� ���׷�JT��DR�m�LAB��ݥ9 FGGRO� ݒ=l� B_�1�u���}��`�����ޥ��qa��AND�����qa� �Eq��1��A@��� �NT$`��c�VEL�1��m��1u���QP��m�NA[w�(��CN1� ��3줙� �SERVEc���p+ $@@d@���!��PO
�� _:�0T ! ����p,  $.TRQ�b
(�2 -DR2,+"P~�0_ . l"@�!�&ERR��"Ip� q���~TOQ�����L�p]�e���0G���%�����R}E�@ / ,��/I -��RA� �2. d�&�! 0�p$�&��2tPM� OC|�A8 1  p�COUNT�� ��qFZN_CFG�2 4B �f�"T��:#��Ӝ� x��`�s3 ���M:0�R�qC@��/�:0��FA1P��?V�X������r���� �P:b��HEL�pe4 5���B_BAS�cRSSR�f @�S�!�QY 1�Y 2|*3�|*4|*5|*6|*72|*8�L!RO������NL�q �AB����0Z ACK��I-NT_uUS`�Pta9_PU�>b%ROU��PH@�h9#��u`w�9�TPFWD�_KAR��ar R�E���PP��A]@QUE�i&��	�f�>`QaI`��9#�j3r��f�SEME��6��PA�STY4SO�0�DI'1�`���18�rQ_TM�cM�ANRQXF�EN�D�$KEYSWITCHj31:A��4HE	�BEATmM�3PE�pLE�(�1��HU~3F�42�S?DDO_HOM�BPO:a0EF��PARr��*�v�uC�@�O�Qo �OV_Mtϒ��Eq�OCM��d�7� �8%HK�qG5 D��g�Uj��2M�p�4R��FO�RC�cWAR����p8%OM�p 6� @�Ԣ�v`U|�P��p1�V'p�T3�V4���	#O�0L�R7<��hUNLOE0h-dEDVa ���@�d8 <pAQ9�>l1MSUPG�Ua�CALC_PLA5Ncc1��AYS1�1�, �@�9 � X`��P �q;a�� ��w��2��j�M$P��`���fyt$��rSC�M�pm�q ���aq���0�tYzZzEU�Q�b�� T!�Hr�p�PvNPX_AS�f: 0g ADD|��$SIZ%a�$VA��MULTIP�"]pq�P�A�Q; � A$T9op�B���rS���j!C~ �vFRIF��2S�0�YT�pN=F[DODBUX�B�0�u&�!���CMtA������������\|Z ��< � �pƛTEg�����$SKGL��T��X�&{𷃥㰀��STMT<e�ЃPSEG�2���BW���SHOW�؅�1BAN�`TP�O���gᣥ���������V�_G�= ��$PC���O�kFB�QP\�SP�01A&0^� VDG���>� �cA00�����P���P��P�P���P��5��6��U7��8��9��A�� �P���P��w᧖��!F����h���1��v�Th�י1�1�1��U1�1�1%�12�U1?�1L�1Y�1f�U2��2��2��2ʙU2י2�2�2��U2�2�2%�22�U2?�2L�2Y�2f�U3��3��3��3ʙ3י3�3���Ȫ�3�3%�32�3�߹3L�3Y�3f�4���4��4��4ʙ4�י4�4�4��4��4�4%�42�4�߹4L�4Y�4f�5���5��5��5ʙ5�י5�5�5��5��5�5%�52�5�߹5L�5Y�5f�6���6��6��6ʙ6�י6��6�6��6��6(�6%�62�6�߹6L�6Y�6f�7���7��7��7ʙ7�י7��7�7��7��7(�7%�72�7*߹7L�7Y�7f�OR�V�`_UPD��?s �c 
������@ x $gTOR�1T�  �caOP �, ZQ_7�RE^��� J��S�sC�A��_Ux�p�7bYSLOA"A � �u$�v���w�@���@��bVALUv10�6�=F�ID_L[C:�HI5I�R$FI�LE_X3eu4$��CQP�SAV��B� hM �E_BL�CK�3�ȁ�D_CPU��p��p5�hz�pY��R3R �C � PW���� 	�!LAށ�SR�#.!'$RUN�`G@%$D!'$�@ G%e!$e!'%HR03$؇ '$��T2Pa_L}I�RD  � �G_O�2�0P_�EDI�R@�T2SPD�#E�"i0�ȁ�p	� �DCS�9@G)F � 
$JPC71q�� �S:C;C9$7MDL7$5P>93TC�`@7UF�@?89S� ?8COBu �@Q�"|�L�G�P;�;� 9:; }� ABUI_�!�L�HGb�% F\B3G$�3A�s�R�LLB_AVA�I�BPP�3�!��I� $� SEL� N�Ẽ�@RG_D Nܙ�Ta���4SC��PJ �1/ABb�PT�R`�1_M]`�L�K \M f/QLI_��FMj��PGi��U9R�6��PS_J�P\� �p�EE7B��TBC2�eL a���``�`b$�!�FT�P'T�`TDCg�� BPLp�sNU&;WTH��qhTg�tWR�2$�pERVE.S�T;S�Tw�R�_ACkP MX -$�Q�`.S�T�;S�PU@�`IC�`L�OW�GF1�QR2�g�`��p�S�ERTIA�d^0iP�P�EkDEUe�LAC�EMzCC#c�V��BrpTf�edg�aTCqV�l�adgTRQ�l �e�j|�Scu��edcu�!J7_ 4J!��RSe@qde�Q2�0`���1�PRcuPJKlvVK<�~qcQ~qw�sp�J0��q�sJJ�sJJ�sAAL�s�p�s��p�v���r5sS�`N�1�l�p�k�`5dXA_�́0QCF�BN{ `M GROU (��bh�NPC0sD�?REQUIR�R� GEBU�C�Q�6g0 2Mz��Pd�Q�SGUO�@�)A�PPR0C7@� 
u$� N��CLO� "ǉS^U܉Se
Q�@]A�"P �$PM]Pp�`�`sR�_MGa!�C���+��0�@,��BRK*�NOLD�*�SHORTMO��!m�Z��JWA�SP �tp`�sp`�sp`�sp`P�sp`�A��7��8sQ�!�QTQ� �m��R.Q�cQ�PATH�*� �*��Xh&���P�NT|@aA�"p��� �IN�R�UC4`a��C�`U%M��Y
`�)p���>�Q��cP���p��P�AYLOAh�J2�L& R_Am@�L� �����+�R_?F2LSHR�T/�LO���0���>���ACRL0z�p�y�ޤrsRH5b$H+�^��FLEX����JVR P��_._Е_�_QJ�US :�_�Vd`0�G���_tQd`�_�_lF1 G��ũ�o0oBoTofoxo��E�o�o�o�o�o �o�o ����wz3 lt����3EWF�^z	T!��X�'qju� �uu~�W؁���p �u�u�u�u����s 	��(�T �P`5�G�Y�' AT��l�pEL0�_B��s��J�Sz�JEW�CTR7B`NA��d�HAND_VB��Q��TUO@`4+�`TSW�=A��A�V� $$M��e G�AV�Qs�De�oAA���@�	$�A5�G�A�U�Ad�� 6��G�D*U�Dd�PD�G/ -CSTI�5V�5Ng�DYF ��+�x��� �P&�G�&�A��lw�o�Q�k�P������ʕ�ӕܕ�RJUWc 7 �� ��x3%�?!ASYMT��m�T�V�o�A�t�_SH�~�������$����Ưد�J�񬢐�#39"���_�VI��`8�q0V_UNIrS�4��.�Jmu�2��2A��4X� �4�6a�pt�������D&E_�������E���CH( X �̱���TOc�P�P�VsSvD�US�RU�P�����z@�D�A}@_5�U��P�EyAa���RPROG_NA���$�$LAS9T���CANs�IS~z@XYZ_SPu�@�DW]R@Ͱ,VSV@��E1QENc��DCU�R�H����HR_TF��YtQ9SЄd��O�T�uP?�SZ ��I�!A�D ���Q���#�S����#��3�vP [ � -ME�O��R4#B�!T�PPT0F@1�a��̰� h�1a%iT0� $DUMMY1���$PS_��RF���% $lfװFLA*�YP�bc$GLB_TI ��U�e`ձ#�LIF�(!\����g`OqW�P��eVOL#q�b �a_2��[d2 �[`����b�P�cZ`�TC��$BAUYDv��cST��B�2�g`ARITY0sD�_WAItAIyC,J2�OU6�ZqyyTLANS�`�{S��SZc��BUF_��r�fиx�PyyCH�K_�@CES��V� JO`E�aA<�x�bUBYT��� ��r�.�.� ��aA���M�������Q]c Xʰ����ST�����SBR@M2�1_@��T$SV�_ER�b����CL��`��A1�O�BpPG�Lh0EW(!^ 4� $a$Uq$�q$W�9�At�@R�� �Ӄ�Uم_ "��Dw$GI��}$ف ^�Ӄ�(!�` L�.��"}$�F�"E6�NEAR���B$F}��T�QL���J�@R� �a7�$JOI�NTa�o�&ՁMS�ET(!b  +�Ec�2�^�Se�҄^�(!_c�  ��U��?���LOCK_�FO@� �PBGLmV��GL'�TE�@sXM���EMP���:�K��b�$U�؂a�2_���q��`<� �q�^��C�E/�?��� $KA�Rb�M�STPDRqA܀����VECX������IUq�av�H=E�TOOL����V��REǠIS3d��6��ACH̐�m b^QONe[d3����IdB�`@$R�AIL_BOXE:a���ROB�@D��?���HOWWA�R0Aa�i`-�ROLMtb��$�*���T��`ܱ���O_FU�!>��HTML58QS��� e�`ӂ�(!dF��
��@�(!e�x��������Ӄ�}p(!f t��m�^`a��t��B�PO�%�AIPE�N����O����q��AOR�DED�m �z�XIT`��A)mSP�O�P g D �`OB�����ǯ�Ucp�`��� ��SYS��ADR��pP`U@^ � h ,"��f$A��E��E�Q�PVWVA�Qi� � �@ق�UP�R�B�$EDI|�Ad�VSHWRU�z���IS�Uq�p�ND�P7���G�HECAD�! @���!i�3KEUqO`CP)P�֗JMP��L�U R�ACE�Tj����IL�S��C��N�E���TICK�!MKQ&��H=Nr�k @���HWC��PHVF��`S�TYeB+�LO�aC����[�C�l3��
�@�F%$A��D=:��S�!$�1�p� a�e�q�ePv HVS3QU��#LO�b_1�TERC`"�T=S?�m 5���@R�m@3���ܡ��O`�	c IZ�d�A�e@ha�qtb}�hA}pP~rN��_DO�B�X�p9SSQ�SAXI�q��!v�bS�U�@TL��ƞREQ_ܠ��E�T���`�CY%��FdY'��Af\!\d�9x�P �SR$$nl-�w �@����c
�uV
Qh(�A���dC`�A��	�Y���D��p�E"�	CC�C��/�/�/	4ޣ�TSSC�` 7o h��DSmడf[`SP�@�AT� �
R��L��XbAD�DR�s$Hp� IyF�Ch�_2CH����pO����- �TU�k�Ir p�CQUCp��V��I�RAq�4���c��
K��
�^ ���Pr \z�D����|,K� P�"CN��*CƮ��!��TXSCREE��s�Pp@�INA˃<�4�DmQ����`t Tᫀ�b�� ��O Y6���º�U4h�RR�������R1�UvÐUE��u �j ��qz`Ś��RSML��U����V�1tPS_��6\��1�9G�\���C��2@4 12��0Ov�R���&F�AMTN_FL�*�`Q��W� ��PB�BL_/�WB`�PwS ����BO ��B�LE"�Cg�R"�DR7IGHtRD��!OCKGRB`�ET��|�G�AWIDTHs@���RB��a�r�0I��sEYհRx d��ʰ�����`y�BACCK���>U���PsFO��QWLAB��?(�PI��$�URm�~Ph�P�PH�y1 y 8 $�PT_��,"�R�PRUp�s5�da��Q)O%!t�zV�ȇ�p�U�@�SR ���LUqM�S�� ERVJ��SP��T{ � " GE�Rh� ��&��LPAeE��)^g�lh�lh�ki5ik6ik7ikpP`@�Z�x����$u1���p�Q zQU{SRل| <z�b�PU2�a#2�FOO .2�PRI*m9�[��@pTRIPK�m��UNDO��}�)���Yp��y��� q�h����p ~�R\p�qG ��T����-!�rOS2��vR ��2�s�CA��X���r`� �sUIaCA����3Ib_�s�OFFA�D@���Ob�r���L�t��GU��Ps�������+QSUB`� }��E_EXE���VeуsWO� e�#��w��WAl��p΁fP
 V_CDB���pT�p�O�V░���3OR�/�5�RAU@6�T�K���__����s |j �OWNj�>34$SRC�0`����DA���_MPFqI����ESP��T�$0��c��g�8n�z�E!� `%�ۂr34J���COP��$`��p_���/�+�6���CT�Cہ铸ہ�D�DCS��P�4�COMp�@�;��O`�=���K�^�/��VT�q'���Y٤Z��2���@p�w#SB����2�\0˰�_��M��%!]�DI�C#��AY�3G�P�EE�@T�QS�VR�1���eQL�� a� �P�D ��f�z��f� > ���6�QA�t�b#� �L2SHAD�OW��#ʱ_UNgSCAd�׳OWD��˰DGDE#LE�GAC)�q'�V�C\ C��� Av����だm�RF0�7���7d`C2`7�D�RIVo���ϠC��A]�(�` ���MY_UBY�d?Ĳ��s ��1��$0������_ఆ���L��BMv�A$�DEY	�cEXp@C�/�MU��1X��,��0US����;p_R"1�0p#�2��GPACIN*���RG��c�y�:�`y��sy�C/�RE�R�"!�q�y�D@�S L !�G�P�"H��p�R�pD@�&P��Px1Q��	.���RmE��SWq�_Arђ�+�{�Oq�AA(/�3�hEZ�U����g n��HK����PJ��_/�Q0{�EAN��ۀ2�2�0�MRCVCA�; �:`ORG��Q��dR	��L�����REFoG�����!�+` 	�p��������<���q�_����r��� S�`C��Ú�ҁ�@D� ��0�!��#q��š�OU����?� g��Վ2�J@00� 1�*p�����0 UL�@�f�CO�0)��� NT�[��Z�Qf�af% L飏����Q��a�VI�Aچ� �ÀHD<7 6P$JO�`oB��$Z_UP|o��2Z_LOW���$�QiBn��1$EP�s�y�� 1�!f ��0æ4�� 5�PA�A� �CACH&�LO�w�В�1B�*��Cn�I#F^��qTm����$HO2�B32{��Uÿ2O�@ ���Ro��=a��Ɛ�VP���@A"_SI	Z&�K$Z$�F(�G'����CMPk*FAIjo�G��AD�)�/�MRE���"P'G�P�0е�9�ASY�NBUFǧRTD��%�$P!�COLE_'2D_4�5W�sw��~�UӍQO��%EwCCU��VEM��xv]2�VIRC�!5�#�2�!_>�*&�p�Wp��AG	9R�X#YZ@�3�W���8���4+Qz0T"��I�M�16�2P�GR�ABB�q��;�LE�RD�C ;�F_D��F�f50MH�PEP�R��0����l�JR�LAS�@��[_GEb� �H൑~23�ET����"���b¨�I�D�ҙ6m�BG�_LEVnQ{�PK�|Л6\q��GI�@N\P4�[�P��!gI�dr�S� �NRTOm�VLʁc�Ų���#a��c"!D�qDE����Xа�X����q�2��d��p�zZ���d�c���DR4q��q2pT��U&��� $�ITPr�9p[Q��ՓV�VSF$�d�  fp/�f��UR��QaMZu9�dr��ADJ`C�v� ZDVf� D�X�AL� � 4 P�ERIKB$MS7G_Q3$Q!o%����p'��dr:g�qxQ� �XVR\t���B�pT_\��R_�ZABC"�����Sr���
X�aAC�TVS' � �� $|u�0�cCgTIV�Q!IOu�s&D�IT�x�D�Vϐ
x�P��4�!���pPS����� �#��!���q!L�STD�!�  �_}ST�	 wrvq�CHx�� L-� @��u�Ɛ*���P GNA#�C�!q��_FUN��  ��ZIPu��LHR�$L����p��ZMPCF"���`bƀ�rX�ف��LN�K��
��M�#�� $ !��ބ�CMCMk�C8�C�"����P{q '$J8�2�D6!>� O�H���T���2������M���UX�1݅UXE1Ѡ��1C���Y���ੑ����˗7�FTFpG>������Z��C�s@�j���$��YD'@ � �8n�R� Uӱ$�HEIGHd�:h?(! 'v��@���� � Gd����$B% � E��SH�IF��hRVn�F�`�HpC� 3�(� 8H`O�ѡ�C��+%YD	�"�CE�pV�1}�SPHERs� � ,! M�c��u� �$POWEORFL 4Q|�����|�p�RG�`��������_�A�  ��?�p����pd��NSb �����?�  Bz|� >l�  <@�|�Z�|�%���˃���8�ŵ�� 2ӷ��� 	H`pl&����>���A� |��t$���*��/�� **:@���p�ϥ��͘���F������ɘ�� |�����5������� %ߟ�I�[߉�ߑ�� ����������w�!�3� a�W�i��������� ��O����9�/�A��� e�w�������'���� �=O}s �������k 'UK]��� ���C/��-/#/ 5/�/Y/k/�/�/�/? �/�/?�/?�?1?C? q?g?y?�?�?�?�?�? �?_O	OOIO?OQO�� 	 �O�O�O_ �E��3_���O`_�O�_��_÷PREF �Ӻ�p�p
��I?ORITY p|�d���p����pSPL`z����WUT�VqÈ�gODU~����Y�_?�OG��Gx���R��,fHIBqO�y�|kTOENT �1��yP(!A�F_b�`�o�g!�tcp�o}!�ud�o)~!�icm�0bXY�̳�k �|�)�� �����p� ���u����� �N�5�r�Y��������̏�����*/c̳�ӹ���E�W�|�>�+���F��/��4����|��,�7�A��_,  ��P�����%�|�'���Z@��h�z�����|���ENHANCE S	#�7�A9�d��<���  �,f�T�
�_�S����POSRTe�rb�@�U���_CARTR�EP�Pr|brSKS�TAg�kSLGS6�`�k����@�Unothing������Ϳ>��P�b�To��TEMPG ?isϨE/��_a_seibanm_��i_�����0� �T�?�x�cߜ߇ߙ� �߽�������>�)� N�t�_������� ������:�%�^�I� ��m�����������  ��$H3lWi ������� D/hS�w���uϪ�VERS�I�P=g  disable���SAVE �?j	2670H�705��k/!`�m//*�/ 	�(H%b�O�+�/�Se? 6?H?Z?l?z:%<�/�?4�*'_j` 1
�kX �0ubuE�?xOqG�PURGE��1Bp`�ncqWF<@�a�TӒ*fW�`]Daa��WRUP_DELAY z�f�B_HOT %?e�'b��OnER_NORMAL�HGb�O%_�GSEMI_*_i_��QQSKIP�3.��3x��_��_�_ �_�]?eo+goKo]o oo5o�o�o�o�o�o�o �o�o5GYi �}������ �1�C�U��y�g��� ������я����-��?�7%�$RACF�G �[ќ�3��]�_PARAMr�Q3y��S @И�@`�G�42Cj۠��2��CbFzB�B]�BTIF����J]�CVTMOUړ����]�DC�R�3�Y ���Q@�B���B�e@���@B�<W{B��]���1���ᑿl'����eN�߾K��_��o ;e��m���KZ;�=�g;�4�<<����f@����� �5�G�Y�k�}��������ſ׿���xUR�DIO_TYPE�  �V�5��ED_PROT_a�&g>��4BHbC�EސSǆQ2c� ��B�ꐪϸ� ��ϐ����&�ݹ� W�V_~�o����߱� ��������A�O�m� r���9������� �������=�_�d��� ������������� ��'I�Nm�� �������# EJi+k�� ����//4/F/ /g//�/y/�/�/�/ �/�/	?+/0?O/?c? Q?�?u?�?�?�?�?�?�?;?,O��S�INT� 2�I���l�G;� jO|K��鯤O�f�0 �O�K�? �O�?___N_<_r_ X_�_�_�_�_�_�_�_ �_&ooJo8ono�ofo �o�o�o�o�o�o�o" F4j|b�� �������B��O�EFPOS1 �1"�  xO��o×O����ݏ 鈃���Ϗ0��T�� x����7���ҟm��� �����>�P����7� ������W��{���� �:�կ^�������� ��S�e��� ��$Ͽ� H��l��iϢ�=��� a��υ�� ߻���� h�Sߌ�'߰�K���o� ��
��.���R���v� ��#�5�o������� ���<���9�r���� 1���U����������� 8#\����? ��u��"�F X�?���_ ��/�	/B/�f/ /�/%/�/�/[/m/�/ ?�/,?�/P?�/t?? q?�?E?�?i?�?�?O (O�?�?OpO[O�O/O �OSO�OwO�O_�O6_ �OZ_�O~_�_+_=_w_ �_�_�_�_ o�_Do�_�Aozocf�2 1 r�o.oho�o�o
o .�oR�oO�#� G�k����� N�9�r����1���U� ���������8�ӏ\� ��	��U�����ڟu� ����"����X��|� ���;�į_�q����� �	�B�ݯf����%� ����[���ϣ�,� ǿٿ�%φ�qϪ�E� ��i��ύ���(���L� ��p�ߔ�/�A�Sߍ� ������6���Z��� W��+��O���s��� ������V�A�z�� ��9���]������� ��@��d��#] ���}�*� '`���C� gy��&//J/� n/	/�/-/�/�/c/�/ �/?�/4?�/�/�/-? �?y?�?M?�?q?�?�? �?0O�?TO�?xOO�O<�o�d3 1�oIO [O�O_�O7_=O[_�O __|_�_P_�_t_�_ �_!o�_�_�_o{ofo �o:o�o^o�o�o�o �oA�oe �$6 H�����+�� O��L��� ���D�͏ h�񏌏�����K�6� o�
���.���R���� �����5�ПY���� �R�����ׯr����� ����U��y���� 8���\�n������� ?�ڿc�����"τϽ� X���|�ߠ�)����� ��"߃�nߧ�B���f� �ߊ���%���I���m� ��,�>�P������ ���3���W���T��� (���L���p������� ����S>w�6 �Z����= �a� Z�� �z/�'/�$/]/ ��//�/@/�/�O�D4 1�Ov/�/�/ @?+?d?j/�?#?�?G? �?�?}?O�?*O�?NO �?�?OGO�O�O�OgO �O�O_�O_J_�On_ 	_�_-_�_Q_c_u_�_ o�_4o�_Xo�_|oo yo�oMo�oqo�o�o �o�o�oxc�7 �[����>� �b����!�3�E�� ��ˏ���(�ÏL�� I������A�ʟe�� �������H�3�l�� ��+���O���ꯅ�� ��2�ͯV����O� ����Կo�����Ϸ� �R��v�Ϛ�5Ͼ� Y�k�}Ϸ���<��� `��τ�߁ߺ�U��� y���&�������� ��k��?���c���� ��"���F���j���� )�;�M��������� 0��T��Q�%��I�m��/�$5 1�/���mX ���P�t�/ �3/�W/�{//(/ :/t/�/�/�/�/?�/ A?�/>?w??�?6?�? Z?�?~?�?�?�?=O(O aO�?�O O�ODO�O�O zO_�O'_�OK_�O�O 
_D_�_�_�_d_�_�_ o�_oGo�_koo�o *o�oNo`oro�o�o 1�oU�oyv� J�n����� ��u�`���4���X� �|�ޏ���;�֏_� �����0�B�|�ݟȟ ���%���I��F�� ���>�ǯb�믆��� ���E�0�i����(� ��L���翂�Ϧ�/� ʿS�� ��LϭϘ� ��l��ϐ�ߴ��O� ��s�ߗ�2߻�V�h� zߴ�� �9���]��� ���~��R���v�����#�	6 1 &������������� ��}���<��` ����CUg� �&�J�n	 k�?�c��/ ���	/j/U/�/)/ �/M/�/q/�/?�/0? �/T?�/x??%?7?q? �?�?�?�?O�?>O�? ;OtOO�O3O�OWO�O {O�O�O�O:_%_^_�O �__�_A_�_�_w_ o �_$o�_Ho�_�_oAo �o�o�oao�o�o�o D�oh�'� K]o�
��.�� R��v��s���G�Џ k�􏏏���ŏ׏� r�]���1���U�ޟy� ۟���8�ӟ\����� �-�?�y�گů���� "���F��C�|���� ;�Ŀ_�迃������ B�-�f�ϊ�%Ϯ�I� �����ߣ�,���P�<6�H�7 1S��� �I��߲������� 3���0�i���(�� L���p�����/�� S���w����6����� l�������=���� ��6���V�z � 9�]�� �@Rd��� #/�G/�k//h/�/ </�/`/�/�/?�/�/ �/?g?R?�?&?�?J? �?n?�?	O�?-O�?QO �?uOO"O4OnO�O�O �O�O_�O;_�O8_q_ _�_0_�_T_�_x_�_ �_�_7o"o[o�_oo �o>o�o�oto�o�o! �oE�o�o>�� �^�����A� �e� ���$���H�Z� l�����+�ƏO�� s��p���D�͟h�� �����ԟ�o�Z� ��.���R�ۯv�د� ��5�ЯY���}�c�u�8 1��*�<�v� ��߿��<�׿`��� ]ϖ�1Ϻ�U���y�� �ϯ�����\�G߀�� ��?���c����ߙ�"� ��F���j���)�c� ���������0��� -�f����%���I��� m������,P�� t�3��i� ��:���3 ��S�w /� �6/�Z/�~//�/ =/O/a/�/�/�/ ?�/ D?�/h??e?�?9?�? ]?�?�?
O�?�?�?O dOOO�O#O�OGO�OkO �O_�O*_�ON_�Or_ __1_k_�_�_�_�_ o�_8o�_5ono	o�o -o�oQo�ouo�o�o�o 4X�o|�; ��q����B� ���;�������[� ������>�ُb������!�������MA_SK 1 ��������ΗXNO � ݟ���MOT�E  ���S�_C�FG !Z����N�����PL_RA�NGV�N������O�WER "���Ϡ��SM_DRY�PRG %����%W��եTART� #Ǯ�UME_PRO���q����_EXEC_EN�B  ����GScPDJ�������gTDB����RMп���IA_OPTI�ON������~�NGVERS���`�řI_�AIRPUR�� �R�+���ÛMT_�֐T X���ΐO�BOT_ISOLEC����������/NAME8��H�Ě�OB_CATEG�ϣ,��S�[�.��ORD_NUM �?Ǩ��H705  N��ߨߺ�ΐPC_T�IMEOUT�� �xΐS232s�1�$��� L�TEACH PENDAN��o���)���V�T�M�aintenance ConsN��&�M�"B�P�No Use6�r�8�������̒��N�PO$��Ҏ�"�^��CH_LM�Q�朕	a�,�!U�D1:��.�RՐVgAILw��粥�*�SR  t�� ���5�R_INoTVAL����� ���V_DAT�A_GRP 2'|���� D��P�������	�� ����B0 RTf����� �/�/>/,/b/P/ �/t/�/�/�/�/�/? �/(??L?:?p?^?�? �?�?�?�?�?�?O O "O$O6OlOZO�O~O�O �O�O�O�O_�O2_ _ V_D_z_h_�_�_�_�_ �_�_�_o
o@o.oPo�vodo�o��$SA�F_DO_PUL�SW�[�S���i�SC�AN�������S�Cà(/��0���S�S�
������(q�q�qN� �L ^p���5��`� ��$��+�E�r2M�qqdY��P�`�J�	t/� @��������ʋ|���� r ք��_ @N�T ��'�9��K�X�T D�� X���������ɟ۟� ���#�5�G�Y�k�}��������䅎������Ǧ  "�;�oR� ����p"�
�u���Di���q$q�  � ���uq %�\�������ҿ��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6�H�Z����珈��� ����������g�;� D�V�h�z��������� ������(�Ӣ0�r� i�y���$�7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/?r�+?=? O?a?s?�?�?�?�?�? 8��?OO'O9OKO]O oO�O��$�r�O�O �O�O	__-_?_Q_c_ u_�_�Y�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o�o "4FXj|�c�路g������ �0�B�T�f�x�����@����ҏ�������:�Ҧ��y��3�	�	1234�5678��h!�B!�� \��p0���� Ο�����(�:�@� �c�u���������ϯ ����)�;�M�_� q�����R���ɿۿ� ���#�5�G�Y�k�}� �ϡϳ����ϖ���� �1�C�U�g�yߋߝ� ����������	��-� ��Q�c�u����� ��������)�;�M� _�q���B�������� ��%7I[m �������� !3EWi{� ������// //�S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?D/�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O*����O	_�E�?5_G_�Y_�yCz  A}��z   ��x�2�r }��)�
�W�/  	�*�2�O�_��_ oo"l�#\� �_hozo�o�o�o�o�o �o�o
.@Rd v����Mo�� ��*�<�N�`�r��� ������̏ޏ����&�8�J��X #P$P�Q:�R<u� k��Q?  �������S�P���Q�Qt C �PÙ۟�P(� `,b����]�P�Fl�$SCR_G�RP 1*0+�04� �� �,a ��U	 v��~������d����%���ɯ���h]���P�D1� �D7n��3��Fl�
CRX-10i�A/L 2345_67890�Pd�i r��Pd�L ��,a
1o�������-�[ ¶~�+fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@�R��d�t���H�~�Ă�m��ϴ��� ���ϼ��,a��1�P��U�[�G�imXhuP�,[��	ӛ�B�  BƠߞҷԚ�9A�P��  @1`��暡@����� ?����H����ښ�F?@ F�`A�I� @�m�X��|����� ������������:�0%�7�I�[�B�i��� ��������������- Q<u`��En �ٯ���W�P�"+f@_�5��1`b���x����ͣ�O�,dA����ߒ��Fa�,a ��#!"/4/E-!pZ(f/x/G/ (�P�!(� �/�/�/��/�/?#9b����S7�س�M�ECLVLw  ,a��ݲ��Q@f1L_DE�FAULTn4b1��1`�3HOTSTR�=��2�MIPOWERF�m0pU�5�4WF�DO�6 �5L�E�RVENT 1+�u1u1�3 L!DUM_EIP#?�5H�j!AF_�INE�0SO,d!�FT)O�NIO�O!����O ��O�O!�RPC_MAI�N�O�H��O>_SV�IS_�I�-_�_!OPCUf�_�W�y_�_!TP&�PPU�_<Id�_"o�!
PMON_POROXY#o?Feo�no�R<o8Mf]o�o!�RDM_SRV�o<Ig�o!RȠ�"=Hh�oR!
�PM�o9LiA�!RLSYNC���y8��!R3OS(O��4�6��!
CE�PMTC�OM7�?Fk%���!=	K�CONS��>G�lq�Ώ!K�WA'SRC�o?Fm���;!K�USB�=H�n	�f�!STM�0��;JoU����O֟��c����CICE_�KL ?%K �(%SVCPR#G1��G�1�2G�L�"6�3o�t�6�4����"6�5��į6�6��6�7��6���W�R�	9_�d�3���6� 9���6�a�ܿ6���� 6���,�6�ٯT�6�� |�6�)���6�Q���6� y���^����^�ʿD� ^��l�^�ϔ�^�B� ��^�j���^����^� ��4�^���\�^�
߄� ��2���6��/��� �V��<�'�`�K��� o������������� &J5nY�� ������4 F1jU�y�� ���/�0//T/ ?/x/c/�/�/�/�/�/ �/�/??>?)?P?t?�_?�?
�_DEV �I�MC�:�84���4GRP 2/E�0+��bx 	� W
 ,@�0
�?OD!OKODdOvO ]O�O�O�O�O�O�O�O _�O_N_5_r_Y_�_(�_/CE�0�_�_ �_o�_'ooKo]oDo �oho�o�o�o�o�o�o��o�o5Y�_D�0i@���� ��� �=�$�a�s� Z���~��������؏ �lD�Q9O'�	A�~�1O������ן
� ������U�<�y��`�������ӯ*�B	 ����3���W�>�P� ��t��������ο� �/�A�(�e�Lωϛ� 6���v��_�ϐ����� ���'߅�v�]ߚ߁� ���߷������*�5� N��r������� �������&�8��\� C���g�y��������� ��g�4-jQ �u����� B)fx_� ���)��/,/ /P/7/t/[/m/�/�/ �/�/�/?�/(??L?�^?E?�?�7d �[~
�6 s���A;*=� �6?�=���D��>�����g�:�0��ī���|@�-�@��5_�eA�5�-�=BG+h��&���6)A�B�m�����`x��=�?7O%TELEOP8O�cN[~y��5��o�ʾTF������������|��ҝ�����E�1��E@�*�A`��~�n�!��$��A���M�Y�<T�������C=�J�?���Gc��McO���IJO/_�[~���6r _�1<��׻��y;��	A`�ʛ1�bP��N	V�A��&@в@�?��@)E�]�1������0ד�� x���Q���U?�Q���O�__ _oDU��NU9��6>�ߔ�E�bQ�2�]�j_ ���rAS�AT��@��@G$��_ ��yC�� �Pr}��Q� 2i?�R�_`�o�_�_�oDU�K�5���l�������S���`
��� 3>v����M@�@�V��@�%@���Ŀ�q���]�V�N��N�!C�(uµ���� �®��ɒow�o�o�DU��b�5?���T�@O�P�%��*�-�����N�PA�����
Q@����q�A����M�{�B&��br'C9r�t�1��^с�fK��������pm�5>���@�«��͙~��E�A�����c�N'pA(��AC8AD�����A��y�Nd�A���R��ֺ������s��`_��^��\�n�S�BW�c��v"��?/����H?��4@� �+79���$ΏA8	�AAlܾc`��f�@�c+�Ne�?6A�z2���LQ� f��t?���`�D��p2�D�)�DT�m��6�M�W�1�������F0�<
u���8�N�W`@�^}A1N�u@X�ƿP��A%��N�j�!��g(�E��uB��y�!F�`G�/������:�p��6
������\��w�������kuf�@�In_�PI3��@K�@�"����P������NuN�A���Q¸!C=�������º�����ٯ�п;�t2��0�Bq̾���?P�������lG-���~�u�AR���@&G Az����:�AX����NzQBA������V�����uC���׿�����ϒ��I �I����������*�P�%���y�hoR߬� ���߾������Z�?� ~��r������� ����2��V���J�8� n�\�~�������
��� .���"F4jX z������� B0f��� VxR���// >/�e/�./�/�/�/ �/�/�/�/?X/=?|/ ?p?^?�?�?�?�?�? �?0?OT?�?HO6OlO ZO�O~O�O�?O�O,O �O __D_2_h_V_�_ �O�_�O|_�_x_�_o 
o@o.odo�_�o�_To �o�o�o�o�o< ~oc�o,���� ����V;�z� n�\���������ڏ� ��ʏ�Ə4�j�X� ��|����ٟ���� ����0�f�T���̟ ���z��ү���� �,�b�����ȯR��� ���ο���j��� aϠ�:ϔςϸϦ��� �� �B�'�f���Z��� jߐ�~ߴߢ������ >���2� �V�D�f�� z��������
��� .��R�@�b������ ��x�������* N��u�>`:� ���&hM� �n����� �@%/d�X/F/|/ j/�/�/�/�//�/</ �/0??T?B?x?f?�? �/?�??�?O�?,O OPO>OtO�?�O�?dO �O`O�O_�O(__L_ �Os_�O<_�_�_�_�_ �_ o�_$of_Ko�_o ~olo�o�o�o�o�o�o >o#bo�oVDzh ������� ��R�@�v�d���� �� �������� N�<�r�����؏b�̟ ���ޟ ���J��� q���:�����ȯ��� گ��R�x�I���"�|� j�����Ŀ���*�� N�ؿB�ԿR�x�fϜ� �������&ϰ��� >�,�N�t�bߘ��Ͽ� �ψ�������:�(� J�p�ߗ���`���� ����� �6�x�]�o� &�H�"����������� P�5t���hVx z����(L �@.dRtv� � �$�//</ */`/N/p/���/� �/�/�/??8?&?\? �/�?�/L?�?H?�?�? �?O�?4Ov?[O�?$O �O|O�O�O�O�O�O_ NO3_rO�Of_T_�_x_ �_�_�_�_&_oJ_�_ >o,oboPo�oto�o�_ �o�o�o�o�o:( ^L��o��or� ��� �6�$�Z�� ���J�����؏Ə� ���2�t�Y���"��� z�����ԟ�:�`� 1�p�
�d�R���v��� ��Я���6���*��� :�`�N���r����Ͽ �����&��6�\� Jπ�¿���p����� ����"��2�Xߚ�� ��H߲ߠ��������� �`�E�W��0�
�x� ���������8��\� ��P�>�`�b�t����� �����4���(L :\^p���� � �$H6X ����~��� � //D/�k/�4/ �/0/�/�/�/�/�/? ^/C?�/?v?d?�?�? �?�?�?�?6?OZ?�? NO<OrO`O�O�O�O�O O�O2O�O&__J_8_ n_\_�_�O�_�_�_�_ ~_�_"ooFo4ojo�_ �o�_Zo�o�o�o�o�o B�oi�o2� �������\ A��
�t�b������� ��̏"�H��X��L� :�p�^���������ߟ ������"�H�6�l� Z���ҟ�������د ����D�2�h����� ίX�¿���Կ
��� �@ς�gϦ�0Ϛψ� �Ϭ������H�-�?� �����`ߖ߄ߺߨ� �� ��D���8�&�H� J�\��������� �����4�"�D�F�X� �������~����� ��0@������� f�����, nS���� ���/F+/j� ^/L/�/p/�/�/�/�/ /?B/�/6?$?Z?H? ~?l?�?�?�/�??�? O�?2O OVODOzO�? �O�OjO�OfO�O
_�O .__R_�Oy_�OB_�_ �_�_�_�_o�_*ol_�Qo�[�P�$SE�RV_MAIL + �U�`��Qvd�OUTPUT�h��P@vdRoV 20f  �`� (a\o�ovdS�AVE�l�iTOP�10 21�i d 6 s�P_6r _�P:p�a2o`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟�`����0�B���u�YP�cFZN_�CFG 2e��c�T�a�e|�G�RP 23��q ,B   AƠ~�QD;� BǠ��  B4�S�RB21�fHELL�4ev�`�o���/�>�%RSR>�?�Q���u����� ҿ������,��PϠ;�t�_Ϙϩ����  �¼���(�Ϸͻ��P�&Ҧ'�ސW��2�Pd���g��HK 15�� ,ߡ߫� ����������@�;� M�_���������������OMM �6��?��FTOV_ENB�d�au��OW_REG_U�I_��bIMIOFWDL*�7.�ɥ��/WAIT\�`ٞ�ȼ��`���d��TI�M������VA��`����_UNIT�[�*yLCy�TR�Y��uv`ME�8���aw֑d ���9� ���j��<��X�Pxڠ6p`?�  �`�o+=`�VL�l�fMO�N_ALIAS k?e.��`heGo ������/)/ ;/M/�q/�/�/�/�/ d/�/�/??%?�/I? [?m??�?<?�?�?�? �?�?�?!O3OEOWOO {O�O�O�O�OnO�O�O __/_�OS_e_w_�_ �_F_�_�_�_�_�_o +o=oOoaoo�o�o�o �o�oxo�o'9 �o]o��>�� ����#�5�G�Y� k��������ŏ׏�� ����1�C��g�y� ����H���ӟ���	� ��-�?�Q�c�u� ��� ����ϯᯌ���)� ;��L�q�������R� ˿ݿ��Ͼ�7�I� [�m��*ϣϵ����� �ϖ��!�3�E���i� {ߍߟ߱�\������� ����A�S�e�w�� 4����������� +�=�O���s������� ��f�����'�� K]o��>�� ���#5GY�}����l��$SMON_DE�FPROG &������ &*SYS�TEM*���R�ECALL ?}�� ( �}3�xcopy fr�:\*.* vi�rt:\tmpb�ackT!=>19�2.168.56�.1:16260� z"�/�/�/�,}4K%aS/e/w%�/?#?�5? }8L$s:o�rderfil.dat�,�/?�?�?��?}/L"mdb: �/o?| {?OO0O�$ J/�/n/ O�O�O�O�/ YOkO�/_!_3_F?X? �?�?�_�_�_�?�?q_ �?oo/oBO�O�OxO �o�o�o�O�Oco�O +>_P_�_t_�� ��_�_i�_��'� :oLo�opo�����8� �o[�m����#�5�H Z���������a� �|���1�D�׏� z�������S�e��� 	��-�@�R�۟v��� ������Пk����� )�<�N��r��ϕϧ� ��̯]����%߸� J�\�� ߑߣߵ�ȿ c��~��!�3�F��� ��|ύ�����U�g� ����/�B�T���x� ����������m��� +>�P���t�� �����_��' :�L�^����8 ��e���/#/5/H ��~�/�/�/�W/ i/�??1?DV� z�?�?�?��/o?� 	OO-O@/R/�/v/�O �O�O�/�/aO�/__ )_<?N?�?�O�_�_�_ �?�?g_�?�_o%o7n��$SNPX_A�SG 2:����Va� � b%�7o~o � ?�GfPARAoM ;Ve`a� �	lkP>T�DP>X�d� ���I`OFT_K�B_CFG  �CS\eFcOPIN_�SIM  Vk��b+=OYsI`R�VNORDY_DOO  �eukr�QSTP_DSB�~�b�>kSR �<Vi � & TELEO�e��{v>TW`I`TOP_ON_ERRx�Gb�PTN zVeP��D:��RING_PRM�'��rVCNT_GOP 2=Ve�ac`x 	���DP��яؼ���BgVD�RP' 1>�i�`�Vq ؏0�B�T�f�x����� ����ҟ�����,� >�e�b�t��������� ί���+�(�:�L� ^�p���������ʿ� � ��$�6�H�Z�l� ~ϐϷϴ��������� � �2�D�V�}�zߌ� �߰���������
�� C�@�R�d�v���� ������	���*�<� N�`�r����������� ����&8J\ n������� �"4[Xj| �������!/ /0/B/T/f/x/�/�/ �/�/�/�/�/??,? >?P?b?t?�?�?�?�?��?�?�?O�PRG�_COUNT�f9�P�)IENBe�+E�MUC�dbO_UPD� 1?�{T  
ODR�O�O�O�O�O __A_<_N_`_�_�_ �_�_�_�_�_�_oo &o8oao\ono�o�o�o �o�o�o�o�o94 FX�|���� �����0�Y�T� f�x����������� ���1�,�>�P�y�t� ��������Ο��	�� �(�Q�L�^�p����� �����ܯ� �)�$� 6�H�q�l�~������� ƿؿ���� �I�D��V�"L_INFO {1@�E�@��	 yϽϨ������?=ք?����>G�q=�>a�����3���@o��<Q�=��7� �D/  � � D1� C4 � ´j�|�-@YS�DEBUG:@�@��o�d�I��SP_PwASS:EB?�ۿLOG A��.�A  o�i�v��  �Ao�U�D1:\��}���_MPC�ݚEk�}�A�&�� �AK�SAV B��IA#��l*�i�1�SVB��TEM_TIME� 1C���@ _0  6nĦi��;�q����MEM�BK  �EA��������X�|�@� R��� ����������h�,9
�� #�@�` r�������� �@R dv�����
Le�//(/:/L/^/ p/�/�/�/�/�/�/�/� ??$?6?H?Z?��SKV�[�EAj��?�?�?V���@f]2��|�?i�  0 o� ^
:O.@R�O�O�O}N�o�� ��OBD)O_&_8_,M2�Y_�_�_�_�_�_o�U�_�_� o'o9oKo]ooo�o�o �o�o�o�o�o�o#�5GYk_?T1SVGUNSPD��� '����p2M�ODE_LIM #D��Ҋt2�p�q�E�݉uABUI_DCS H}5���0�G�0��D���|-�X�>���*���� 
��e��iđ��r�i������uEDIT I���xSCRN �J���rS�G �K�.�(�0߅SK_OPTION�и^����_DI��ENB  /�����BC2_GRP 2L���MP�C�ʓ�|BCCF2/�N���� ����F`�>�W�B�g� ��x�����կ����� ���S�>�w�b��� ������Ͽ����� =�(�a�Lυϗ�Ň�� ��������v��
�/� U�@�yߧ��`�iМ� �߰�����
���.�� >�@�R��v����� �������*��N�<� r�`������������� ��̀4FX�� |j������ �B0fTv x�����/� ,//</b/P/�/t/�/ �/�/�/�/�/�/(?? L?d?v?�?�?�?6? �?�?�?O O6OHOZO (O~OlO�O�O�O�O�O �O�O __D_2_h_V_ �_z_�_�_�_�_�_
o �_.oo>o@oRo�ovo �ob?�o�o�o�o <*Lr`��� �����&��6� 8�J���n�����ȏ�� �ڏ��"��F�4�j� X���|��������֟ ��o$�6�T�f�x��� ������ү������ �>�,�b�P���t��� �����ο��(�� L�:�\ς�pϦϔ��� �������� ��H�6� l�"��ߖߴ�����V� �����2� �V�h�z� H������������ ��
�@�.�d�R���v� ������������* N<^`r�� �����&8� \Jl����� ���"//F/4/V/ X/j/�/�/�/�/�/�/ ?�/?B?0?f?T?�? x?�?�?�?�?�?O�? ,O�DOVOtO�O�OO �O�O�O�O�O_ V4P��$TBCSG_�GRP 2O U��  ��4Q 
 ?�  __q_[_�__�_�_��_�_�_o%k8R?SQ~F\d�HTa�?4Q	 HA��}�#e>���>$a��\#eAT�̓A WR�o�hdjma�OG�?Lfg�bp�o�n�ffhf���ȼb4P|j��o*}@���Rhf�ff>�#33pa#e<qB�o+D=xrRp�qUy�rt~��H�y rIpTv�pBȺt~	xf	x (�;���f���N�`�Ю�ˏڋ����	�V3.00WR	�crxlڃ	*@��3R~t��HH�ư� \�.�]�  cC.�����8Q+J2?SRF]�����CFG T UePQ SPܚ���r�ܟ1�� 1�W�e�	Pe���v��� ��ӯ�������� Q�<�u�`��������� Ϳ�޿��;�&�_� Jσ�nπϹϤ����� ��WRq@�0�B��� u�`߅߫ߖ��ߺ��� ���)�;�M��q�\� ������4Q _���O  ���J�8�n�\��� �������������� 4"XFhj|� �����. TBxf��nO� ���//>/,/b/ P/�/t/�/�/�/�/�/ �/�/?:?(?^?p?�? �?N?�?�?�?�?�?�?  O6O$OZOHO~OlO�O �O�O�O�O�O�O __ D_2_T_V_h_�_�_�_ �_�_�_
o�_o@o� Xojo|o&o�o�o�o�o �o�o*N`r �B������ �&��6�\�J���n� ����ȏ��؏ڏ�"� �F�4�j�X���|��� ğ���֟���0�� @�B�T���x�����ү 䯎o���̯ʯP�>� t�b������������ ��Կ&�L�:�p�^� �Ϧϸ��τ������  �"�H�6�l�Zߐ�~� �ߢ����������2�  �V�D�z�h���� ���������
�,�.� @�v�������\��� ����<*`N ����x�� �8J\(� �������/ 4/"/X/F/|/j/�/�/ �/�/�/�/�/??B? 0?f?T?v?�?�?�?�? �?�?OO��2ODO��  O�OtO�O�O�O�O�O _�O(_:_L_
__�_ p_�_�_�_�_�_ o�_ $oo4o6oHo~olo�o �o�o�o�o�o�o  D2hV�z�� ���
��.��R� @�b���v���&OXO֏ 菒�����N�<�r� `�������̟ޟ🮟 ��$�&�8�n����� ��^�ȯ���گ���  �"�4�j�X���|��� ��ֿĿ����0�� T�B�x�fψϊϜ��� ��������>�P��� h�zߌ�6߼ߪ����� �����:�(�^�p�� ��R������� ����  &�*� �*�>�*��$TBJ�OP_GRP 2�U��� � ?���C�*�	V�]�Wd������X?  *���� �, �� ���*� @�&�?��	 �A������C�  D�D�����>v�>�Ϗ\? ��aG߮:�o��;�?�AT������A�<��MX�����>��\)?����8Q�����L���>�0 &�;ikG.��Ap< x� F�A�ff��v��� ):VM�.�� S>o�*�@��R�C��	���������ff�:�6/ފ?�33�B   ��/������>):�S����� �/�/@��H�%&/�/��==� <#�
*���v�;/�ڪ!?���4B�3?'?2	 ��2?hZ?D?R?�?�? �?F?�?�?�?�?OAO O�?`OzOdOrO�O�O�*�C�*���A��	�V3.00{�ocrxl��*P��%�%c5Z �F� JZH �F6� F^ �F�� F�f �F� G� �G5 G<
 �G^] G� �G���G�*��G�S G�; 7G��ERDu�\�E[� E� �F( F-� �FU` F}  �F�N F� �F�� Fͺ �F� F�V �G� Gz �Ga 9ѷ$�Q�LHefJ4�o
,b*�0c1���O�H�ED_TCH cXd�+X2S�&���&�d$'X�o�o�*�1F�TESTPARS  ��cV�HRpABL�E 1Yd�  N`*�����g$j�g��h�h)�1��g	��h
�h�hHu*���h�h�h%vRDI0n�GYk}��u	�O�#�-� ?�Q�c�u�)rS�l� �z6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z���I�� �m�Fwͩ��ȏڏ� ������x)r���NUM  ��Un���2� Ep��)r_CFG �Z��I���@V�IM?EBF_TTqD�:�e޶VER���z��޳R 1[8{O 8�o*�%�2Q� ��د  9�K� ]�oρϓϥϷ����� �����#�5�G�Y�k� }��ߡ߳��������� ��1���E�W�i�{� ������������� �/�A�S�e�w����� ����������+H=O�_���@���`LIF \&��D`����tDR�(FP
�!p��!p� d� ��M�I_CHAN� �� DBGLV�L��fETHERAD ?u
��0`1�_}��ROUT�!Ǝj!��SN�MASKY�j255.%S///�A/S�`OOLOF/S_DIp�C�ORQCTRL C]8{��1o�-T�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�?�OL�/6O%OZOcPE_DETAI7��*PGL_CON?FIG c�������/cell�/$CID$/grp1^O�O�O�O
__|���G_Y_k_}_ �_�_0_�_�_�_�_o o�_CoUogoyo�o�o ,o>o�o�o�o	- �oQcu���: �����)����_�q���������׮} N����%�7�I�a�KOq�P��M�����ʟ ܟ� �G�$�6�H�Z� l�~������Ưد� �����2�D�V�h�z� �����¿Կ���
� ��.�@�R�d�vψϚ� )Ͼ��������ߧ� <�N�`�r߄ߖ�%ߺ� ��������&��J� \�n����3����� �����"���F�X�j��|��������@��User Vie�w �I}}1234567890�� ��+=Ex �e����2��B�� ����`r��3�Oas����x4>//'/@9/K/]/�~/x5� �/�/�/�/�/?p/2?x6�/k?}?�?�?�?�?$?�?x7Z?O1O�COUOgOyO�?�Ox8 O�O�O�O	__-_�O�N_TR l?Camera���O��_�_�_�_�_�_˂E �_o)o;n��Uogoyo0�o�o�o�)  mV�	 �_�o#5GY o }���o������F_�mV=�k� }�������ŏl��� �X�1�C�U�g�y��� 2�D��"�ן���� �1�؏U�g�y�ğ�� ����ӯ�����D��k ��E�W�i�{�����F� ÿտ�2���/�A� S�e��nUY9������ ������	߰�-�?�Q� ��u߇ߙ߽߫���v� D�If��-�?�Q�c� u�ߙ�������� ��)�;���D��I�� �������������� )t�M_q���N�`�93�� 0B��Sx�1 �����//�J	oU0�U/g/y/�/ �/�/V�/�/�/�? -???Q?c?u?/./tP v[?�?�?�?OO(O �/LO^OpO�?�O�O�O �O�O�O�?oU�k�O:_ L_^_p_�_�_;O�_�_ �_'_ oo$o6oHoZo _;%N��_�o�o�o�o �o �_$6H�ol ~����moe�� ]�$�6�H�Z�l� �������؏����  �2��e&�ɏ~��� ����Ɵ؟���� � k�D�V�h�z�����E� e��5����� �2� D��h�z���ׯ��¿�Կ���
ϱ�  ��9�K�]�oρϓ���Ϸ���������   ��5�G�Y�k� }ߏߡ߳��������� ��1�C�U�g�y�� �����������	�� -�?�Q�c�u������� ��������);pM_q�  
���(  �-�( 	 ����� ��#35G}�k����
� �Y�
//./��R/ d/v/�/�/�/����/ �/�/A/?0?B?T?f? x?�/�?�?�??�?�? OO,O>O�?bOtO�O �?�O�O�O�O�O_KO ]O:_L_^_�O�_�_�_ �_�_�_#_ oo$ok_ HoZolo~o�o�o�_�o �o�o1o 2DV h�o�o���	� �
��.�@��d�v� �������Џ��� M�*�<�N���r����� ����̟�%���&� m�J�\�n�������� ȯگ�3��"�4�F� X�j�����������ֿ �����0�w���f� xϊ�ѿ���������� �O�,�>�Pߗ�t߆� �ߪ߼�������� ]�:�L�^�p������@ ������������ ��"f�rh:\tpgl�\robots\�crx!�10ia?_l.xml��D� V�h�z�������������������0B Tfx����� ����,>Pb t������� �/(/:/L/^/p/�/ �/�/�/�/�/��/? $?6?H?Z?l?~?�?�? �?�?�?�/�?O O2O DOVOhOzO�O�O�O�O �O�?�O
__._@_R_ d_v_�_�_�_�_�_�O �_oo*o<oNo`oro��o�o�o�o�o�n ��6� ���<<w 	� ?��k !�o;iOq� �������� %�S�9�k���o������я����(�$T�PGL_OUTP�UT f����;�� �&� 8�J�\�n��������� ȟڟ����"�4�F� X�j�|�������į��p�ր2345678901���� �1�C�K����r��� ������̿d�п��&�8�J��}T�|ώ� �ϲ���\�n����� 0�B�T���bߊߜ߮� ����j�����,�>� P����߆������ ��x����(�:�L�^� ��l�����������t� ��$6HZl z�������  2DVh � ������/./ @/R/d/v//�/�/�/��/�/�/�/ۂ $$��ί<7*?\? N?�?r?�?�?�?�?�? �?OO4O&OXOJO|O nO�O�O�O�O�O�O_�O0_"_T_}�an_�_ �_�_�_�_�]@�_�o	z ( 	 V_Do2ohoVo�ozo �o�o�o�o�o
�o. R@vd��� ������(�*��<�r�`���ܦ�  <<I_ˏݏ �������:�L�֪ ��}���)���ş���� ���k��C�ݟ/�y� ��e������������ �-�?��c�u�ӯ]� ����W���Ϳ��)� ����_�q��yϧρ� ������M��%߿�� [�5�Gߑߣ�߫��� s����!���E�W�� ?���9�������� �i���A�S���w��� c�u����/����� =)s���� �U���'9 �!o	[��� ��K�#/5/�Y/ k/E/w/�/�/�/�/ �/�/?�/?U?g?�/ �?�?7?�?�?�?�?	O�O��)WGL1�.XML�_PM�$�TPOFF_LI�M ���P��{�^FN_SVf@�  �TxJP_�MON g���zD�P�P2ZIS�TRTCHK �h��xFk_aBVT?COMPAT�HQ�|FVWVAR �i�M:X�D R�O R_�P�BbA�_DEFPROG� %�I%T�ELEOPi_�O_DISPLAYm@��N�RINST_M�SK  �\ ~�ZINUSER_��TLCKl�[QU?ICKMEN:o�ToSCREY`��~Rtpsc�T�at`yixB�`_�iS�TZxIRACE_�CFG j�I�:T�@	[T
?�~�hHNL 2k�Z���aA[ gR-?Q�cu����z�eI�TEM 2l{� �%$1234?567890 ��  =<
�0�B�J��  !P�X�dP ���[S���"��� X�
�|���W���r�֏ ����.��0�B�\�f� ����6�\�n�ҟ���� ����>���"��� .�����ίR����Ŀ ֿ:��^�p�9ϔ�T� ��xϊ���d��� H��l��>�Pߴ�\� ������v� ������ h�(�ߞ߰�4�L��� ������@�R��v� 6���Z�l������� ��*���N��� ���� ��������X�� �J
n��� b����"4F �/|</N/�Z/� ��//�/0/�/?f/ ?�/�/e?�/�?�/�? �?�?,?�?P?b?t?�? �?DOjO|O�?�OOO (O�O�O^O_0_�O<_ �O�O�_�O�__�_�_@H_�_l_~_Go�dS�b�m�oLj�  ��rLj �a�o�Y
� �o�o�o�o{j�UD1:\|���^aR_GRP 1�n�{� 	 @�PRd{N�r����~��p����q+��O�:�?�  j�|�f������� ���ҏ����>�,� b�P���t����������	e���\cSC�B 2ohk  U�R�d�v����������Я�RlUTORIAL phk�o-��WgV_CONFIG qhm�a�o�o���<�OUTPUT� rhi}�����ܿ� ��$�6� H�Z�l�~ϐϢϴ�z� ɿ���� ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� �����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/��/ �/??0?B?T?f?x? �?�?�?�?�/�?�?O O,O>OPObOtO�O�O �O�O�?�O�O__(_ :_L_^_p_�_�_�_�_ �_f�x�ǿoo,o>o Poboto�o�o�o�o�o �o�O(:L^ p�������o  ��$�6�H�Z�l�~� ������Ə؏���  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x���� ����������,�>� P�b�t�����������������X��� #��N�_r� ������ &8J��n��� �����/"/4/ F/X/i|/�/�/�/�/ �/�/�/??0?B?T? e/x?�?�?�?�?�?�? �?OO,O>OPOa?tO �O�O�O�O�O�O�O_ _(_:_L_^_oO�_�_ �_�_�_�_�_ oo$o 6oHoZok_~o�o�o�o �o�o�o�o 2D Vgoz����� ��
��.�@�R�d� u��������Џ�� ��*�<�N�`�q��� ������̟ޟ����&�8�J�\�k��$T�X_SCREEN� 1s% �}�k�����ӯ���	���Z�� I�[�m�������,� ٿ����!�3Ϫ�W� ο{ύϟϱ�����L� ��p��/�A�S�e�w� �� ߭߿�������� ~�+��O�a�s��� �� ���D�����'� 9�K������������ ����R���v�#5G�Yk}����$U�ALRM_MSG� ?�����  �n���	:- ^Qc������� /�SEV  ��2&�EC�FG u��  n�@� � Ab!   B�n�
 /u����/ �/�/�/�/�/??%?�7?I?W7>!GRP �2vH+ 0n�	� /�?� I_B�BL_NOTE �wH*T�G�lu���w�T ~�2DEFPRO� =%� (%�O�w�	OBO-BTELEOPGO#O�O�O�O �O�O�O�O_�O&_�?��0FKEYDAT�A 1x���0p W'n��?�_�_0z_�_�_�Z,(�_o�n�(POINT� ERon  I�RECT@oko�PN�DUo�oOcCHOI�CE]�onTOUCHU`O�o�_ �o7[mT�x ������!���E��Z��/fr�h/gui/wh�itehome.pngQ�������ŏ�׏�h�pointz���/�A�S���  i�direc���������şןf�/iny��"�4�F�X�|�m�choicy�@������ͯ߯�h�touchup��@�/�A�S�e��h�arwrg����� ÿտ�n���(�:� L�^�p����Ϧϸ��� ����}��$�6�H�Z� l��ϐߢߴ������� �ߋ� �2�D�V�h�z� 	������������ �.�@�R�d�v���_� ������������� 2DVhz�� ����
�@ Rdv��)�� ��//�</N/`/ r/�/�/%/�/�/�/�/ ??&?�/J?\?n?�? �?�?3?�?�?�?�?O "O�?4OXOjO|O�O�O �OAO�O�O�O__0_ �OT_f_x_�_�_�_=_ �_�_�_oo,o>o�_�boto�o�o�o�oW���k�b�����o}�o8J$v,6�{.����� ����/��S�:� w���p�����я�ʏ ��+��O�a�H��� l�������ߟ��� '�9�Ho]�o������� ��ɯX�����#�5� G�֯k�}�������ſ T������1�C�U� �yϋϝϯ�����b� ��	��-�?�Q���u� �ߙ߽߫�����p�� �)�;�M�_��߃�� �������l���%� 7�I�[�m�������� ������z�!3E Wi������� ��П/ASe w~������ /�+/=/O/a/s/�/ /�/�/�/�/�/?�/ '?9?K?]?o?�?�?"? �?�?�?�?�?O�?5O GOYOkO}O�OO�O�O �O�O�O__�OC_U_ g_y_�_�_,_�_�_�_ �_	oo�_?oQocouo �o�o�o:o�o�o�o )�oM_q�� �6�����%��7�9�����b�t���^�������,��돞�� ��3�E�,�i�P����� ��ß��������� A�S�:�w�^������� ѯ����ܯ�+�
O� a�s��������Ϳ߿ ���'�9�ȿ]�o� �ϓϥϷ�F������� �#�5���Y�k�}ߏ� �߳���T������� 1�C���g�y���� ��P�����	��-�?� Q���u����������� ^���);M�� q������l %7I[� �����h�/ !/3/E/W/i/@��/�/ �/�/�/�/�??/? A?S?e?w??�?�?�? �?�?�?�?O+O=OOO aOsOO�O�O�O�O�O �O_�O'_9_K_]_o_ �__�_�_�_�_�_�_ �_#o5oGoYoko}o�o o�o�o�o�o�o�o 1CUgy�� ����	���?� Q�c�u�����(���Ϗ ������;�M�_��q�������~ ��}�~ ���ҟ@���Ο�*��,� [���f�������ٯ �������3��W�i� P���t���ÿ���ο ��/�A�(�e�Lω� ��z/���������� (�=�O�a�s߅ߗߩ� 8���������'�� K�]�o����4��� �������#�5���Y� k�}�������B����� ��1��Ugy ����P��	 -?�cu�� ��L��//)/ ;/M/�q/�/�/�/�/ �/Z/�/??%?7?I? �/m??�?�?�?�?�? ���?O!O3OEOWO^? {O�O�O�O�O�O�OvO __/_A_S_e_�O�_ �_�_�_�_�_r_oo +o=oOoaosoo�o�o �o�o�o�o�o'9 K]o�o���� ����#�5�G�Y� k�}������ŏ׏� �����1�C�U�g�y� �������ӟ���	� ��-�?�Q�c�u���� ����ϯ�����0����0���B�T�f�>�����t�,��˿~��ֿ� %��I�0�m��fϣ� ������������!�3� �W�>�{�bߟ߱ߘ� �߼�����?/�A�S� e�w�������� ������=�O�a�s� ����&��������� ��9K]o�� �4����# �GYk}��0 ����//1/� U/g/y/�/�/�/>/�/ �/�/	??-?�/Q?c? u?�?�?�?�?L?�?�? OO)O;O�?_OqO�O �O�O�OHO�O�O__ %_7_I_ �m__�_�_ �_�_�O�_�_o!o3o EoWo�_{o�o�o�o�o �odo�o/AS �ow������ r��+�=�O�a�� ��������͏ߏn�� �'�9�K�]�o����� ����ɟ۟�|��#� 5�G�Y�k��������� ůׯ������1�C� U�g�y��������ӿ ������-�?�Q�c�huχ�^P���^P�������������
���,��;��� _�F߃ߕ�|߹ߠ��� �������7�I�0�m� T����������� �!��E�,�i�{�Z_ ������������� /ASew�� �����+= Oas���� ��//�9/K/]/ o/�/�/"/�/�/�/�/ �/?�/5?G?Y?k?}? �?�?0?�?�?�?�?O O�?COUOgOyO�O�O ,O�O�O�O�O	__-_ �OQ_c_u_�_�_�_:_ �_�_�_oo)o�_Mo _oqo�o�o�o�o���o �o%7>o[m ����V�� �!�3�E��i�{��� ����ÏR������ /�A�S��w������� ��џ`�����+�=� O�ޟs���������ͯ ߯n���'�9�K�]� 쯁�������ɿۿj� ���#�5�G�Y�k��� �ϡϳ�������x�� �1�C�U�g��ϋߝ�@�����������`�����`����"�4�F��h�z�T�, f���^��������� )��M�_�F���j��� ����������7 [B�x�� ���o!3EW ixߍ����� ��///A/S/e/w/ /�/�/�/�/�/�/�/ ?+?=?O?a?s?�?? �?�?�?�?�?O�?'O 9OKO]OoO�OO�O�O �O�O�O�O_�O5_G_ Y_k_}_�__�_�_�_ �_�_o�_1oCoUogo yo�o�o,o�o�o�o�o 	�o?Qcu� �(������ )� M�_�q������� �ˏݏ���%�7� Ə[�m��������D� ٟ����!�3�W� i�{�������ïR�� ����/�A�Яe�w� ��������N����� �+�=�O�޿sυϗ� �ϻ���\�����'� 9�K���o߁ߓߥ߷� ����j����#�5�G� Y���}�������� f�����1�C�U�g��>�i��>������������������,��?& cu\����� ��)M4q �j�����/ �%//I/[/:�/�/ �/�/�/�/���/?!? 3?E?W?i?�/�?�?�? �?�?�?v?OO/OAO SOeO�?�O�O�O�O�O �O�O�O_+_=_O_a_ s__�_�_�_�_�_�_ �_o'o9oKo]ooo�o o�o�o�o�o�o�o�o #5GYk}� �������1� C�U�g�y�������� ӏ���	���-�?�Q� c�u�����p/��ϟ� ����;�M�_�q� ������6�˯ݯ�� �%���I�[�m���� ��2�ǿٿ����!� 3�¿W�i�{ύϟϱ� @���������/߾� S�e�w߉ߛ߭߿�N� ������+�=���a� s�����J����� ��'�9�K���o��� ��������X����� #5G��k}��г������>����� &�HZ4,F/� >/�����	/� -/?/&/c/J/�/�/�/ �/�/�/�/�/?�/;? "?_?q?X?�?|?�?�? ���?OO%O7OIOX mOO�O�O�O�O�OhO �O_!_3_E_W_�O{_ �_�_�_�_�_d_�_o o/oAoSoeo�_�o�o �o�o�o�oro+ =Oa�o���� �����'�9�K� ]�o��������ɏۏ �|��#�5�G�Y�k� }������şן��� ���1�C�U�g�y�� ������ӯ���	��? -�?�Q�c�u������� ��Ͽ���Ϧ�;� M�_�qσϕ�$Ϲ��� �����ߢ�7�I�[� m�ߑߣ�2������� ���!��E�W�i�{� ���.���������� �/���S�e�w����� ��<�������+ ��Oas���� J��'9� ]o����F����/#/5/G/�$�UI_INUSE�R  ����h!� � H/L/_MENHIST 1yh%�  �( u ��(/�SOFTPART�/GENLINK�?current�=menupage,153,1�/0�/??0?�)�/�/13�/|?�?�?�?�'E?W>71l?�?O�#O5O�+�?W5ed�it�"TELEOP�?�O�O�O:O�?�?2k?__*_<_��/>�O148,2A_�_�_�_�_���_�_�_ o o2oDo�_hozo�o�o�o�o��\a�!\o �o/ASVow �����`�� �+�=�O������� ����͏ߏn���'� 9�K�]�쏁������� ɟ۟j�|��#�5�G� Y�k���������ůׯ ��o�o�1�C�U�g� y�|�������ӿ��� ���-�?�Q�c�uχ� ϫϽ�������ߔ� )�;�M�_�q߃�ߧ� �����������7� I�[�m��� ���� ����������E�W� i�{������������� ����ASew ���<��� +�Oas�� �8���//'/ 9/�]/o/�/�/�/�/ F/�/�/�/?#?5? � 2�k?}?�?�?�?�?�/ �?�?OO1OCO�?�? yO�O�O�O�O�ObO�O 	__-_?_Q_�Ou_�_ �_�_�_�_^_p_oo )o;oMo_o�_�o�o�o �o�o�olo%7�I[F?��$UI�_PANEDAT�A 1{�����q  	��}  frh�/cgtp/fl�exdev.st�m?_width�=0&_heig�ht=10�p�pi�ce=TP&_l�ines=15&�_columns�=4�pfont=�24&_page?=whole�pm~I6)  rim�9�  �pP�b�t��� ���������Ǐ�� (�:�!�^�E�����{������ܟ�՟�I6�� �     ��J� O�a�s���������ͯ @����'�9�K��� o���h�����ɿۿ¿ ���#�5��Y�@�}���vϳ�&��Ɠs� ����)�;�Mߠ�q� 䯕ߧ߹�������V� �%��I�0�m��f� ������������!� �E�W����ύ����� ������:�~�/A Sew���� �� =$a sZ�~���� d�v�'/9/K/]/o/�/ ��/�/*�/�/�/? #?5?�/Y?@?}?�?v? �?�?�?�?�?O�?1O CO*OgONO�O�/�/ �O�O�O	__-_�OQ_ �/u_�_�_�_�_�_6_ �_o�_)ooMo_oFo �ojo�o�o�o�o�o �o%7�O�Om� ����^_�!� 3�E�W�i�{������ Ï���������A� S�:�w�^�������џ DV��+�=�O�a� ������
���ͯ߯� ��|�9� �]�o�V� ��z���ɿ���Կπ#�
�G�.�k�ޟ�}�|ϵ����������)��4ߧ�#�`�r߄� �ߨߺ�!�������� ��8��\�C���y� ������������������$UI_PO�STYPE  ���� 	� �s�B�QUI�CKMEN  �Q�`�v�D�RESTORE 1|���  ������������mASew� ,������ +=Oan�� ���//�9/ K/]/o/�/�/6/�/�/ �/�/�/�??0?�/ k?}?�?�?�?V?�?�? �?OO�?COUOgOyO �O6?@O�O�O.O�O	_ _-_?_Q_�Ou_�_�_ �_�_`_�_�_oo)o �O6oHoZo�_�o�o�o �o�o�o%7I [�o������oSCRE��?��u1sc��Wu2�3�4�U5�6�7�8���sTATM�� x����:�USER�pd��rT�p�ks����4��5��6��7�8��B�NDO_?CFG }Q������B�PDE���None���v�_INFO 2�~��)���0% �D���2�s�V����� ��͟ߟ��'�9���]�o�R���z��O�FFSET �Q�-���hs��p� ����G�>�P�}�t� ��Я��׿ο��� �C�:�L�^Ϩ���������
����av��WORK �!������.�@ߢ�u�U�FRAME  ����RTOL_�ABRT�����E�NB�ߣ�GRP �1�����Cz  A������ *�<�N�`�r��֐��U�����MSK � �)���N���%!��%z����_'EVN�����+�vׂ3�«
 h��UEV��!�td:\event_user\�Fu�C7z���jpF���n�SPs�x�sp�otweld��!C6��������!���G|'��5 kY����� >���1�U g���/��	/ ^/M/�/-/?/�/c/�/ �/�/�/$?�/H?�/:�J�W�3�����8C?�?�? �?�?�? �?O+OOOOaO<O�O �OrO�O�O�O�O_�O '_9__]_o_J_�_�_��_�$VALD_�CPC 2�« ��_�_� w��qd�R�*o_oqo��hsNbd�j�`�� �i�da{�oav�_�oo o3BoWi{�o�o �o�o��o�P A�0�e�w����� �����(�=�L� a�s�
�������ʏ�� ���$�ޟH�:�o� ��������ڟ؟��� �� �2�G�V�k�}��� ����¯ԯ����� .��R�S�yϋϚ��� �������	��*�<� Q�`�u߇ߖϨϺ��� ������&�8�M�\� q���߶���n��� ���"�4�F�[�j�� �������������� !0�B�Wf�{�� ���������, >teT���� ���/+/:L a/p�/�/./��� ��//'?6/H/?l/ ^?�?�?�/�/�/�/�/ ?#O�?D?V?kOz?�O �O�?�?�?�?�?_O 1_@ORO9_vOw_�_�_ �O�O�O_�__-o<_ N_`_uo�_�o�o�_�_ �_�_o&o;Jo\o q�o����o�o�o � �"7�FXj� ���������� !�0�E�T�f�{����� ��ßҏ����
�,� A�P�b�����x����� Ο�����(�*�O� ^�p���������R�ܯ � ��Ϳ6�K�Z�l� &ϐ��Ϸ���ؿ��� "� �2�G���h�zϏ� �ϳ���������
�� 1�@�U�d�v�]�ߛ� ���������,��<� Q�`�r�������� ������&�;J�_ n����������� ���$F[j| ������� 0E/Ti/x��/ ��/�/�/�//,/ .?P/e?t/�/�/�?�? �?�?�/??(?:?L? NOsO�?�?�O�?�O�O vO OO$O6O�OZOo_ ~O�OJ_�O�_�_�_�O�_ _F_D_V[�$V�ARS_CONF?IG ��Pxa�  F�P]S�\lCMR_GRP 2�xk' ha	`�`�  %1: S�C130EF2 �*�o�`]T�VU�P��h`�5_Pa?_�  A@%pp*`��Vn No9x CVXdv��a��N<uA�%p�q�_R���_R B���#�_Q'��H� �l�;���{�����؏ ÏՏ�e��D�/�A��z�-�����ddIA_WORK �xe�ܐ�Pf,	�	�Qxe���G�P� ���YǑRTS�YNCSET  �xi�xa-�WIN?URL ?=�`�����������ȯ�گSIONTM�OU9�]Sd� ���_CFG ��S۳�S۵�P�` FR�:\��\DATA�\� �� �MC3�LOG@� �  UD13�E�Xd�_Q' B@ ����x�e_�ſx�ɿ�VW �� n6  ���VV��l�q?  =���?�]T�<�y�Y�TRAI�N���N� 
g!p?�CȞ��TK��:�b�xk (g��� ��_���������U� C�y�g߁ߋߝ߯���\���_GE��xk7�`_P�
�P�R,ꋰRE��xe*�.`hLEX�xl`�1-e�VMPH?ASE  xec��ecRTD_F�ILTER 2�.xk �u�0�� ��0�B�T�f�x��� ��VW�������� �$6HZl_iSH�IFTMENU {1�xk
 <�\1%�������� ��=&sJ \��������'/�	LIVE�/SNA�c%v�sfliv��9/�+�� 7�U�`\"menur/w//�/��/�����]��M�O��y��5`h`Z%D4�V�_Q<��0���$WAITDINEND��a2p6OK  �i�<��r�?S�?�9TIM�����<Gw?M�?�*K�?
J�?
J�?�8RELE��:G6p3��<�r1_ACTO 9Htܑ�8_<� �ԙ��%�/:_af�BRD�IS�`�N�$X�VR��y��$oZABC�b1�S;� ,��j�I�2�B_ZmI1�@VSPT� �y��eG�
�*�/o�*!o7o��WDCSCHG ��ԛ(��P\g@m�PIPL2�S?�i��o�o�o�ZMPCF_G 1��ii�0'¯S;Ms�Si��i��p'��g��e2��  ��G�?�t��t�uI�D_/  ��p1�r1������U� ��2�.���a����~>�C4  ´ԏ �ӈ*���*�@�N� x��$�6���5��ןȌTp���o�_C_YLIND�� {� Х� ,(  *=�N�G�:�w�^����� ȟѯ� ��7����<�#�5�r� ����������޿y�_� ���8�ύ�nπ��r�ã wQ �5 �����Sǟ���(��h��X�זr�A���SPHERE 2���ҿ��"ϧ��� ���P�c�>�P�̿t� ��ߪ�����'�� �]�o�L���p�W�i�������������PZZ�F �6