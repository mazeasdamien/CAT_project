��   v��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@���&�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	>4SUSRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  wXKaIRTs1�	o`'2 L1���L2�R�	 %,��?���a1`��b�d~a����� � � ����
 ��a�o�o1CU �oz���� �c�
��.�@�R� �v���������Џ� q���*�<�N�`�� ��������̟ޟm�� �&�8�J�\�n����� ����ȯگ�{��"� 4�F�X�j����������Ŀֿ���`/TPTX������/�` sȄ��$/softpa�rt/genli�nk?help=�/md/tpmenu.dg���Ϩ� ���υ�����&�8� J���n߀ߒߤ߶��� W������"�4�F�X� ��|����������+�a�f�b�� ($p�-����T�?�x���a�a��c���c����l��c�g����a�a�a�ah��a2�h�	f����������`���a��h��_epS��h#h�F�brc Xc�B 1)h�R \ _��� RE�G VED]����wholemod�.htm�	sin�gl	doub~ trip8browsQ �����u�� �//@/���_dev.sl�/43� 1�,	t�/_ �/;/i/??/?�/S?�e?w?�?�?�?�  ��?�?OO%O7OIO0[OmOO�E @�?�O �O�O�O�O_�F�	�? �?;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omooM'�o�o�o �o�o�o+=O as������ ���?>�P�b�t��� ������Ώ���O�� ���L�^�_'_��� ����ş�����6� 1�C�U�~�y�����Ư ��ӯ�o���-�?� Q�c�u���������Ͽ ����)�;�M�_� -��ϬϾ�������� �*�<�7�`�r�A�S� �ߺ�q���i����� !�J�E�W�i���� ����������"��/� ��O�I�w��������� ������+=O as������� ,>Pbt� ��߼���// �����^/Y/k/}/�/ �/�/�/�/�/�/?6? 1?C?U?~?y?�?Y��? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__�R_d_v_ �_�_�_�_�_�_�_��o*o�_o`oro�j��$UI_TOPMENU 1K`��aR 
�d�a*Q)*d?efault5_]�*level�0 * [	 ��o�0�o'rtpio[23]�8tpst[1[x�)w9�o	�=h�58E01_l.�png��6me�nu5�y�p�13�z��z	�4���q��]���������̏ ޏ)Rr���+�=�O��a���prim=��page,1422,1h�����ş ן����1�C�U��g���|�class,5p�����ɯۯ4�����13��*��<�N�`�r���|�53������ҿ�����|�8��1�C�U�g� y����ϯ���������"Y�`�a�o/��m!�`�q�Y�w�avtyl}<Tfqmf[0nl�}	��c[164[w��59[x�qG���/��29��o�%�1�� �{��m��!����� 0�B���f�x������� ��O�����,>����2P���� �\��'9K ������������1��/$/6/H/�Z/��|�ainedi'ߑ/�/�/�/�/���config�=single&>|�wintp���/ $?6?H?Z?	�ߐ??���gl[�<��?�߲08��
A���?,OH2��DO�?cO�O�zl �� �4s�x �O�O�$��Ol�E_W_ i_{_�_�_���_�_�_ �_oo/o�_SoeowoЉo�o�o�$;�$dokub5o��13���&dual�i38���,4�o&�o9 �o�n�o�a8��� Ao����&�8�� \�n���������m�� ���
��.�@�K�d�@v���������Z{? �;�M�sc�_;���As��X�}���e�u�� 0����O_ �J�4p�^�6e�u7���� �ｿϿ���P�)� ;�M�_�qσ�ϧϹ�@���������"�1�M�_�q߃ߕߠ� �����������7� I�[�m��������������!�����6 (�]�o��������$��74������)��C�ߟT�	TPTX[20�=Aw�24#GJ���Bw1 H������8�"H����A#��[�t!v`�R��@2�K�0�11���5S:��$treevie�w3�f3��o}381,26M/_/q/ 0�/�/�/�/�/�/~/ ?%?7?I?[?m?�o/܈5�o5%���?�?�? 
?#O5OGOYOkO}O�?$�? "2�?8"2K��O�O_�O��1�?�E�8f_x_�_ �6_ڀedit�a>_P_�_ �_oˉ/���_�Co oo�o�oB�o�o��o A�o�+=O as��o���� ���(�9���Q�x� ��������ҏO��� �,�>�P�ߏt����� ����Ο]�����(� :�L�^�ퟂ������� ʯܯk� ��$�6�H� Z��l�������ƿؿ �y�� �2�D�V�h� ���Ϟϰ������ϕo �o��o@ߧE�c�u� �ߙ߽߬�����O��� �)�<�M�_�q��� W���������&�8� ��\�n���������E� ������"4��X j|����S� �0B�fx ����O��/ /,/>/P/�t/�/�/ �/�/�/]/�/??(? :?L?��߂?1ߦ?� ���?�?�?�?O$O5O GO�?SO}O�O�O�O�O �O�O�O��2_D_V_h_ z_�_�_�/�_�_�_�_ 
oo�_@oRodovo�o �o)o�o�o�o�o *�oN`r��� 7�����&�� J�\�n���������E� ڏ����"�4�ÏX� j�|�������a?s?� �?�sO_/�A�S�e� w������������� ��,�=�O�a�#_�� ����ο��=��(� :�L�^�pς�Ϧϸ� ������ ߏ�$�6�H� Z�l�~�ߐߴ����� ������2�D�V�h� z������������ 
����@�R�d�v��� ��)����������ƚԔ*defa�ult%��*level8�ٯw����? tp�st[1]�	�y��tpio[23���u����J\menu7�_l.png_&|13��5�{4�y4�u6��� //'/9/K/]/���/ �/�/�/�/�/j/�/?�#?5?G?Y?k?�"p�rim=|pag?e,74,1p?�?��?�?�?�?�"�6class,13�?�*O<ONO`OrOOB5�xO�O�O�O�O�O�# L�O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo]o�oo�o`�$UI_�USERVIEW� 1֑֑�R 
�� �o��o�o[m�o '9K] ��� ��l���#�5� �oB�T�f������ŏ ׏鏌���1�C�U� g�
���������ӟ~� ����v�?�Q�c�u� ��*�����ϯ�󯖯 �)�;�M�_�
��~� �����ݿ���%� ȿI�[�m�ϑ�4ϵ� �������Ϩ�
��.� ��i�{ߍߟ߱�T��� ������/���S�e� w���Fߨ����>� ��+�=�O���s��� ������^����� '����FX��|� �����#5 GY�}���� p���h1/C/U/ g/y//�/�/�/�/�/ �/�/?-???Q?c?/ p?�?�??�?�?�?O O�?;OMO_OqO�O&O �O�O�O�O�O�?�O_  _�OD_m__�_�_�_ X_�_�_�_o!o�_Eo Woio{o�o0h