��   �c�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����DCSS_C�PC_T 4 �$COMMEN�T $EN�ABLE  �$MODJGRP�_NUMKL\�  $UFR�M\] _VTX �M �   $�Y�Z1K $Z�2�STOP_T�YPKDSBIO�IDXKENBL_CALMD��USE_PRED�IC? �ELAY�_TIMJSPEED_CTRLKOVR_LIM? *p D� �L�0�UT�OOi��O���&S. ǰ 8J\TC �u
!���\�� jY0 � � �CHG�_SIZ�$A�P!�E�DIS"�]$!�C_+{#�s%O#J�p 	]$J d#� �&s"�"{#�)�$��'�_SEEX�PAN#N�iG�STAT/ D�FP_BASE_ $0K$4�!� .6_V7>H�73hJ- � q}�\AXS\3UP�LW�7�<���  d4r �< w?�?�?���?�?�//	7EL�EM/ T �&B.2NO�G]@%C�NHA�DF#� $/DATA)��&e0  PJ�@� 2 
&PN5 �� 1U*.n   _VSiSZHbRj0jR(�VyT(��R%S{TROBOT��X�SARo�U�V$CUR_��Rj�SETU4"	� $d P_MG�N�INP_ASSe#�PB!� `CiH �77`e�.fXc1��CONFIG_C;HK`E_PO* }d_SHRST�gM^#�/eOTHERRB�T�j_G]�R�dT�v �ku�dVALDa_7h�e�4hT1r�
0R HLHt� 0 � lt<NerRF!YhH~t�5�1� �r�W�_A$R�� DSPH/ (�G%Q�Q�Q3�?wBOX/ 8 �@F!�F!�G �r���sJTTUIRi@ � ,�F�pE}R%@2 $�po l�_Sf��uUIZN/O 0 IF(@L�p��Z_�0�_�08?wu0  @�QWy�v	*���$$C�L`  ����!���Q��Q�V�ERSION��  XK~2�IRTUAL��0�' 2 ?�Q  (������&@^���ʐ�����ϟ��������d<�9�Cz   P�8���a��������� ׯ�����.�@� R�d�f����������� �Կ	��*�<�N�`� r����ϫϺ�̿��� �߮�8�J�\�n�)� �ϧ߶��ς������ %�4�F�X�~�|ߎߣ� .����������!�0� B�T�f�x������� �������/>�P� b���v��������� �+:L^p �������  /'/9/HZl/�/ ��/����//#? 5?D/V/h/z/�/�?�/ �?�/�/�?
?O1OCO R?d?v?�?�O�?�O�? �?O	_�O-_?_NO`O rO�O�O�O�_�_�O�O o_)o;o�_\_n_�_ �_Mo�_�o�_�_�oo 7IXojo|o�o�o �o�R�o�o�3� E�Tfx����� Տ��ݏ��A�S� b�t���������џ�� ���(�=�O�^�p� ��������ʟ߯� � �$�9�K�]�l�~��� 6���Ưۿ����#� 2�G�Y�h�z������� ��Կ����
��.�C� U�g�vψϚϬϮ��� �����<�-��Q�c� r߄ߖߨߺ������� ��)�8�M�_���� ����q�������� ��4�&[m|����� �������v3 BWix���� ���/>?/ e/w/�����/� �///(/=?L/a?s? �/�/�/�/�/�?�/O ?$?9OH?]OoO�O�? �?�?ZO�O�?�OO O 2OG_VOk_}_�O�O�O �O�O�_�Oo_._Co R_goyo�o�_�_�_�_ �o�_	o*o`oQ@ u��o�o�o�o�o�o ��&8M�\q��� ��������� "�4��X�J������ಏď�����$D�CSS_CSC �25��?Q  P�;� ��Z���~�A�����w� د������ ��D�V� �z�=���a�¿��� �����߿@��d�'� ��KϬϾρ��ϥ�� ��*���N��r߄�G� ��k��ߏ��߳��&� ��J��n�1��U���y�������GR�P 2� ����	�s�^����� ����������'�� 7]H�l��� ����5 2 kV�z���� ��/
///U/@/y/ d/�/�/�/�/�/�/	? �/-??*?c?N?�?r? �?�?�?�?�?�?OO 'OMO8OqO\O�O�O�O �O�O�O_�O%__"_ [_F__�_�_n_�_�_ �_�_o�_oEo0oio��_GSTAT �2�E��<� 6�4����w�?��5�*���`�b� � 5+�E����LD&t�����D)��X`<x�e�a��4��Z�e���` q����e����$4�1�?�|��5p�����,qy���91�d�D�� y4Wݕ� u�mwUq�|qhp�P�oq��^T4� '���1�eC��E9���/Xp���c��,�a<�`�y�q
�`��`���o�o�g ��\�n��P����� ��Џ����o�����  y �N�4�F�h���|� ��̟��ԟ����� J�ďz�������¯�� ����
� �N�4�b�,� j�P�b���������� ο����8�f�h� ���گ��������߼&� ݳ��^4�3�!6p?7�4��ߴ�Ad��տ�31'.�7�C���
����C��s$�\�_�����b*�g4�U#4��ѿ��"w���i�;)�W�X�%�\��?��J��y.����O�?���D��� z��;=Okx?~�i������b��cX��[�? �T�G�ӌ����� ��Y$��C�y��?�SDڌ�]^�ѳ�2�ѹ����K.a3���ϳ1';X�p�D�zL�^�p����� �0�B��.�x���$� rϴ��߼������� 2:hNp�� ���`�(Z�4 ^8J������ ��/�� /N/4/ V/�/j/|/�/�/�/�/ ?�D?v0?z?�? f?�?�?<ߺ���r߄� �ߨߺ�����,��� &�OJ�\�n���� �?�?
O�?�_�_�?�_ �_�_�_o&o�?Po ROXo�olo~o�o�o�o �o�o: 2T ��_���_��� �0�B�8o�l��d� ���������Џ� � ��V�<�N�p���� J����̟�(��L� ^��?V_h_O O2ODO VOhOzO�O�O�O�O4� �O�O
__._@_���� ��@�2�D�:�h�z�T� fϰ���\�������� "���<�j�P�rߠ� �ߨ��߼������� N�`��l��p���� ����"��6� �>�$� 6�X���l��������� ������:<���| ��h�����t� �Ϫ���ί��� �d�:�L�^������ ����ʿܿ0B� �/�/�??�/?L? ^?��F�?��?�?�? �?�?O�?O<O"ODO rOXOjO�O�O4?�O�O .?_2___h_z_p? �O�_�O�_�_�_�_�_ "oo*oXo>oPo�oto �o�o�o�O�_J_ N`:���/�/ FXj|��� / ���l�/0/B/T/ f/x/���xj�|� r������������_ �o$�&�,�Z�@�R�t� ������د������ �(�V�П����ʟ�� ο�������Z�@� n�8�v�\�nϐϾϤ� ��������*��"�D� r�t�ϴ�濠����� �� �2�*�<��� ��*�<�N���r��� �����̏ޏ���� V�h�z���< N(:��0�~�� ������>$ FtZ|���� �l"/4/f@/j/D/ V/�/�/���/
/�/ ?�/
?,?Z?@?b?�? v?�?�?�?�?�?O/ �/PO�/<O�O�OrO�O �OH�����~���� ������8�� �2��_ V�h�z��������O_ _�O�o�o�O�o�o�o �o 2�/O\^_d �x������ ��F�,�>�`��� ��Џ܏����<� N�D��x���p����� ��ȟ��ܟ��,��$� b�H�Z�|�����V�� �د"�4��X�j�`���$DCSS_J�PC 2`��Q ( D������ʴԿaP�� ��ʿܿ1� ��$�y� Hχ�l��ϐ��ϴ�	� ����,�Q� �2߇�V� h�z��ߞ�������� ;�
�_�.�@��d�v� ���������%���I� �m�<�N��������� ��������3W& {J�n���� ���AO4� X�|����/ ��O//0/B/�/f/ �/�/�/�/?�/'?�/ ?]?,?>?P?�?t?�? �?�?�?O�?5OOO XO}OLO^O�O�O�O�O �O�O_�OC__g_6_ �_Z_l_�_�_�_�_	oP�_oʣ��S����ALouo&o�o͠ddo �o�o�o�o	�o-�o Qu<�`r� �����;��_� &���J���n�ˏ��ُ ���ڏ����m�4� ��X���|�ٟ����ğ !��E���0�y��� f�ï��篮��ү/� ��S��w�>���b��� ����������=�� a�(υ�Lϩ�p��ϔ� �ϸ�����%�K��o� 6ߓ�Z߷�~��ߢ��� ��#���1��k�2�D� V�h���������� 1���U��y�@���d� v�����������? c*�N�r� ����� q8�\�����/�%/�FdMOD�EL 2Sk�x��
 <�c� (  � �(�/�/�/�/�/�/�/ �/??d?;?M?�?q? �?�?�?�?�?O�?O NO%O7OIO[OmOO�_ �Oy/�O�O&_�O_\_ 3_E_W_�_{_�_�_�_ �_o�_�_oXo/oAo �oeowo�o�o�o�o �o�o�O�O�O/� ������� �P�'�9�K�]�o��� Ώ�����ۏ���� #�5���Y�k���Se �����������1� C���g�y�Ư������ ӯ���D��-�z�Q� c�u���������Ͽ� .�ɟ۟	�ψ��q� ���ϧϹ������<� �%�7߄�[�mߺߑ� ����������8��!� n�E�W��?�Q�cϑ� ��y�����F��/�|� S�e�w����������� ��0+=Oa ��������� >���]o� �������/ #/p/G/Y/�/}/�/�/ �/�/�/$?�/?Z?1? C?U?+�?O}?�?�? �?�?2O	OOhO?OQO cO�O�O�O�O�O�O_ �O__d_;_M_�_q_ �_�_�_�_�_�?*o�? �_oroIo[o�oo�o �o�o�o�o&�o\ 3EWi{��� ������/�A� o��;oi�{�菿�я �����+�=�O��� s���ҟ����͟ߟ� �P�'�9���]�o��� �����������߯� ^�5�G���k�}���ܿ ��ſ����H��1� Cϐ�g�y��ϝϯ��� ������D��-��� '�U�g���O߽����� ���R�)�;��_�q� ����������<� �%�7�I�[�m����� �����ߝ�����J�� 3EWi{��� ����/| Se������ �0///f/A/ S/�/;/�/�/?�/�/ >??'?t?K?]?o?�? �?�?�?�?�?(O�?O #OpOGOYO�O}O�O�O w/�/�/�O�O�O_1_ ~_U_g_�_�_�_�_�_ �_�_2o	ooho?oQo couo�o�o�o�o�o �o�Ov_?Q '�����*�� �%�7�I�[������ ޏ��Ǐُ����\��3�E���i�{�������$DCSS_PS�TAT �����Q �   �� � (&�K�2�o���� ������ $�˟į֯������ �����'��SET�UP 	�B	ȶ�����X�r�� ��������ۿ��g��T1SC 2
K�����Cz��#�5�|G� �CP R�D$�Dl�Ϥ�^ �����ϻ��"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��� ��~������- �Qcu���� ���//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�__ /_BS_e_w_F_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o'9K] o������� ��#�5�G�Y�k�}� ������ŏ׏���� �1� _U�g�y��_�� ���������	��-� ?�Q�c�u��������� ϯ����)�;�M� _�q���������˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �!�3�E�W�i�{�J� �߱�ğ��������� /�A�S�e�w���� ����������+�=� O�a�s����������� ����'9K] o������� �#5GYk} ��������� /1/C//g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ �!o3oEoX/io{o�o \o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�ok�}� �o^���ů������ �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m���ڨ�$DCSS�_TCPMAP � ������Q @ *���⠽�U����U	�
������W�  U����U���⡪�������� �!��"�#�$�%��&�'�(�)��*�+�,�-��.�/�0�1��2�3�4�5��6�7�8�9��:�;�<�=��>�?�@��U�IRO 2����������� 0BTfx�� �����,���U��y�� �����	//-/ ?/Q/c/u/�/�/�/6 �/Z�/??)?;?M? _?q?�?�?�?�?�?�? �?OO%O7O�/[O�/ O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_��_�_�_NO�_��UI�ZN 2��	 �����(o:oLoR� %ozo�o�oao�o�o�o �o
.�oRdv E������� �*�<�N�`�#����� e���̏ޏ�����&� 8��\�n���C����� ȟ������ӟ4�F� X�'�|�����c�u�֯�请���0��_��U�FRM R�������w��������� ѿ�����+�=�O� a�sυϗϩϻ����� ����'�9�K�\�r��\߄ߖ�qߺ��� �������&�8��\� n�I��������� �����4�F�]�o�|� ��-������������� 0TfA�� w����� >Pg�t�%�� ����/(//L/ ^/9/o/�/�/�/�/�/ �/ ??�/6?H?_l? ~??�?�?�?�?�?�? �? O2OOVOhOCO�O �OyO�O�O�O�O
_�O ._@_W?d_v__�_�_ �_�_�_�_�_o*oo No`o;o�o�oqo�o�o �o�o�o&8O_! n������ ��"��F�X�3�|� ��i���ď�����Տ �0�B�Yf�x���� ����ҟ䟿����� >�P�+�t���a����� ί����߯(�:�Q�