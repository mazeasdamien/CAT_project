��   >��A��*SYST�EM*��V9.4�0107 7/�23/2021 A 	  ������CCHG_�LIM_T  � �
$COM�MENT �$CTRL_STATE  M�IO_TYPX
I�DXXUFRAM�E_NUMxTO�OL�INSID~WMARGINX �$UPP_XY�Z4   �$LOW��/C�FG8� a�$KNOB_MO�UGZ �SE�L�EF�GRIP_wENBOPE� {)CLOSW �)LEVER�L�V_DIR_PY�XBTN_OUT�YeYuONE�_HANDXAV�G_F�� ROT�_^TRNS� T�R �b�uSFD�OD�  �$ORG_PTH�_RES�TOUCH�OC�*��$JNT4MR�G�3$,$�G+C"2a3�U"l(�SP�8u#�)�WPR�*�)�DC���#$R�EC_METHO��'b �$e�$uT�EACH_PAT>#MULTI7�!|�&CUSTO��GEN_TP_PRO= )T�*�� �e=�� ]1DEV��5���_AR� 3  
�K9_2 �K_S0�n�1ENC�SB~�2,$�0_RIGH��/!HDL_MAS�BCV1�A�2�VA�5EG�5E+L=JML+G�1F_�1 �7�FF_VAL�ID_M�MAX�_RUN� + � GAIN��G� �3!�� J(k!�F� SNG�L�R;"��B� P���X�22T�!�0_AR�3�!�PT]1C��CUR_F5PTS�M�@wX�APUSH_F�C�@�Y�U�T�Uħ3;T3S��'$�!�YJ1_R�V�@�j5�[SIMPLE-QXOF�F<a�E3SH� M1OK�^�.RO�RSV Nt� �2sbREA@ܻ�cSTR|a?>�0DEBUG� ���DATA8$ S�6�@ ^�@ �esP�oT�lb.*� rQ3!wrl lc�02�S PRSW�NE��REBO�2�I�T�]dNON_R�ST�FSA/bITgnsORCW ."�r��C."MEAN�zH�DGD_ACTI�VWSAFEM1
��tO�u�r�@�$0�`�X�P PS�T�bNEqp�4 �S�S�xf�S_W�P."EX�{ -�h�,$��@�`�V] ��3!�!��l ���T�� d��d��-���X����SMAL�A���@OCVR���+��FO=���@l H�1G�U�5�G�BE���vAF���wESCAPE��TOP�f$CL�AL�aAlTDDS1BrQ�!TCg � �e�%rQ�)rS�Wꕿ)  Yu�"*z�w���������rQ.XM3?V?uE�gSUBS0GtN�O_M�Ė�DBp=!ߦȦ�WAIXt��jP�A��b�'8�NiT`r�qbT_ϓ:Y�C�DOW3Sm�1N�v�3�FC���1�B�e�1T @�gtfV���jV�2/ MQ0� 6T��P�9Vmd ]l`@0yA`�.���!T�dTL_OR84 �E�AMOMW�2����GRV_OF C2���!�2��`F�ÇRSL��LQu!�F!I�q�$ud��f�����GRP>8 � A
T4� qp��IIO�RL8��1DI��3AP�W�3�5VE IT4SjVR@0MD�'��jІݠQ2v}�:�/ S�\ 9$PAUS������G�ABWҔDAP�5 	Uoq���P�W� WM��@:�FIb��T�U���ERR�f�u�Bd�W���RETRY %�,Q���������(T`HtC�AqpR�A��O�1�3�BՔ�1᠀��]�bC��W�\Tpbp�u�rL�O�b����LOO L���"2����+՘��ɛ�EN�5d���E���]�UaE U� RT�Ǖ3�ONL�SP� OFFG�BLIN�1caĖ`(�� 7B K�7UaALAR���Q�)� q��Ua��zҦk�)'�b8�rn�Ǎd9 �ԻeP���W�m�ӑ�lu�O*�ID1`H��h��OOPERn��I����P�C�_�	$GWIR`p��sPCY���� ��m�CHA�R���VOLTAd(�C҉RI*�IO�;�O�a�Lr0�`0ӑ�lCONNcEC��6OT�` �����Ґ���A�&NE;��3꒼a� U"�&��♛��6.�PcSW����$3PA���T�)6A1776�aIN�p!Z4�0�d4 a7 m3da*3!��PATHҭ�o!"~b�cTt�`�8 �b3�;�:3���3sPH!H�I> �,a@�zʼ2V��ÚaDa1Q\Gm1jH3gK4gK�5gA��$̑SS�������A��Y��� Y�@�PSIO�N�H��XK�AIRTU�`�O�@ܶb�� �HY��AY)�A._@_'_d_XF[��|_B�FV�Vq�P�_�U �_�FU@����PF< �_<�R��Po�S>aCH  A�P2a1@�_Em�R)
��!�G_01�_n�Q�A�?��T
 P1 o�S�]B/`/��E;� �e�a� �`�e�o�o�o�o�o  $6HZl~� ����9��� � 2�D�V�h�z������� ԏ���
��.�@��R�d�FZ�PBΔT�P��T�ӟ�?��3�@ ��  ��X�P�Q���UA����`�����"��3a�Q��+�*�^�`=���*�B+�_=L��?ϕp�P�� B�Q��.bx��������R u0  sЊ���  d:a�>�aw�?��<#�
&�7d�b�U�І���2�_9�K�]�o����� ����ɿۿ"����#� 5�G�Y�k�}Ϗϡ�FX
 W_FR���� ���
��.�W�R�d��vߟ߿A T�!  Y�a����������� ���_�[.�_͖b����FZ������ �&���/�\�S�e��� ������������" f�$��HO�w� ��������) M�q���� ���//ZlI/ [/m//�/�/�/�/�/\�/��MTPS\�'ҡ�-����5?�T*??�?�?���n?�?�?�?�/GRP� 3[2 l��� 	MfnG@T9P��kl0?��P:`\��4!  UFXd�� 3OEI�AUM�GoO�O�O�Ogc3�O(X�O�O�O_gc4*_�XG_Y_k_}_gc5�_ h�_�_�_�_KC6olho1oCoUoKC7no�h�o�o�o�oKC8�oDx�o	-KC9F�xcu��KB1ѠTM��� ���QO��;�M�_� q���O󉧏��ˏݏ �)__��%�7�I�� �_˙��������o 7�����!��mo�� W�i�{�����o�ï կ����E{�/�A� S�e���繛�����ѿKB2�S���+� =�OÉ���sυϗϩ� O���+�������O� a���K�]�o߁�O�͟ ��������O�9�o� #�5�G�Y�Oå���� �����O��G���� �1�O�}���g�y��� ��O��	������	KB3Uϋ	?Qcu ����	����� -�c);M��� �������;) �//%/�q�)[/ m//�/�#��9�/�/ �/�/�#I�93?E?W? i?�#���9�?�?�?�? �#!WIOO/OAO�"4��IwO�O�O�O�C �/Y�O�O__�Ce �YO_a_s_�_�C�i �_�_�_�_�C=/si'o 9oKo]o�C�/�i�o�o �o�o�C?Ky�o# 5�C�?�yk}�� �C�?#������C�YO��C�U�g�y��"5��O������Ӊ�$C�CSHG_CFG ���Y��Y����3����ӄ
֖������Bb����ֆ�ӈ�ցř����ؖɝ� ���<�i�{��X�����ѯ�������+�G���A �Y�0��	12�345679����90������Ϳ�߿���|��  !��2�*�*�<� N�`�rτϖϨϺ�������
��.�@� R�d�.���꯿�������ߴ��+�=�� �ϴ�Z�l�~����