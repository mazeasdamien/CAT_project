��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$VOERSI� � �0�COUPLE]  o	 $�!PP�1CES0�2eG ��PB> �1
 � �$SOFT�T�_ID�2TOTA/L_EQ 0�1�@qN" �@U SPI
 ��0^�EX�3CREt -DdBSIGJ@�dOvK�@PK_�FI90	$T�HKY"WPANE��D � DUMM�Y1dIT1TU4�QQ!Rx1R� � $TIT91� ��� �Td�T0��ThP�T5�V6�V7*�V8�V9�W0�W�W@OQ�U�WgQ�U�W1�WU1�W1�W1�W2�R~OASBN_CF�![@$<!J� �; ;2�1_CMNT��$FLAGS�]�CHEK"$�b_OPTJB6 � �ELLSETUP�  `@HO,8@9 PR�1%�c#��aREPR�hu0D�+�@��b{uHM�9 MN�B;1 U�TOBJ U��0 49DEV�IC�STI/@� � �@b3�4pB�d�"�VAL�#ISP_�UNI�tp_DOxcv7�yFR_F�@�|%u13��A0s�C�_WA�t,q�zOF�F_T@N�DEL��Lw0dq�1�Vrc?^q�#S?�o`�Q"U�t#*�QTB����MO� �E' � [M������REV�BI�L���XI� v�R_  !D�`~��$NOc`AM�|���ɂ/#@ǆ� ԅ���1X�@}Ded p E �RD_E��h�$�FSSB6�`KBoD_SE�uAG� G�2Q"_��2b�� V!�k5p`(��CO@�0q_ED� � G� t2�$!S�p&-D%$� �#�B9�ʀ_OK1��0] P_C� ʑ0t���U �`LACI�!��a�Y�� �qCOM9M� # $D
� ���@���J_\R���BIGALLOW�� (Ku2-B�@VAR���!�AB B_�BL�@� �� ,K�q���`S�p�@M_O]˥���CCFS_U	T��0 "�A�Cp'���+pXG��b�0 =4� IMCM ��#�S�p�9���i �_D�"tk���M�1� h$�IMPEE_F�s��s��0� t����D_���J��D��F�� �q_����0 T@L��L�DI�s@G�^� �P��$I�'����CFed X@G�RU@��Mb�NF�LI�\Ì@UIR�E�i42� SWIYTn$`0_N�`S 2�CF�0M� 	�#u�D��!��v`(����`J�tV��[ �E��.p�`�ʗELBOF� �շ �p`0���3����� F�2T��A`�rq1�J1��z _To!@��p��g���G�� �r0WARNM�p#tC�v`�ç` �� COR-UrF�LTR��TRAT�9 T%p� $AC�CVq��� ��r$�ORI�_&�RTr��S<�m�CHG�0I���TW��A�I'�T��!D��� �202�a1���HDR�2��2�2JP; S���3��4��U5��6��7��8���9 1��׀
 �2� @� TRQ�$�vf��'�1�<�_U�<�G��Oec  <� P�b�t�53>B_�LLEC��!~�MULTI�4�"u�Q|;2�CHILD���;1ذO�@T� "'�STY92	r��=��)2���ױ��ec# |r056$J ђ��`���u�TO���E^	EX�Tt����2��2�2"�0����$`@`D	�`&��p������ %�"��`%�a�k�����s�����& '�E�Au��Mw�9 n�% ��TR�� ' L@U#�9 ���At�$JO�B����PM�}IG��( dp���� ��^'#j�~�x�p{OR�) t$�3FL�
RNG%Q@�TBAΰ �v&r�* `1t(��0 �x!�0�+�P�p�%Q!��*��͐U��q�!�;2MJ�_R��>�C<QJ�8&<J D`5CF9���x"�@?���P_p�7p+ \�@RO"pF�0��I9T�s�0NOM��>Ҡ�4s�2�� @U<PPTgў�P8,|Pn�ć0�P�9�͗ RA����l�?C�� �
$�TͰtMD3�0TD��pU�`�΀+AYHlr>�T1�JE�1 \�J���PQ��\Q��hQ�CYNT�P��PD'BGD̰�0-���PU6$$Po�|�u��AX����TAI�sBUF,���A�1�. ����F�`PIV|�-@PvWMuX�M�Y�@�VFvWSI�MQSTO�q$7KEE�SPA��  �?B�B>C�BذP��/z�`��MARG��u2�FACq�>�SLEW*1!0����h
�N�s�CW$0'����pJB�Ї�qD�ECj�eG�?�dbV%1 Ħ�C�HNR�MPs�$G_@�gD�_�@s���1_FP�5�@TC �fFӓC�Й���qC���+�VK�*��"*�JR|x���SEGFR$`�IOh!�0STN�L3IN>�csPVZ�cb�A�D2����r 2���hr�rz�P��3` +^?���եq�` ��q|`�����t��|aSIZ#�!� ��T�_@%�I��qRS �*s��2y{�Ip{��pTpLF�@�`��C3RC����CCTѲ��Ipڈ�a���b��MI�N��a1순���D
<iC �C/���!uc�0OP4�n j�EVj���UF��_!uF��N�����|a��=h?KNL�A�C2�AVSC�A�@A�� ��1��4�  cSF0�$�;�Ir �4�@�05��	D-Oo %g��,,m����ޟ���BRC�6� �n���sυ�U��Rޝ0HANC��$L�G��ɑDQ$t�NYDɖ��AR۰N��`aqg��ѫ�X�ME��0^�Y�[PS�RAg�X�CAZ�П���rEOB�FCT��A��`�2t!�Sh`0ADI��O ��y�s"y�n!����Ј��~#C�G3t!��BMPmt@�Y�3�af�AES$�����W_�;�BAS#XYZ'WPR��*�m!���	 ��U�87 � ƀI@d���8�\�p_C:T���#�abR_L
 � 9 %���C�/�(zJ�KLB�$�3�D�<�5�FORC�b�w_AV;�MOM*�q�SaԫBP`Ր�yӐHBP�ɀE�F����A�YLOAD&$EAR�t&3�2�Xrp��!� �FD�� : T`I�Y3���E�&��Ct��MS�PU
$(kpD�&�9 �b�;�B�	7EVId�
�!�_IDX   $���B@X�X<&v�SY5� ���_HOPe�<��AL�ARM��2W�rY�R9_�0= hb P�nq�`M\qJ@$PiL`A&�M#�$�` ��� 8�	���V�]�0�U��U�PM{�U���>�TITu�b
%�![q�BZ_;�.��? �B pQk���6NO_HEADE^az��}ѯ��`� �����dF�ق�t�P����@�@��uCIGRTR�`��ڈL���D�CB@4�RJ�� 1�[Q���A�2>�&��OR�r��O����F`UN_OO�Ҁ�$����T������I�VaCnpb`DBP�XWOY���B�P�$SKADR��DB]T�TRL��C���րfpbDs��~�DIJj4 _�DQ}���PL�qwbWA���WcD�A��A�=�2�UMMY�9��10�a�D�B����D;[QPR~�� 
��DМZ���E O�Y1�$�a$8���L)F!/����0G�G/���PC�1H�f/���PENE�A@Tf�I�/�$�C�OR`"JH �@ �E$L�#F$#PR���+jp��nq��_D$�qPROSS]�
���R�r�` u�$TRIG96P�AUS73ltETU�RN72�MR:�U2 0Ł0EW$��`?SIGNALA�QR�$LA�З5�1G{$PD�H$Pİ"�AI�0�A�C�4�C��DO�D�2�!��6GO_AWAY�2MOZq�Z�W D{CS��CSCBg��K Իa#���ERI�0Nn�T�`$������FCBPL�@QBGAGE���P��ED|B0D�wA[CD�OF�q[F�0�FoC��MPMA�B0XoC�$FRC�IN��2Dk��@���$NE�@�FDL|8�� L� ��@��=��Rw�_��P� OVR10���l�~��$ESC_�`>uDSBIO����pTe�E�VIB�� �`s��Z��V��pScSW��$�VL��:�Lk��X���ѣ�bQ�����USC�P��A8=�	Q�MP1%e&S�*`�(bt`'c5۳ESUd��-cWg&SWg ?cWd����Wd��Wd.���AUTO$�Ya҃�ac�SB����-d���&SwB[��GB�f$/VOLT�g ��  �GAOD!�qr���@:�ORQҀ�Kra�$DH_THE&0�Rgp� qtnwALPHnt��o���w0 Vp]�$�.�R a�[��s�5�`r�CQ#RBUD�S� F1M�B�sV
��;��Lb��tk���BRTHR���L��T`�Z���Vɖ��DE  �1��2�⋅�� ������kѯ�aәT t0V�ꆸ������̈ Я�-�"�N~��sxS2����INHB��ILTG0ɡ�T?��3 $�w��E��PqQxQ�ThqPe��0Y�AF}�O�ນ��ڗ�� qPڳē����bPܙ����PL?���3���TMOU��ēS���� ���s�/�S18���O�A�ܙ��I����CDI8Ƒ˩o�STI��գ��O:ҋ�,0���AN��Qg�S��+r��#x$�����w�_�����PRA�P`pvC����MCNeQ�e�����VERSP��r�oPIw�FP�åǲШ۷G.�DN"��G>�����F�2ŤǷ�M�7�F��_
�MN�D̠,����d �{ƭa����OB��`�U˱z���DI�� ��#���3�����A����w�Fx���3�ONp�5��Q��VAL�{CR[�_SIZ��8b�;Qn�REQ�Rb�`�]2b���CHq� ΂�ڃ�Ռ�����:��n�S_U��X��wWF�LG���wU$�CV�iMGP�QδFLXP�923R�u���&EAL�P-�C	�F
+rT��W��� �R�cx���NDMS7�d ��K>S�P_M'0h�STWv�������AL�P���Q���pU���U�IAG,��o��d�U�-�T"A-`� ���A������H`��Q`��6��Pq_D&��1s��.�P��F�>2�T�� ?7 1A>��#�t#L��?_0=i @@>LD�c�F�0�FRI�0 �`Ѐ��1}ѲI�V\1�*�^1�UP�`��a��C�LW��
`L=S&-c&&S�C.w�� L����!����d�Q$w�҇��$w���8�
�P�5RSM��(�V0h � r��d6^2AW�a_TRp}��8@NS_PEA�����< ��$�SAV�G�8�6G]%���CAR �`�!�$���"�CRa���$ d�#E8�@��"STD���!qFpo��'QOF���%��"RC���&RC۠�(F�2A�R#7��X�%, gMA�Q_�a���
QQ��al2��u4Ib�r7I�R�9wQH�7�8M/��!Cp�R�  �p�2F�<�SDN�a0 ���W2QM P $Mi��s$cA� $C�cm�9���4�A�T�0CY_ wN LS!IG1x'�yB��y@@H2Y�N�O����SDEV�I�@ O@$n�RBT:VSP�3�CuT�DBY|�A	W|`3CHNDGDAwP H@GRP�H	E iXL�U��VS�F�x2� DL1p Q06ROp��FB�\]�FEN�@��S��C�hAR d�@DO<d�PMCSb�P�薇P�R��HOTS�Wz42�DMpELE��1/ex\8`�RS T��@���r� hf��`OL�GHA�Fk�Fs���|�C�A@T �� $MDLUb 2S@�E���q�6@�q	0�i�c�e�cJ��	uݢ�#~5t+w�PTO��� �b��e�SLAVS� U;  ��INP �	V��ЊyA_;�ENU�AV $R�PC_�q�2 1bL�wpp�b�pSHO+� WA ���A�a�q�2�r��v�u�vcB_CF�� X` ,f��r�OG gE��%XD�h�{PC�Iߣ�i�MA��D�x AYr?�W� p�NTV	��D�VE�0@�SKIB��T�`g?Ň2��" JZs�! Cꆻ���f�_SV/ �`X�CLU��H���O�NL��'�Y�T��O=T:eHI_V,11 �APPLY��HI�4`;�U�_ML�� $VRFY8��	�U�M{IOC_�I���J 1/��߃O��@X�LSw"`@$?DUMMY4����ڑ�Cd L_TP����kC��^1CNF f���E��@T�y� 	D_#UQ_��ݥ�YPCP��=�� �������uJ �� Ys +�
0RT_;P���uNOCCb 3Z�r�TE����=�פ DG�@[ �D�P_BAe`3kc�!��	_��H��u��� \�pAb=cA7RGI�!$���`�[ �tSGN�A] ��`U��I�GN�Տ��� ���V������ANNUN��&�˳�EU�J'�ATCH��J���pt�rA^ <`@g�����:c$Va��������AE�F] I�� _ �@@FͲITb�	$TOTi �C�O��c�c@EM�@NIF�a`tB��c��ùA>���DAY@CLOAD�D\�n���� ��EF7�X�I�Ra��K���O�%��a�ADJ_)R�!@b��>�H2��"[�
 c�%��`a�͠MPI�J��DR�qA��?�Ac 0� �х�� ��Z�ϡ��Ui ��CTRLܖ Yp d��TR�A8 ?3IDLE_�PW  �Ѡ��Q��V��GV_���`c ��o�;Q@e� �1$��6`<cTAC�-3��P�LQ�Z�Rdz\ A-u:ɰSW;�A\���/Jղ�`b�K�OH�(OsPP; �#IRO� ��"BRK��#AB  �O������� _ ���F���`d͠, j@�S�RQDW��MS��P6X�'z��IF�ECAL�� 10^tN��V��豊�V�(0��CP
��Nr� Yb�0FLA_#f�OVL ��HE��>�"SUPPO��ޑ�\�L�p��&2XT�$Y-
Z-
W-
���/��0GR�XZl�q�$Y2�CO�PJ�SA�X2R��*r�!���:��"~RI�0)��f `�@CACH�E��c��0�s0L}AZ SUFFI, C��{Q\��哹6�%�MSW�g� 8�KEYIM[AG#TM�@S���n
2j�r��r�OC�VIE��~�h ��aBGL����`�?��@���0�i��6!`STπ!�����������EMAI�`N��`Ac@NZ�FAU� �j�$"{Qa��U�3"��u E}�k< �$I#�US�� �IT'�BUF`�r�DNB���SUBu$��DC_���J"��"SAV�%�"k�������';��P�$�UOR	D��UP_u �%��8OTT��_B`��8@�LMl�F4��C7AX�@Cv���Xu 	��#_uG��
�@YN_��R�l6���D�E��UM����T��F���caC�DI`BED%T)@C��~�m�rI��G�!c�&��l`����A�P��FZP n (�pSV� )d\��ρ���A��o�� ����>"$3C_R�IK��kB���hD{pRfgE.(AD�SP~KBP�`�II�M�#�C�Aa�A��UЂG���iCM! IP`��KC��� �DTH� ȷS�B*�T��CHS�3�CBSC��� ���V�dYVSP�#[T_D^rcCONV�Grc�[T� �Fu F�ቐd0�C�0j1��SC5�e�]CMER;dAFBgCMP;c@ETBc� p\FU D�Ui ��+�~�C�D�I%P702# �E	O���qWӏ�SQ��1QǀSU��MSS�1j�u�4`�Tr�Aa��A>�1r� "�Й��4$ZO@s���"l�U6�&��eP���e�CNc�l��l�l�iGGROU�W)��S c�MN�kNu�eNu�e NpR|b|�i�cH�pi�8�z
 �0CYC���s`�w�c��zDEL�3_D��RO�a�� �qVf���v{�O�2� ��1��t��:R�ua�.#�� ��AL� �1s@ˢI1¡�J0�PB�� A4?`R^�T�Gbt ,!@��5膁aGI1LcR1s �
PC������1u ���������P����EC�	������2���J0�0vH *	�LU�1#J�Q��V
� [�7Az���z��z�Ѡz��z�Fz�7w�8Bw�9w���y���1��U1��1��1��1ĚU1њ1ޚ1�2���2����2��2��2���2Ě2њ2ޚ2*�3��3��3����U3��3��3Ě3њ�3ޚ3�4��GBX	TF��1w6�.(�0�f��0�U�0ŷ�e%�FD�R5�xTU V�E��?1���SR��R�E�F���OVM�~C)�A2�TROVf2�DT� R�MXa��IN2���Q�2�IN	Dp�r�
���0�0�0�Gu1��[�G`��{�D_�[�RIV�P��oGEAR~AIOr�	K"N�0�y�p��5`@�a�Z_MCaM� �����UR�R�yǀ��!? ���p?nЋ�?En�ER�v�3���!��P��zE@:�PXq�B�RI0% �#ET�UP2_ { ����#TDPR�%T�Bp������E!�"BAC�2| T��"�4E)�:%	`^B��p�WIFI��� Mc����.�PT��DMA��FLUI�}c � ��K UR�c!���B�1SPx E�ESMP�p�2$��S^�?x��Jق0
3�VRT���0x$S�HO��Lq�6 AS�ScP=1��PӴBG_�����<�FORC��g㶙d~)"FUY�1��2\�2
Eh� p�� |��NAV�a)�������S!"��?$VISI��#�SCM4SE����:0jE�V�O��$��X�M���$��I���@�FMR2>��� �5` �r�@�� �2�PI�9 F�"�_���?LIMIT_1�d�C_LM������D�GCLF����DY&�LD����5���Ϥ���M�Fc���~u	 T�FS0Ed� P��QC�0$EX_QhQ�1i0�P�aQ3�5��GoQ��� �l���RSW�%ON�PX�EBUG��'��GRBp�@U�SBKv)qO1L� ��POY 
)��P��eM��OXta`SM���E�"�ю��`_E �� �0F���T�ERMZ%�c%Dp�'ORI�1_ �c%�KSMepO��_ �c%OXK��`�(�c%���UP>� �g� -���b����q#� ���G�*� E�LTO��p�0�PFIrc�1Y��P�$�$߆$UFR��$��1L0e� OT�Y7�PT4q�k3NS]T�pPAT�q4OPTHJ�a`EG`8*C�p1ART� !5p� y2$2REL�:)ASHFTR1�1��8_��R�Pc�& � $�'@�� ��H�s�1 @I�0�U�R} G�PAYLO�@�qDYN_k���.bp�1|��'PERV�� RA��H��g7�p�2�0J�E-�J�RC����ASYMFLTR��1WJ*7����E �ӱ1�I��aUT�p bA�5�F�5P�PlC��Q1FOR�pM�I!���W��/&��0F0�a.H��Ed�� �m2N���5`OC�1!?�$OaP����c���,��bRE�PR.3�1Xa�F��3e��R�5�e�X�1(�e$PWaR��_���@R_�S0�4��et$3UD��NܟQ72 ���$�H'�!�`ADDR
�fHL!G�2�a�a�ar��R��U�� H��SSC����e-��e���e��SEE���HSCD��� )$���P_�_ B�!rP������HT�TP_��HU�� (�OBJ��b(�[$�fLEx3Us>�� � ����J��_��T?#�rS�P���z�KRN�LgHIT܇5��P���P�r��`�����PL��PSS<��ҴJQUERY_�FLA 1�qB_W�EBSOC���HQW�1U���`6P�INCPU���O h��q����d���d������IHMI_{ED� T �R�H�?$��FAV�� d�Ł �IOL]N
� 8��R��@$SLiR$�INPUT_(i$
`��P�� ؁wSLA� ����5�1��C��B�a{IO6pF_AS7��$L%�}w%�A��\b.1�����T@HYķ�������h�UOP4� ` y�ґ�f�¤�������`PCC
`����#�|��aIP_ME��n��� Xy�IP�`<�U�_NET�9����Rĳs�ѱ�D�SP(�Op=��BGȞp��M�A��� �l�:CTAjB�pAF TI�-U��Y ޥ��0PSݦBUY IDI�rF ��P�s񘬢 �y0�,�����Ҥ�NQ�Y R���IRCA�i� ך ěy0�CY�`EA�����񘼀�CC����R�0�A�7Q�DAY_���NTVA����$��5 ����SCAd@��CL����� p���𵁛`8�Y��2e�o�N_�PACP�q��ⱶ��,� N����
�xr���:p<�N� 2��Ы��(ᵁ����xr۠L�ABy1��Y ��UN�IR��Ë ITY�듭��e�R#�5�|��R_URL��o�$AL0 EN�Шҭ� ;�T��T_}U��ABKY_z���2DISԐ�AT��Jg����P�$���E��g�R��З �A�/���J����F�Ls��7 Ȁ���
��UJR� ��pF{0G��E7���J7 O R$J8I�7��R�d��7��E�8{�H�AP�HIQS��D�eJ7J8B��L�_KE*�  ��K��LM[� 7� <X�XRl�u����WATCH_V�A�Qo@D�tvFIE�Lc��cySp��4�� � o1Vx@��-�C�T[�9�m�����LGH��� �$��LG_SIZ��t�z�2y�p�y�FD��Ix���+!��w� \ ����v��S���2 ��p�������\ ���A4�0_gCM]3NzU
RFQ\vv�rd(u�"B��2�p����I ��+ �\ ��v�R� _�0  �Z�IPDUƣ�qLN=��ސ�p�z@6���f�>sD�PLMnCDAUiEAFp0���TuGH�Rp��|�BOO�a�g� C��I�IT+����`��RE���ScCR� �s��DI���SF0�`RGIO"$D�����T("�t|�	S�s{�W$|�X���JGM^'MNCHL;�|�FN��a&K�'�uЅ)UF�(1@�(F�WD�(HL�)STP�*V�(%Г(��(�RS9HIP�+��C�[T�# R��&p:'^9U =q�$9'�H%C𜓚"Gw)�0PO�7�*�`�#W}$���)EX��TUI�%I���Ï����rCO#C� *�$S��	)��B@v�NOFANA|��Q
�AI|�t:��EDCS��c�C�c�BO�HO�GS���B�H9S�H(IGN�����!O���DDEV6<7LL����-�ҭЦ(�;�T�$@��2�p������#A���(�`�{�Y��PWOS1�U2�U3�Qp	��2�@�Ш ��{�PtD����&q`)��0�d��VSTӐ�R�YU�B@ ` /�$E.fC.k�p�<p=fPf���4�ѩ LRТ� ��x�c�p���<�Fp�dSp?"�_ �����Kq&ü��c��MC7�� ��pCLDP|Ӑ��TRQLI#���ytFL��,r��5s8�D�5wS�LD85ut5uORG��91�HrCRESERV ���t���t���c�?� � 	u95�t5u��PTp��	�xq�t�vRCLMC�������q̐�M��k������$�DEBUGMASP��ް��?U8$T@���Ee�g��M�FRQՔ� �� j�HRS_R%U7��a��A��k5�FREQ� �$</@x�OVER���n��V#�P�!EFI�%�a��g�ǒ����t� \R�ԁd�s$U�P��?�p��PS�P��	߃C ��͢a��U\�l��?( 	R�I;SC� d@�QkRQ��	��TB �� Ȗ0A՘AX����ؗ�EXCE�Sj�oQ��M��\���;�����	᫒SC>�P � H��̔�_��Ƙǰ]����MKHԳK�J� �m�B_K�FLIC��dB�QUIREG3MO��O˫3���ML�`MGմ @�`��T���a#NDU�]��>���k�G�Df��INAsUT���RSM>�a��@N�r]3-��p�5�PSTL\�� �4X�LOC�VRI�%��UEXɶANGtuBu�S�ODA�����������MFO����Y�b@�e84�2k�SUP�eQ��FX��IGG� � ��p�c�� �cQ6�dD�%�b|�!` ��!`��|��3w�ZWa�CTI��p;� M��n[�� t��MD��I�)֟@���qHݰM��DIA�����W,!�wQ�1�D�)��O���]��� 0�CU��VPP��pu��O!_V��ѻ ���S�X�&5������P��04N���P��KES2����-$B� ����N�D2����2_T=X�dXTRA�C?��/��M�|q�`��Pv��XҰ�Pt SyBq`�USWCS���T��	���PULS,��A�NSޔ��R��JOIN��H��~`j�=��b��b�����P=��$��b$���TA����S���S�4HS�E��SCF���J��R��PLQ� 7��LO���1�.���^����8ᾊ�����0�RR2>��� 1��e�A�q d$��I$ΐ+�G�A2+/�� �PRIN܍<$R SWq0"�a/�ABCȇD_J%�¡u��_�J3�
�1SPHܠe�u�P��3�(�р`u��J/����r�qO8QIF��CSKP"z{�{�	J���QL2LBҰ_AZ�r�~�ELQ��OCMaPೕ�T���RT������1�+���P1Ѿ�>@�Z�SM�G0��=�JG�`S�CL�͵SPH_D�@��%;0u� RTER`  �< SA_�@G1"�A�@�c��\$DI�
"2{3UDF  ǀv~ LW�(VELq�IN�b)@� _BL �@u��$G�q�$�'�'p�%`<�� ECHZR�/�TSA_`� %���E}`<����5��Bu� 1}`_�� �)5D2d%��A4I�1�N9t&pPDH�A�:��ÀP$V `�#>A$��ł�+$Q�pR}ӆ���H �$BE�Lvᵆ<!_ACC�E�!c��7/��0IR�C_] ��pNT<T��S$PS�rL� d�/Es��F{�@F
��9gGCgG36B���_�Q�2�@�A����1_MGăD1D�A]"łFW�`��`�3�EC�2�HDE�K�PPABN>G��SPEE�B�Q%_pB��QY�Y��11$US�E_��,`Pk�CTEReTYP�0�q P�YN��Ae�V)�B�QM���ѷ��@O� YA�TINCo�ڱ�B��DՒ�WG֑ENC�����u�.A�2Ӕ+@INPOQ�I6Be���$NT�#�%NT2c3_�"�2IcLO� �2_`��I�_�if� @_�k�? �` ej�C400fMOSI�A������A䃔�PERCH#  �c��B" �g� �c��lb=�����oUHu@�@	A6B(uLeT 	~�1eT�ljgv�fgTRK@%�AY�� "sY��q6B�u�s۰�8]��RU�MOMq�Ւ�Y�MP�^��C0�s�CJR��DUF �B�S_BCKLSH_C6B)����f���S�t�H��RR��QDCLALM-d���pm0���CHK���GLRTY���d��Y�8��)Üd_UM]�ԉ�C��A!�=PLMT� _L�0��9��E�.� ��#E)��#H� =��Q3po�xP	C�axHW�頿Eׅ�CMCE��@�GCN�_,ND�Ζ�SF�1�iVoR��g<!���6B���CATގSH)�,�DfY��f`��7A���܀PAބ&�R_P݅�s_ ��v���s����JG��T]���Y�����TORQUaP��c�yPOU��b��P%�_W�u�t��1D��3�C��3C�IK�IY�I�3F�6�����@�VC�00RQ�t��1࿾�@ӿ��ȳJRK������UpDB Ml��UpMC� DL�1BrGRVJ�Cĭ3C��3$�H_��"�j@q��COS~˱~�LN ���µ�ĭ0����� u����̓��Z���f$�MY��؊��˾>�THET0reN�K23�3hҧ3��C�Bm�CB�3C! AS� ��u��ѭ3��m��SB�3��x�GTS$=QC�������<����$DU��Kw��B�%(��%Qq_ ��a��x�{�K���b(��\�A`Չ��p�{�{�LPH~�g�Aeg�Sµ��������g������֚�V��V���0��V��V��V���V��V	�V�V%�H��������G������H��H��H	�H��H%�O��O��OTV	��O��O��O��UO��O	�O�OցFg���	�����S�PBALANCE�_-�LE��H_`�SP!1��A��A>��PFULCEl�Tl��.:1��U�TO_����T1T2��22N���29` �!�qnL�=B�3�q�TXpOv 
A4�IN�SEG�2�aREV8��`aDIF�uS9�1�8't"1�tpO!B.!t�M��w2�9`���,�LCHWARLRCBAB�� ��#��`-ФQ 5�X�qP�R��&��2�� 
p�""��1eROB͠�CR6B5�� ��C�1_��T �� x $WEgIGH�P`$��d?3àI�Qg`IFYQN�@LAG�Rq�S�R� �RBILx5OD��p�`V2ST�0V2P!t�W0�01�&1/0��30
�P�2�QA � 2řd[6DEB�Ug3L_@�2�M'MY9&E Nz�D�`$D_A�a$��0��O� ����DO_@A.1� <B0�6�m�Q�IB�2�0N-cdH_p`�P��2O�� �/� %��T`"a���T/!�4)@TICYKh3| T11@%�C� ��@N͠�XC͠R�?��Q�"�E�"�E8@P�ROMP�SE~� $IR��Q��8R;pZRMAI)��Q4�R4U_r02S; t�q�PR8�COD�3sFU�Pd6ID_[��vU R!G_SU;FFu� l3�Q;Q�BDO�G �E�0�FGRr3�"�T�C �T�"�U�"�Uׁ�T8D��0�B0Hb _FIv�19*cORD�13 50�236V�+b|�Q1@$ZDT}U�s0�1;E�4 *:!L_NAmA�@�b>�EDEF_I�h�b �F�d�E�2�F�4�F�c�E�e�FISP��PAKp�Ds�C�d��44בi��2D�"�It��3D�O#OBLOCKEz��S�O�O�Gq�R�PUM�U�b�T �c�T�e�T!r�R�s�U �c�T�d�R�6�q�S � ���U�b�U�c�S�Z��X�@P` t�@qDe�)@W�x���soa�TE�<D�( }l1LOMB_���ɇ0V2VIS;�I�TYV2A��O�3A�_FRI��a SIq�QR�@��@R�3�3V2W��W��4����_e��QEAS^3�Rϡ��_�[p:R��4�5�6_3ORMULA_Iz����THR^2 �EGtg�30f��<8�5COEFF_O�A�	 ��A��GR�^3S�g0BCAnO/C$l��]3��BGRP�� � � $h�p�YBX�@TM~w����u�B�s��bCER�, Tttsd�0�  ��LL�TSpS~�_�SVNt�ߐ���0ʸ���0� ��SwETUsMEA*P��P��W0�1+b/0� g� h��  @�ڐo�l�o�cqz��bH�@cqq`tP�G��R�� Q\p*q[p��t>�c NPREC>a�t���MSKy_$|�� PB1?1_USER�e"��{ ���VEL@���{ 0�$Ō!I]`���MT�ACFG>���  �@@ =O�"NORE-0l@,o�V�SI.1�d��6��"UXK�fP!��D�E�� $KE�Y_�3�$J3OG�� SV���0���!��}�SW�"�ah\aS�ՐT|�GI����| ^�� 4 �h��'d2�!XYZ�c���31�_ERR#�� 8Ԡ�A�fPV�d��1����/$BUF��X��p`��MOR|�� HB0CUd�lA�!��GQ�\aB�,"!a$�� ���a�����_�?�G~�� � �$SIՐ���V�O��T� OBJE<_��ADJU)B�ŏELAY���%�DR�OU.`=ղВQ0b=��T���0���;BDIR���; 8I�"0DYNW�#���T��"R���@�0��"�OPWORK����,%@SYSsBUy�SOP�H��ޑ�U�; P�pN�<�PA�t�>�"V��OP�PUd!0��`!��l�IMAGbw�B0y�2IM��ƕ�INe�d��RGOVRD��-��o�Pq��0��J�Os����"L�pBa���o�P�MC_Ee`���1N"y M A�21�2����SL_��� � $OVSL����?q�`��2�" -�_��k�P��k�Pu���2�C� �`��x����_ZER��D��$G�� �2=���� @h*���%O~PRI��� 
JP8+u�T=!/�L��ح�T� ަ0ATUS��TRGC_T���sB�� }fs�9s�1Re`���� DFAm����L����"��0a� ޱ��X�Ew{�����C0vUP��+p	qCPXP�j�43 ^� �PG\���$SUBe�%�q�e9JMPWAI�T z}%LO��F<�A�RCVFBQ�@�x"�!R�� �x"AC�C� R&�B�'IG�NR_PL9DB�TB�0Pqy!BW�bP�$w�Uy@�%IG�T�PI��TNLND�&2R��rL�NP���PEED \HADOW�06�w���E[q4jO!�`SP]DV!� LbAz�p�`�07�3UNIr�ȡ�0"!R��LY�Z`� ou�PH_�PK��e�RETGRIE9{�q�/��0'PFI"�� �xG`�0D 2�g��DBGLV�#LO�GSIZ��EqKT��!U��VDD�#$0_)T�G�MՐCݱ���|@eMRvC}�3�CH�ECK0���P�O�V!�k�I��LYE(!��PArpT�2�K�W��@P2V!� h $ARIB iR� c�a/�O�P8�ӐATT��2�IF`|@z�Aq4S�3UX��̊�2LI2V!� y$g���ITCHx"Z[�W �AS9��wSLLBV!��_ $BA�DYs��BAM!���Y9��PJ5��Q��R6|�V�Q_KNOW�C4b��U��AD�XV��0D�+iPAYL#OAt��Ic_��Rg��RgZOcL�q��P�LCL_�� !�7��b�QB��d��
�fF�iC֠�js��d
[�I�hRؠ�g�Ңd�B����J��q_Jt�a#���AND���Ĳ.t�b�a�q�PL~0AL_ �P��0���QրC��D:NcE���J3CpWv�� TPPDCK�������P�_ALPHgs�sBE��g�y| �K�1�� �� ���HoD_1jOj2ydDP�AR��*��;�&���TIA�4U�5U�6��MOM��a���n���{�Y�B� ADa���n���.{�PUB��R��҅ n�҅{�O2�Wp��W _�  PMsb�T� �BxQ���� e$PI�� 81��TgJ��niJ�IV�Id�Ir��[��3!��>!��r��8��U3HIG�SU3 �%�4얎4�%� ����"����!
��!�%SAMP���^��_��%�P4s ю��� [ 	ӝ�3 ���0��� &�C�����^��Sp��H&0	�IN�SpB� ���뤕"��6��6�^V�GAMM�Sy�I�� ETْ��;�D��tA�
$ZpIBRt!62IT�$HIِ!_���C�˶E��ظ1AҾ���LWͽ� 
���7���rЖ,0�q�C�%CHK��" 7�~I_A��� ��Rr�Rqܥ�Ǚ��������Ws �$^�x 1���I7_RCH_D�!� cRN{��#�LE��ǒ!,��x���90M�SWFL�$�SCR((100��R@��3]B��ç��a����ټ�0��PI3A9�METHO����%��+AXH�XX0԰N62ERI��^�3��IR�0$u	��pF{�$_���?ⲣ1�L�qL�_�a�OOP��p��wᲡ��APP:���F���@{���أRT�V�OBp�0T�`���;��� 1�I�`�� ��r���RA�@�MGA1���SSV�-��P�CUR�g�;�GRO[0S�_SA�Q��Y�#NO�pC!"�tY� �Zolox�������!bX����&�DO�1A�� �A����Х��A���A`"�WS�c �q�wPM)�� � F��YLH�qܧ��ASrZ�]B�o�=�Pq�õq_�C1�N�M_W���g����c�M� �`Vq�$p�x1o�3"�P9MJ�,�� �'A� d9�!Wi:�$�LWQ|ai�tg�tg �tg{t� �N`��(�S��SpX�0O�sRq�Z��P� *�� �
��M���������� ����X��� ��@!��q_~R� |�q#(Y� ���&n��&{�Y�Z��'��&t��Q��qU�"0��ҏ }`�$PQ�P�MON_QUc� �� 8�@QCO�U��%PQTH��H�O�^0HYS:PES�R^0UEI0O��@]O|T�  �0PG�õz�RUN_TO�� �0ْ.�� �PE`�5C��A<�I�NDE�ROGR�AH�� 2g�NEg_NO�4�5IT���0�0INFO�1�� �Q�:A��e��1IB� (��SLEQݖFAѕF@�6�eOSy�T� =4�@ENAB��0�PTION.S%0ERVE���G��A0zCwGCF�A� @R0�J$Rq�2���R��H�O�GqPxA_EwDIT�1� �vR�K�ޓʱE�sNU0W*XAUTu�-UCOPY�ِN\����MѱNXP\[qƯPRUT9� _RN��@OUC�$G��2�T��$$sCL`?0����k��a�a� �Pr�S�@�X�P�XK�QIRTU���_�PA� _WRoK 2 e�@� 0  �5��QMoYhJo|m |l	�`�m�oa�B`��o�o�f�e�l }�aI[ct'`sBS�*� 1�Y� <7 �������&� 8�J�\�n��������� ȏڏ����"�4�F� X�j�|�������ğ֟ �����0�B�T�f� x���������ү��� ��,�>�P�b�t����������srCC��L�MT?0���s  dѴINڿ�дPRE_EXE��)�Ƅ0jP��zaV'`DV��S�@e�)�%sele�ct_macro࿿��kϤ�qtIOC�NVVB�� ��P���USňw���0Vw 14kP $$p���a�|�`?� ��߰>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p�������� ��$�ѰL�ARMRECOV� ^�����L�MDG ��Ь�LM_IF ���d  Y�ST-040 O�peration� mode AU�TO S��ed �(TELEOP) �� ����9�K�]��o��, 
 ����#�8� ǘL�INE 6ǑقP�A��DǙJOINT 100 %�����$��1�@��$�@��ATAǒ0ǐ3���������  clear�䀪���ί��NGT�OL  @� 	� A\���ѰP�PINFO �� f�L�^�p����  ������k� ��ۿſ�����5��`Y�C�iϏ�%���ٯ ����������'�9��K�]�o߁ߓߙ�PP�LICATION� ?t���|�Han�dlingToo�lǖ 
V9.�40P/17\��
883ǀ����F90�	�549����|����7DF5�м��ǓNone���FRA�� �ؒ��,�_ACTI�VE1�  �� � s ��ڀMOD���������CHGAoPONL�� ��OUPLED 1	��� >�B�T��f���CUREQ �1
��  Tp�
p�p�	�������� l�������������xi3l�p�g���^H���A�t
HTTHKY�FXv|�� *<N`�� ������// &/8/J/\/�/�/�/�/ �/�/�/�/�/?"?4? F?X?�?|?�?�?�?�? �?�?�?OO0OBOTO �OxO�O�O�O�O�O�O �O__,_>_P_�_t_ �_�_�_�_�_�_�_o o(o:oLo�opo�o�o �o�o�o�o�o $ 6H�l~��� ����� �2�D� ��h�z�������ԏ ���
��.�@���d��v�����������TO������DO_CL�EAN���E�NMw  �� p��������ɯۯv�DS�PDRYRL���H	I��o�@��G�Y�k� }�������ſ׿���8�ϻ�MAX��,�����=�X,���9�|����PLUGG,�-�9���PRC��B�m�q�6�(ϗ�Ox����SEGF�K���� �m��G�Y��k�}ߏ�����LAP $�7ޡ������+� =�O�a�s�����> �TOTAL_ƈɾ �USENU$��1� ������RGDISPMMC�ed�C�O�@@��1�O"�D��-�_�STRING 1���
�M���S��
��_I�TEM1��  n ��������� $ 6HZl~��������I�/O SIGNA�L��Tryout Mode���InpNSim�ulated���Out`OV�ERR!� = 1�00��In c�yclT��Prog Aborj���JStatu�s��	Heart�beat��MH� Faul��Aler�!/!/3/�E/W/i/{/�/�/�/ (���(����/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O84OFO�/WORИ� ~A�/XO�O�O�O�O�O  __$_6_H_Z_l_~_��_�_�_�_�_�_�^PO���"`�KoEo Woio{o�o�o�o�o�o �o�o/ASepw��bDEV%n �p9o����#�5� G�Y�k�}�������ŏ�׏�����1�C�PALT�-j��OD� ������ȟڟ���� "�4�F�X�j�|�����p��į֯X�GRIB� ������6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�z�����R�-��&������� ���"�4�F�X�j�|� �ߠ߲����������<��PREGn�W� ��0�~�������� ����� �2�D�V�h��z���������$�$�ARG_~@D ?�	�����  	�$$	[]��$:	��SBN_CONFIG��XWqRC�II_SAVE � $zm��TC�ELLSETUP� 
%  O�ME_IO$$%?MOV_H� ���REP��#��U�TOBACK� �	tFRA;:\D� .D�z '`�D�w� �s  �25/11/2�9 20:26:16D�;D���#//h��C/j/|/ �/�/�/�/D�X/�/ ??(?:?L?�/p?�? �?�?�?�?�?g? OO $O6OHOZO�?~O�O�O�O�O�O�O���  �c_F_\ATB�CKCTL.TM��)_;_M___q_8INIm��j~C?MESSAG� �Q�z �[ODE_D(� �j�XO�p�_�@PAUS6` !�� , 	��; :oHg,		2oloVo�ozo�o �o�o�o�o�o 
D�.Pz}d`TSK�  mw}_CUgPDT�P�Wd�p��VXWZD_ENqB�Tf
�vSTA�U��u��XISX UONT 2�vwy �� 	 �:�� �� �,�i�> ��`�y_D�R����0������ ���m�����R�����k\�;�� B� ����╏�yp����.�1�MET���2@��y PQ�A��Q�A��A�`%�A�Ah�A�����>��>iHw�>yK�?
0[�?��?	�8�5�SCRDCFG� 1Y; �� ���%�7�I�pD�Q ��ݟ������Я��� [���<�N�`�r���`����7���FGR9���p�_ԳPNA� �	FѶ_ED��P1��� 
 ��%-PEDT�-¿ R�v���E��<�GE�D�;�9/�>���  ����2�����B� ��ˀ�{�����j�����3 ��#� �G�Y���G����6�����4����� �Yި��Z�l������5K������Y�t�@��&�8���\���6 ��d��Y�@����(��7�S0w Y�w��f���!8�W��{�IZ��@C/��2/���9{/��//LZݤ/?V/0h/�/�/��CR�� �?�?Tn?�? ?2?�?�V?԰!�NO_DE�L�ҲGE_UN�USE޿дIGALLOW 1��   (*SYSTEM*
��	$SERV_�GR[�@`REGƜE$�C
��@NU�M�J�C�MPMU|?@
�LAYK��
�PMPAyL�PUCYC1����L4]P!^YSUL�SU_�M5Ra�C�Lo_�TBOXOR=I�ECUR_�P�M�PMCNVV��P10I^�PT4�DLI�p�_�I	*�PROGRA�D?PG_MI!^KoF]`AL+ejoTe]`�B�o�N$FLU?I_RESU9W�o�O�o�dMR�N�@�<�?�;M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3��E�W�2BLAL_OUT �K���WD_ABOR:P�cO��ITR_RT/N  �$�빸�?NONSTO��� lHCCFS_UTIL ��̷CC_AUXA�XIS 3$� h}�j�|�����ƽ�CE_RIA_IL`@�נ��FCFG $��/�#��_LIMv�B2+� �8p7� 	��B\���$�8p
Ԡ��)�Z��%�/����� [�����.R���!����	�L��(
5������PA�`GP 1H�����A�S�e��w�6�CC� C7���J��]��p�������� C����������������ê��̩�ձ�ߩ��*�������;���PSCk����������U���������ɱ���������� �D� D!�j!�!�!� ��&�?��HE@ON�FIpC�G_Pv�P1H� +E H��ߟ߱���������|�C�KPAUS�Q31H�ף b� S�H�A��e���� ����������E�+�@i�{�a���A?I�ץ�MؐNFO �1��� �3��$4�A��A_�e�T���?3�L�����* �D58o�G���C˃]�3�����n�����bPb�O� �� ��LLECT�_�!�����E�N+`�ʒ���ND�E�#�/��1234567890�"�A��$/ҵHw��#)j� �<i{��;��/ ��/`/+/=/O/�/ s/�/�/�/�/�/�/8? ??'?�?K?]?o?�?��?�?�?O�?��$ο ��IOG &��"S�`�O�O�O�O`GTR�2'DM(��^�?�N�N�(oM Z��_�MOR)q3)H�� 7ىU3��Y�_�_�_�_��_�[bR�kQ*H�,�S�?<�<Ѡ<c8pK(Fd���P,��;ϒo�o�o˿�o�o(œh�UY@E�o�S �sj]a�PDB.����4cpmidbag3��Рs:��>�uqpz��v  �CAx��}`.��}�`��|�<�CmgP���t��~f�������@ud1�:�?��XqDEFg -��zC)*��cO�buf.txAtJ��|K�[`�/DM=��>���R�A6��MCiR20_{RC�d���hS21����G���CzA�d4��EI�jA��]�C-]�G/X"B�e;F]��H�j�C1�a�F�%J��i�E&�mI؂��LڒYF���I�!oN���mH�?aMSo<����>׼_N��6f23DLD�	>�	P!� 2��}���yc
�@x9� C}�Ĵ  D4G��E���  E�%q�F�� E�p�u�F�P� E��fF�3H ��G�M����?5�>�3#3��?�xn9�q@�Q5����Rp�A?a��=L��<#�QU�@,�C������RSMOFS�T +i�����P�_T1Ɠ4DMA� =ք�MODE 35dm�@��	Q�M;��%��?����<�M>���Ͷ�TESTRc�2i�`�R�6�O�K�CN�AB���n�E 8��\�n�Cd�B���Cpp�����	P:d�QS ��� ������*4�I7>���>B�8m5$�RT_�c�PROG %�j%��d�1�h@NU�SER��x�KEY_TBL  e������	
��� !"#$%�&'()*+,-�./(:;<=>�?@ABCc�GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������>��͓���������������������������������耇����������������������4A8�LCK���F�y��STAT���2�X�_ALM������_AUTO�_DO�E�F�DR 3:i�2�h&q[~�� �BUOSYST�-322 Aut�o status� check t�ime out ����i�$TE�LEO8�i� ���)qA�ʜ�@Ĭ������?�ڛMs�B�õ�?*�?��?Mf�=�o�TR���-���D�.�B���C����B�N�*p��4�N4�J5Hj5H��>�i�IBJ�d�BF�	PZ��[~�bbt��p��5/�M*F��B�GA+$����@R���J�}BQ�H�����������2>���@�@����&�CBxH�CKH<B��6 >Tbt��/���u�US�H?Z?l?i�$ 7?�?:�� mϸ?�?p ���?�?OO�?,OfO xO�M6?�O�O�O~?�O 	_�?*_$_BOD_6_p_ ~_T_�_�_�_�_�Oo )o;o�OLoqo_�o�o �_�o�o�o�o�o�o FXo��No� ��o����@� N�$�b�x�����n� �����A��b�\� z�|�n�������ʟ�� �(�֏O�a�s���� ��T�ʯį��֯� ���2�H�~���>��� ɿۿ���ϼ�2�,� J�L�>�xφ�\Ϛϰ� ���Ϧ��1�C��T� y�$Ϛߔ߲ϴߦ��� ������N�`�߇� ���V߼������� ���H�V�,�j��� ����v�����$ I��jd���v� ����0��W i{&��\�� ���/&/�:/P/ �/�/F�/�/�/��/ ?�:?4?R/T?F?�? �?d?�?�?�? O�/'O 9OKO�/\O�O,?�O�O �?�O�O�O�O�O
_ _ V_h_O�_�_�_^O�_ �_�O
oo"_$ooPo ^o4oro�o�o�o~_�o 	�_,Q�_rl �o�~����� &�8��o_�q���.�� ��dڏԏ��� � .��B�X�����N�ǟ ٟ럖���!�̏B�<� Z�\�N�����l����� �����/�A�S���d� ��4�����¯Ŀ��� ��Կ�(�^�p���� �ϻ�f����Ϝ��� *�,��X�f�<�zߐ� ���߆����#���4� Y��z�t�ߔ���� �������.�@���g� y���6����l����� ������(6J` ��V������ )��JDbdV� �t���/�7/ I/[/l/�/<�/�/ ��/�/�/?�/?0? f?x?&/�?�?�?n/�? �?�/OO2?4O&O`O nODO�O�O�O�O�?_ _+_�?<_a_O�_|_ �O�_�_�_�_�_�_ o 6oHo�Ooo�o�o>_�o �ot_�o�oo�o0 >Rh��^o� ���o�1��oR�L� jl�^�����|���Џ ���?�Q�c��t� ��D�����ҏԟƟ � ��"�8�n���.��� ��˯v�ܯ���"�� :�<�.�h�v�L����� ֿ迖��!�3�ޯD� i���τϢ��ϖ��� �ϴ����>�P���w� �ߛ�FϬ���|����� 
����8�F��Z�p� ���f��������� 9���Z�T�r�t�f��� �������� ��G Yk�|�L��� �����*@ v�6���~� 	/�*/$/BD/6/p/ ~/T/�/�/�/�/�? )?;?�L?q?/�?�? �/�?�?�?�?�?�?O FOXO?O�O�ON?�O �O�?�O�OO__@_ N_$_b_x_�_�_nO�_ �_o�OoAo�Obo\o z_|ono�o�o�o�o�o (�_Oaso� �To���o��� ��2�H�~���>�� ɏۏ����2�,� J�L�>�x���\����� ������1�C��T� y�$������������ �į��N�`���� ����V���ῌ���� ���H�V�,�jπ� ����v����߾�$� I���j�d߂τ�v߰� �ߔ������0���W� i�{�&ߌ��\����� �������&���:�P� ����F���������� ��:4R�TF� �d��� ��' 9K��\�,�� ������
/ / V/h/�/�/�/^�/ �/�
??"/$??P? ^?4?r?�?�?�?~/�? 	OO�/,OQO�/rOlO �?�O~O�O�O�O�O�O &_8_�?__q_�_.O�_ �_dO�_�_�O�_�_ o�.ooBoXo�otc�$�CR_FDR_C�FG ;re��Q
UD�1:�W�P�aJ�d � �`�\�bHISoT 3<rf  �`  ?�RW@tAtB�bWC�P1pDtUEtItg�Pp�otw�_��bIN_DT_EN6p�T?�q�b�T1_DO  ��U�u�sT2��wV�AR 2=�g�p hq  o8s��s��R6�t(4�t(�m[�z�RZ�`STOP���rTRL_DEL�ETNp�t ��_�SCREEN �re�rkcs�c�rUw�MMEN�U 1>��  <�\%�_��T ��R��S/�U���e� w�ğ������џ�	� B��+�x�O�a����� ������ͯ߯,��� b�9�K�q�������� ��ɿ����%�^�5� Gϔ�k�}��ϡϳ��� �����H��1�~�U� gߍ��ߝ߯������� 2�	��A�z�Q�c�� ����������.�� �d�;�M���q�������������YӃ_M�ANUAL{��rZCD�a?�y�rG� ���R�fx"
�"
?|(��P�dTGRP 2@:�y�B� � �s��� �$DwBCO�pRIG����v�G_ERRL�OG A��Q��I[m �N_UMLIM�s���u
�PXWOR/K 1B�8����//�}DBT;B_�� C%����S"� �aDB__AWAY��Q�GCP �r=���m"_AL�F�_�Yz����p�vk � 1D� , 
��/"�/%?/(c_M�pqw,@�=5�ONTIM���f�t�_6�)
�0~�'MOTNENFp�F�;RECORDw 2J� �-?�SG�O��1�?" x"!O3OEOWO�8_O�O �?�OO�O�O�O�O�O (_�OL_�Op_�_�_�_ A_�_9_�_]_o$o6o Ho�_lo�_�o�_�o�o �o�oYo}o2�oV hz��o��C �
��.��R��K� �������Џ?��ߏ �*�����+�b�t�� ������Ο=�O��� ��:�%���p�ߟ񟦯 ��O�ǯ�]������ H�Z���������#��5����ϩ�i"TO�LERENCv$B�ȿ"� L��� C�SS_CCSCB� 2K�\0" ?"{ϰϟ���7�� 
����@�R�d�3߈���"�x�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C�Ugy��� �������R�LL]�La�m1T#2� C�C�p�F�^ A�C�%pC���#�0�? 	 A����B���?�  ��$����\0����0��B��`#sߠK/]/o/�ϓ/��/�/s/�/�/�K��:�L��q����e;��9|?�AȦ��/�Q�/`?;�@���O?�?�?�?Ȏ0A0F��?{F�A OO��7�1���9M	AB 
AZOdBAE�9$O�O�O��Oi:P��`�@0��DJCA� @5��
X-.
[$h=�� M?�>O�ڴ �q_�_�_�_:W�A<,19\<ǲ/o�/�_+oPobotoǦeACHC�V�WB$�Dz�cD�`�a=/��o�oo�oW�a.+�!��2=t,yCE{�YqBf��I? �-t�s�js�w�yj �������Q���@`��$���� �A����Bމ�o�� '�9��_]�o�N���r� ��ɟ۟_�B�ʄ���YZ>`�$v B��w�Be�@��Z�>R�ҹ�x�Z�l�~����`_м¯��� 
���̯9�,�]�o���  �H�����ٿ뿊�� ƿ3�E�W�iϬ���$� ������ Ϟ����/� A�S߶�w�V�h߭ߌ�0�S���ߐ�_�f 	��H�?�Q�~�u�� ����������� D��-�g�q������� ������
@7�Icm��߾�  �����) M@qdv��� ����//I/P� m/�v/�/�/�/�/�/ �/�/?3?*?<?i?`? r?�?^/�?�?�?�?�? O/O&O8OJO\O�O�O��O�O�O�O�O�g	 � Q�P��s �PC4
p*p�p6U6P\�C9p/p��Q ]V^PM]�6P�:P��>P�VJ_�^P��bP�fP�Vr]v��Tp Q
k���_oob�id1Q&oNo ;o�_co�oˏUUA  � �o�k1Q@�  ��o�k�b������Up �� 1��b6�1C���C�cP�fL��?#�c>�/{���`�cP��@@�d��r�`BȲcP>�s�qC��p���b�t<�o�?�PH�)S�B�tq�q�p�r�`CB���eIC�&��Q�4( �oz�UU�D��xz9���=�@>R�����zQ�-R������EE��_�B��3�b��`ځ`  ?�p��<�U�[?���}t���$���$DCSS�_CLLB2 2=M��p�P��^?�NSTCY �2N���  ������� ʟ؟���� �2�D� Z�h�z�������¯ԯ���SA�DEVIC/E 2O��!�$��4&V�h������� ˿¿Կ���
�7�.� [�R�ϑϣϵ������4(A�HNDGD 3P��*�Cz�A�_LS 2Q��_� Q�c�u߇ߙ߽߫����?�PARAM �RP��1�`�&�RB�T 2T�� �8�P<C�'p ��qi�l��s@"��R��(qI�X��0��pB CW  ��B�\x�N��`Z����	%��)���X�j��p�����zq�����B �(s,�F�p�V��`q���b��B ��4&c �S�e�l�4+�����H1~����=D�C�$Z��b����A,� 4��u@�X@���^@w���]B�B�cP%���C4�C3:^�C4��nЬ ���p8�-B{�B��A����� l��C��C3�JC4�jC3��yn+��3 Dff 2�GA PB W4+@:� ]o�W���� �/�/P/'/9/K/ ]/o/�/�/�/�/?�/ �/�/?#?5?�?Y?k? �?�?�o�?�?O�?6O !OZOlOWO�O�Es�? �?�?�O�O_�O�OL_ #_5_G_Y_k_}_�_�_ �_ o�_�_�_oo1o ~oUogo�o�o�o�o�o wO D/Aze ����O�o�o
��o ��R�)�;���_�q� ���������ݏ�<� �%�r�I�[�m����� ���ǟٟ&�8��\� G���k�������گů �����F��/�A� S�e�w�Ŀ������ѿ �����+�x�O�a� �υϗϩϻ�����,� ��b�t�ﯘ߃߼� ����������:�� C�U߂�Y�k���� ��������6���l� C�U�g�y��������� �� ��	-?Q ������� @+dvQ�� ������*// /%/r/I/[/�//�/ �/�/�/�/&?�/?\? 3?E?�?i?{?�?�?U �?�?"O4OOXOCO|O gO�O{��?�O�?�O �O0___f_=_O_a_ s_�_�_�_�_�_o�_ oo'o9oKo�ooo�o �o�o�o�o�O:% ^I�������H�$DCSS_�SLAVE U����	����z_4D  �	��AR_ME_NU V	� ��j�|�������ď�B�Y�� ��~?�SHO�W 2W	� � �b�aG�Q�X�v� ��������П֏���� @�:�d�a�s��� �������߯��*� $�N�K�]�o������� ̯ɿۿ���8�5� G�Y�k�}Ϗ϶����� ������"��1�C�U� g�yߠϝ߯������� �	��-�?�Q�c�� s������������ �)�;�M�t������ ����������% 7Ip�m������ ����!3Z Wi���J�� ��//DA/S/e/ ��/��/�/�/�/�/ ?./+?=?O?v/p?�/ �?�?�?�?�?�??O 'O9O`?ZO�?�O�O�O �O�O�OO�O_#_JO D_nOk_}_�_�_�_�_ �O�_�_o4_.oX_Uo goyo�o�o�o�_�o�o �ooBo?Qcu����o:���C�FG X)��3�3q5p�F�RA:\!�L+�%04d.CSV|�	p}� �qA- g�CHo�zv�P	����3q������́܏� ���4��GJP����qp�1� �RC_OUoT Y���C��_C_FS�I ?i� .�������͟ �����>�9�K�]� ��������ίɯۯ� ��#�5�^�Y�k�}� ������ſ����� 6�1�C�U�~�yϋϝ� ���������	��-� V�Q�c�uߞߙ߽߫� �������.�)�;�M� v�q��������� ���%�N�I�[�m� ���������������� &!3Eni{� ������ FASe���� ����//+/=/ f/a/s/�/�/�/�/�/ �/�/??>?9?K?]? �?�?�?�?�?�?�?�? OO#O5O^OYOkO}O �O�O�O�O�O�O�O_ 6_1_C_U_~_y_�_�_ �_�_�_�_o	oo-o VoQocouo�o�o�o�o �o�o�o.);M vq������ ���%�N�I�[�m� ��������ޏُ��� &�!�3�E�n�i�{��� ����ß՟������ F�A�S�e��������� ֯ѯ�����+�=� f�a�s���������Ϳ �����>�9�K�]� �ρϓϥ��������� ��#�5�^�Y�k�}� �ߡ߳���������� 6�1�C�U�~�y��� ���������	��-� V�Q�c�u��������� ������.);M vq������ %NI[m �������� &/!/3/E/n/i/{/�/��/�/�/�/�/�/3��$DCS_C_F�SO ?����71 P ??T?}?x? �?�?�?�?�?�?OO O,OUOPObOtO�O�O �O�O�O�O�O_-_(_ :_L_u_p_�_�_�_�_ �_�_o oo$oMoHo Zolo�o�o�o�o�o�o �o�o% 2Dmh z������� 
��E�@�R�d����� ����ՏЏ���� *�<�e�`�r������� ��̟�����=�8��J�\�������?C_RPI4>F?��� ����3?�&�o���,�� >SLү@d��� ���%�7�`�[�m� Ϩϣϵ��������� �8�3�E�W߀�{ߍ� ������������� /�X�S�e�w���� ���������0�+�=� O�x�s����������� ��'PK] o������� �(#5Gpk} �����Q���/ 6/1/C/U/~/y/�/�/ �/�/�/�/?	??-? V?Q?c?u?�?�?�?�? �?�?�?O.O)O;OMO vOqO�O�O�O�O�O�O ___%_N_I_[_m_ �_�_�_�_�_�_�_�_ &o!o3oEonoio{o�o �o�o�o�o�o�o FASe�������>�NOCOD�E ZU���?�PRE_C�HK \U��pA� �p�<� ��pU�]�o�U� 	 <Q�������� ۏ�Ǐ�#����Y� k�E�����{�şן�� ß����C�U�/�y� ����s���ӯm���	� ��?��+�u���a� ������ɿ�Ϳ߿)� ;��_�q�K�}ϧϝ� �����ω���%���� [�m�Gߑߣ�}߯��� �����!���E�W�1� c��g�y�������� �����A�S�-�w��� c������������� +=asM_� �����'� ]o	��� ���/#/�G/Y/ 3/e/�/i/{/�/�/�/ �/?�/?C?9Ky? �?%?�?�?�?�?�?	O �?-O?OOKOuOOOaO �O�O�O�O�O�O�O)_ ____q_K_�_�_a? �_�_�_�_o%o�_Io [o5oGo�o�o}o�o�o �o�o�o�oEW1 {�g���_�� ��/�A��M�w�Q� c����������Ϗ� +���a�s�M����� ����ߟ���'��� 3�]�7�I������ɯ ۯ�������G�Y� 3�}���i���ſ���� ����1�C���+�y� ��eϯ��ϛ������� ��-�?��c�u�Oߙ� �߅ߗ��������)� �M�_�U�G���A� ������������I� [�5����k������� ������3EQ {q���]�� ��/AewQ �������/ +//7/a/;/M/�/�/ �/�/�/��/?'?? K?]?7?�?�?m??�? �?�?�?O�?5OGO!O 3O}O�OiO�O�O�O�O �O�/�O1_C_�Og_y_ S_�_�_�_�_�_�_�_ o-oo9oco=oOo�o �o�o�o�o�o�o_ _M_�ok�o� �������I� #�5����k���Ǐ�� ӏ��׏�3�E��i� {�5c���ß����� ӟ�/�	��e�w�Q� ������ѯ㯽�ϯ� +��O�a�;������� �Ϳ߿y����!� K�%�7ρϓ�mϷ��� ����������5�G�!� k�}�W߉߳ߩ����� �ߕ��1���g�y� S���������� �-��Q�c�=�o��� s����������� ��M_9��o� ����7I #mYk��� ���!/3/)/i/ {//�/�/�/�/�/�/ �/?/?	?S?e???q? �?u?�?�?�?�?OO �?%OOOE/W/�O�O1O �O�O�O�O__�O9_ K_%_W_�_[_m_�_�_ �_�_�_�_o5oo!o ko}oWo�o�omO�o�o �o�o1UgA S������	� ���Q�c�=����� s���Ϗ�o������ ;�M�'�Y���]�o��� ˟����۟�7�� #�m��Y��������� ���!�3�ͯ?�i� C�U�������տ��� ����	�S�e�?ω� ��uϧ��ϫϽ�������$DCS_�SGN ]	��E��-����30-NOV-2�5 19:W����29R�20:2�7_�x�x� /[}�t��q�т��xҚك�JѨ�E���Þ� ������  1�HOW �^	�� x�/�VERS�ION =�V4.5.2���EFLOGIC �1_���  	�����C��R�%��PROG_ENB  ��:�{�s�ULSE  X����%�_ACCL{IM������d��WRSTJN�T��E��-�EM�O|�zя�$���IN�IT `2�����OPT_SL �?		�	�
 	�R575��]�7�4b�6c�7c�50��1���C���@�TO  L���� �V�DEX��d�E�x�PATHw A=�A\�k}��HCP_CLNTID ?�:� D�ռ���IAG_GRP� 2e	�����z�	 @��  
ff?a�G���B�  2��/�8[I�@c�ς!�7�@�z�@^��@
�!��m�p2m15 89�01234567�����  �?��?�=q�?��
?޸R�?�Q�?���?�����(��?�z���x�@o�  A_�Ap ,!7A�88_�;B4�� ��L��x�
�@�@���\@~�R@�xQ�@q�@�j�H@c�
@�\��@U�@Mp��//'$��; �O)H��@C�t >d 9��@4��/\)@)� #�t {@���/�/�/�/�/P'?�/��?���_ �?}p�?u�?n{?s ?\�Q�? ?2?D?|V?h8�
=?��鎌0w5�z�H�?p�h��?^�R�?�?�?�?�?h8���t0���,@�?��0�;@ &O8OJO\OnOP'�$_ �_Y_k_�O?_�_�_ �_�_�_s_�_�_1oCo !ogoyoo�o��Bj"�� �2{1�@"?�Ś�f�t0�d"5!{�
u4V��u@"�B3t�A>u��?�@[q��@`,=q��=b��=��E1>�J�>��n�>��H"<w�o �z�s�q���� �x�C�@<w(�Uz� 4i�� ����A@x�?*�o��m*�P�b� ��tn���2���Ώ��x���i>J��&��bN2�"��GI�N��o@�@v���0y����@ffr9!l ��33����(��"C�� �ƒI�CH�)�C.dBت "8"����'��� "~�A?�&"K����pf�B��@�p��������p��? �����	=������곿��Z�ơ5�g����D�58o�G��C˃]x�> �������0��N�T������3����n����b���� ÿ���ҿ��Ϥ���<�o��CT_C�ONFIG f���|�e�gY��STBF_TTS��
�������}���1�MAU�������MSW_C5F��g�  # �ڿOCVIEW��h!�-���s߅� �ߩ߻��ߟ�a���� �,�>�P���t��� �����]�����(� :�L�^���������� ����k� $6H Z��~����� �y 2DVh �������v�KRC�i���!� ��/S/B/w/f/�/�/��/��SBL_FA?ULT j*6�>�!GPMSK���'���TDIAG ik��-�������UD1: 6�78901234A5I2��=1�Ǥ�P\� �?�?�?�?�?�?�?O O'O9OKO]OoO�O�O �Od696���r
t?�O>|�TRECP"?4:
B44_[7��s?p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�O��O�O�o7�UMP__OPTIO=��.F�aTR����)u�PME��Y_T�EMP  ÈW�3BC�gp�B�QtUNI����gq��YN_BRK �lL�7�EDITO�R�a�a@�r_
PE�NT 1m) � ,&TELGEOP^P ����p�PSNA�:�&MTPG�p+�=� �/��I�z�����ۏ ����5��Y�k�R� ��v���ş���П� ���C�*�g�N�v��� ���������ޯ���?�Q���EMGDI_STAzuV�gq��uNC_INFO� 1n!��b����X���������n�1o!� ��o���
�
�d�oU�g�y� �ϝϯ���������	� �-�?�Q�c�u߇ߙ� �߽��� u����
�� *�B�*�P�b�t��� �����������(� :�L�^�p��������� 2�������9�C Ugy����� ��	-?Qc u�������� //1;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?��?�?�?O)/O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�?�?�_ �_o�_3O=oOoaoso �o�o�o�o�o�o�o '9K]o�� ��_�_����+o 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y��������ӟ ���	�#�-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� �7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߹��� �������%�/�A�S� e�w��������� ����+�=�O�a�s� �������������� �'9K]o�� ������# 5GYk}�	�� ����/1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?��?�?�?�? /O)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�? �_�_�_�_O�_!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew��_�_��� �o�+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o���� ���ɟ۟���#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� ���߹���������� %�7�I�[�m���� �����������!�3� E�W�i�{��߇����� �����/AS ew������ �+=Oas ����������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?���?�? �?�?��?OO1OCO UOgOyO�O�O�O�O�O �O�O	__-_?_Q_c_ u_�?�_�_�_�_�?�_ oo)o;oMo_oqo�o �o�o�o�o�o�o %7I[m�_u� ���_���!�3� E�W�i�{�������Ï Տ�����/�A�S� e��������u�� ����+�=�O�a�s� ��������ͯ߯�� �'�9�K�]�w����� ����ɿ�����#� 5�G�Y�k�}Ϗϡϳ� ����������1�C� U�g߁��ߝ߯���ۿ ����	��-�?�Q�c� u����������� ��)�;�M�_�y߃� ������������ %7I[m�� �����!3 EWq�c����� ����////A/S/ e/w/�/�/�/�/�/�/ �/??+?=?O?i{ �?�?�?�?��?�?O O'O9OKO]OoO�O�O �O�O�O�O�O�O_#_ 5_G_�?s?}_�_�_�_ �?�_�_�_oo1oCo Uogoyo�o�o�o�o�o �o�o	-?Qk_ u����_��� ��)�;�M�_�q��� ������ˏݏ��� %�7�I�cQ������ ���ٟ����!�3� E�W�i�{�������ï կ�����/�A�[�� �$ENETM�ODE 1p����  
k�k�f�����j��OATCFG �q�����Ѵ��C���DAT�A 1rw�Ӱ�.��*	�*��'�9�K�]�l�dlύ�e��ϻ�������� �'ߡϳ�]�o߁ߓ� �߷�1���U����#� 5�G�Y����ߏ��� ��������u��1�C� U�g�y������)��� ����	-����c�u�����j�RPOST_LO��	t�[
׶#5�Gi�RROR_P-R� %w�%L��XTABLE  w�ȟ�����RSEV_NUM� ��  ����  �_AUT�O_ENB  ����X_NO5! �uw���" W *�x �x �x 	�x + +w �/�/�/�Q$FLTR=/O&H�IS#]�J+_A�LM 1vw� e�[x,e�+�/�Q?c?u?�?�?�?�/_\"W   w�v!����:j�TCP_V_ER !w�!x޻?$EXT� _R�EQ�&�H)BCSsIZKO=DSTKhI�f%�?BTOL�  ]Dz�"��A =D_BWD��0�@�&�A���CDI�A wķ���]�KSTEP�O�Oj�>POP_DO�Oh��FDR_GRP s1xw��!d 	�?x�_��yPs�Y�Q�'�M"����l��T� ����VyS�_�]��TA�IZ�Rg���@���A^���_�P��PA8{��eAS��o Eo�_Bo{ofo�o�o�o��o@ICm@���?�=�����n
 M;�q a�a]?&:<  !�4:�o^I��X�A@�P�t@S33�uh}@�q�g��yPF@ ��|yP�G�  @�Fg��fC�8RL��}?�pi��~6�X�����875t���5���5`+���~3wM��q�� 
g ".���bY ��FEATURE� y���@���HandlingTool ��]Engli�sh Dicti�onary�4Dw St��ard���Analog �I/O>�G�gle� ShiftZ�u�to Softw�are Upda�te�matic Backup����ground �Edit ��Ca�meraU�FY�CnrRndIm����ommon calib UI���nˑ�Moni�tor$�tr�R�eliabn��D�HCP �[�ata Acquis3�~\�iagnos���R�v�isplay~ΑLicensZ��`�ocument? Viewe?�^��ual Chec�k Safety���hancedh���s�Frܐ��xt. DIO� /�fi��@�en]d�Err>�L���\�4�s[�rP�K� ��@
�FCTN M�enu��vZ���T�P In��fac<ĵ�GigE־��Đp Mask �Exc�g=�HT�԰Proxy S�v��igh-S;pe�Ski�� ����O�mmunicn��onsV�ur���q�V�ײconn�ect 2��nc=rְstru!��ʒ��eۡ��J��X�K�AREL Cmd7. L�ua��ÿRun-Ti<�E�nv�Ȟ�el +:��s��S/W�ƥ����r�Book(System)
�MACROs,M�?/Offseu�p�aHO���o�u�MR8��4���MechSt�op+�t����p�im�q���x�R������odo�witch��ӟ�.��4�Op�tmF��,�fil�䬳�g��p�ult�i-T�Γ�PC�M fun�Ǽ�o���������Regi�e�rq���riݠF����S�Num S�el��/�:� Ad�jua�*�W�q�h�t�atu��ߪ�R�DM Robot>�scove'����ea��<�Freq� Anlyq�Re�m��O�n5�����S�ervoO�!��S�NPX b-�v�SN԰Cliܡ?r��Libr&�_�� ���q +oJ�t��sGsag��X�@ �����	�@/Iս�M�ILIB��P OFirm���P���AccŐ͛TPT9Xk��eln��������orqu>o�imula=��|u(�Pa&��ĐtX�B�&+�ev.�成ri��TUSB port ��iPf�aݠ&R �EVNT� nexcept�����X%5��VC�rl�c���V���"�%q��+SR SCN�/S�GE�/�%UI	�Web Pl��>���A43��ۡ��ZD?T Applj�
�{1EOAT����x&0?�7Grid�񸾡�=�?iR�".�5� F���/גRX-�10iA/L�?A�larm Cau�se/��ed(�A�ll Smoot�h5���C�scii<+�V�Load䠌J�Upl�@w�toS� ��rityAv�oidM(�s7�t�@�ycn�����_�CS+���.3 c��XJo��� -T3_H�.RX��U����Xcollabo����RA�:�.9D���in���NR�THI
�On��e Hel����ֿ������1trU�ROS Eth$��A������;,�G �B�,�|HUpV�%�W�t ԰�_iRS�ݐ��64MB DRA9M�o�cFRO���L8F FlD�����22M �A:�opm�ԕ1ex@V�
�sh�q�"�wce�u��p��|�tyn�sA�
�%�r ����J��^�.v� P)Q/sbS�`���O�N��mai��U�h��R�q�T1�^cFC+Ԍ%̋Fs9�pˌk̋��Typ߽�FC%�hױV�N Sp�ForްK��Ԭ��lu!����cp�PG� j�֡�RJ�[L`Sup"}��֐�f��crFP��lu�� ��al�����r ��i�
q�4@а��uest,IMPLE ׀6*|HZ�p��c0�BTea(�8|���$rtu���V��9HMI�¤��U;IFc�pono2D�BC�:�L�y�p��� ������ʿܿ	� �� ?�6�H�u�l�~ϫϢ� ����������;�2� D�q�h�zߧߞ߰��� �����
�7�.�@�m� d�v��������� ���3�*�<�i�`�r� �������������� /&8e\n�� ������+" 4aXj���� ����'//0/]/ T/f/�/�/�/�/�/�/ �/�/#??,?Y?P?b? �?�?�?�?�?�?�?�? OO(OUOLO^O�O�O �O�O�O�O�O�O__ $_Q_H_Z_�_~_�_�_ �_�_�_�_oo oMo DoVo�ozo�o�o�o�o �o�o
I@R v������ ���E�<�N�{�r� ������Տ̏ޏ�� �A�8�J�w�n����� ��џȟڟ����=� 4�F�s�j�|�����ͯ į֯����9�0�B� o�f�x�����ɿ��ҿ �����5�,�>�k�b� tφϘ��ϼ������� �1�(�:�g�^�p߂� ���߸������� �-� $�6�c�Z�l�~��� ����������)� �2� _�V�h�z��������� ������%.[R dv������ �!*WN`r �������/ /&/S/J/\/n/�/�/ �/�/�/�/�/??"? O?F?X?j?|?�?�?�? �?�?�?OOOKOBO TOfOxO�O�O�O�O�O �O___G_>_P_b_ t_�_�_�_�_�_�_o ooCo:oLo^opo�o �o�o�o�o�o	  ?6HZl��� ������;�2� D�V�h�������ˏ ԏ���
�7�.�@�R� d�������ǟ��П�� ���3�*�<�N�`��� ����ï��̯���� /�&�8�J�\������� ����ȿ�����+�"� 4�F�Xυ�|ώϻϲ� ��������'��0�B� T߁�xߊ߷߮����� ����#��,�>�P�}� t����������� ��(�:�L�y�p��� ������������ $6Hul~������  �H552��2�1R7850�J614AT�UP'545'6�VCAMCR�IbUIF'28ncNRE52VwR63SCH�LIC�DOCV��CSU869z'02EIOC��4R69VES�ET?UJ7UR{68MASK�PRXY{7OCO#(3?+ &m3j&J6%53��H�(LCHR&OP�LG?0�&MHCuRS&S�'MCS>�0.'552MDS�W+7u'OPu'MP�Rv&��(0&PCMzR0q7+ 2� ��'51J51�80nJPRS"'69j&�FRDbFREQnMCN93&�SNBA��'SH�LBFM1G�82�&HTC>TMI�L�TPA�T7PTXcFELF� ��8J95n�TUTv'95j&wUEV"&UECR&wUFRbVCC
X�O�&VIPnFCS�C�FCSG��I�WEB>HTT�>R6��H;RVC�GiWIGQWIPGmS�VRCnFDGu'�H7�7R66J5t'R�8R51
(�6�(2�(5V�J8�86�L=I% ږ84g662R6�4NVD"&R6n�'R84�g79�(�4�S5i'J76�j&D0�gF xRT�SFCR�gCRX�v&CLIZ8ICMqS�Sp>STYnG6)7CTO>���7�NNj&ORS��&C &FCB�F�CF�7CH>FC�R"&FCI�VFCR�'J�PO7GBfM�8�OLaxENDS&L]U�&CPR�7LW�S�xC�STxTE�gS60FVR6�IN�7IHaF� я�����+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯۯ��� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q����������� ��%�7�I�[�m�� �������������� !3EWi{�� �����/ ASew���� ���//+/=/O/ a/s/�/�/�/�/�/�/ �/??'?9?K?]?o? �?�?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_ �_�_�_�_	oo-o?o Qocouo�o�o�o�o�o �o�o);M_ q������� ��%�7�I�[�m���������Ǐُ� � H552���21�R78��50�J614��ATUP7�54�57�6�VCAM��CRI��UIFv7�28��NRE��52v�R63�S�CH�LICƚDwOCV�CSU��8697�0F�EI�OCǛ4�R69�v�ESETW�u�J�7u�R68�MA{SK�PRXY��]7�OCO��3W�h���6�3�J65��536�H$�LCH^ƪOPLGW�0��MHCRǪS��MkCSV�0��55F��MDSW���OP���MPR���6�0n6�PCM��R0E˰��F���6�51f�5u1��0f�PRS���69�FRD��FwREQ�MCN�{936�SNBAכ^%�SHLB�ME�t�ּ26�HTCV��TMIL�6�TP�AV�TPTX��ELړ�6�8%�#��wJ95��TUT���95�UEV��U�ECƪUFR��V�CCf�O��VIP��CSC��CSGtƚ$�I�WEBV�7HTTV�R6՜��lS���CG��IG��oIPGS'�RC���DG��H7��R6�6f�5�u�R��R�51f�6�2�5�v�#�J׼��6��L�U�5�s�v�4��66�F�R64�NVDv��R6��R84�k79�4��S5嫷J76�D0uFnRTS&�CR�wCRX��CLI&̎e�CMSV�sV�S�TY��6�CTOhV�#�V�75�NN��ORS����6�FC�BV�FCF��CH�V�FCR��FCI�F�FC��J#��G�
M��OL�EN�DǪLU��CPR���Lu�S�C$�SvtTE�S60��FVRV�IN��IH���m??�?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� ������������ '9K]o��� �����#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s����������͏ߏ��STD�LANG���0�B� T�f�x���������ҟ �����,�>�P�b� t���������ί�� ��(�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢ� ����������� �2� D�V�h�zߌߞ߰����RBT
�OPTN ������'�9�K�]� o�����������DPN	���)�;� M�_�q����������� ����%7I[ m������ ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ� ����������'�9� K�]�o߁ߓߥ߷��� �������#�5�G�Y� k�}���������� ����1�C�U�g�y� ��������������	 -?Qc�f�������99���$FEAT_�ADD ?	����  	�#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙπ�Ͻ��������D�EMO y   �L�B� T߁�xߊ߷߮����� ������G�>�P�}� t����������� ��C�:�L�y�p��� ������������ ?6Hul~�� ����;2 Dqhz���� �� /
/7/./@/m/ d/v/�/�/�/�/�/�/ �/?3?*?<?i?`?r? �?�?�?�?�?�?�?O /O&O8OeO\OnO�O�O �O�O�O�O�O�O+_"_ 4_a_X_j_�_�_�_�_ �_�_�_�_'oo0o]o Tofo�o�o�o�o�o�o �o�o#,YPb �������� ��(�U�L�^����� ������ʏ���� $�Q�H�Z���~����� ��Ɵ����� �M� D�V���z�������¯ ܯ��
��I�@�R� �v���������ؿ� ���E�<�N�{�r� �ϱϨϺ������� �A�8�J�w�n߀߭� �߶���������=� 4�F�s�j�|���� ��������9�0�B� o�f�x����������� ����5,>kb t������� 1(:g^p� ������ /-/ $/6/c/Z/l/�/�/�/ �/�/�/�/�/)? ?2? _?V?h?�?�?�?�?�? �?�?�?%OO.O[ORO dO�O�O�O�O�O�O�O �O!__*_W_N_`_�_ �_�_�_�_�_�_�_o o&oSoJo\o�o�o�o �o�o�o�o�o" OFX�|��� ������K�B� T���x�������ۏҏ ����G�>�P�}� t�������ןΟ��� ��C�:�L�y�p��� ����ӯʯܯ	� �� ?�6�H�u�l�~����� Ͽƿؿ����;�2� D�q�h�zϔϞ����� �����
�7�.�@�m� d�vߐߚ��߾����� ���3�*�<�i�`�r� ������������� /�&�8�e�\�n����� ������������+" 4aXj���� ����'0] Tf������ ��#//,/Y/P/b/ |/�/�/�/�/�/�/�/ ??(?U?L?^?x?�? �?�?�?�?�?�?OO $OQOHOZOtO~O�O�O �O�O�O�O__ _M_ D_V_p_z_�_�_�_�_ �_�_o
ooIo@oRo lovo�o�o�o�o�o�o E<Nhr �������� �A�8�J�d�n����� ��яȏڏ����=� 4�F�`�j�������͟ ğ֟����9�0�B� \�f�������ɯ��ү �����5�,�>�X�b� ������ſ��ο��� �1�(�:�T�^ϋς� ���ϸ������� �-� $�6�P�Z߇�~ߐ߽� ����������)� �2� L�V��z������ ������%��.�H�R� �v������������� ��!*DN{r ������� &@Jwn�� �����//"/ </F/s/j/|/�/�/�/ �/�/�/???8?B? o?f?x?�?�?�?�?�? �?OOO4O>OkObO tO�O�O�O�O�O�O_|_0]  'X F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ����������
��.�  /�)�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o�o "4FXj|�� �������0� B�T�f�x��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@� R�d�v߈ߚ߬߾��� ������*�<�N�`� r����������� ��&�8�J�\�n��� �������������� "4FXj|�� �����0 BTfx���� ���//,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�?�? O O$O6OHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Rodovo�o�o�o�o�o �o�o*<N` r������� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P� b�t���������ο� ���(�:�L�^�p� �ϔϦϸ������� �(�$�4�8�+�N� `�r߄ߖߨߺ����� ����&�8�J�\�n� ������������� �"�4�F�X�j�|��� ������������ 0BTfx��� ����,> Pbt����� ��//(/:/L/^/ p/�/�/�/�/�/�/�/  ??$?6?H?Z?l?~? �?�?�?�?�?�?�?O  O2ODOVOhOzO�O�O �O�O�O�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ� ����������
��.� @�R�d�v����� ��������*�<�N� `�r������������� ��&8J\n �������� "4FXj|� ������// 0/B/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?t?�?�?�?�?�? �?�?OO(O:OLO^O pO�O�O�O�O�O�O�O� __$_6Y�$FE�AT_DEMOIoN  ;T�fP��<PNTINDE�X[[jQ�NPIL�ECOMP z�����Q�iRIU�PSETUPo2 {�U�R?�  N �Q�S�_AP2BCK �1|�Y  �)7Xok%�_8o<P�P&oco9U�_�oo �oBo�o�oxo�o1 C�og�o��,� P�����?�� L�u����(���Ϗ^� 󏂏�)���M�܏q� �����6�˟Z�؟� ��%���I�[���� ����D�ٯh������ 3�¯W��d������ @�տ�v�Ϛ�/�A� пe����ϛ�*Ͽ�N� ��r���ߨ�=���a� s�ߗ�&߻���\��� ���'��K���o��� |��4���X������ #���G�Y���}���� ��B���f�����1t�Y�PP�_ 2�P*.VR8���*��������l PC���F'R6:�2�V�TzPz�w��]PG���*.F�o/��	�:,8�^/�STMi/�/ /�-M/�/�H�/?�'?�/�/g?�GIFq?�?�%�?pD?V?�?�JPG�?�O�%O�?�?oO�
JSyO�O��5C�OMO�%
JavaSc�ript�O�?CS�O&_�&_�O %�Cascadin�g Style ?SheetsR_���
ARGNAME�.DT�_��� \@�_S_�A�T�_�_�P�DISP*�_����To�_�QLaZooCLLB.ZIwo,2o$ :\�a\�o�i��ACollab�o�o�o
TPEI?NS.XML�_�:\![o�QCus�tom Tool�barbiPAS�SWORDQo��FRS:\�dB`�Password Config� ��/��(�e���� ����N��r����� =�̏a������&��� J���񟀟���9�K� ڟo�������4�ɯX� �|���#���G�֯@� }����0�ſ׿f��� ���1���U��y�� ϯ�>���b���	ߘ� -߼�Q�c��χ�߫� ��L���p��ߦ�;� ��_���X��$��H� ����~����7�I��� m���� �2���V��� z���!��E��i{ 
�.��d�� ��S�wp �<�`�/�+/ �O/a/��//�/8/ J/�/n/?�/�/9?�/ ]?�/�?�?"?�?F?�? �?|?O�?5O�?�?kO �?�OO�O�OTO�OxO __�OC_�Og_y__ �_,_�_P_b_�_�_o �_oQo�_uoo�o�o :o�o^o�o�o)�o M�o�o��6� �l��%�7��[� ���� ���D�ُh� z����3�,�i��� �����ßR��v�������$FILE�_DGBCK 1�|������ < ��)
SUMMAR�Y.DG!�͜M�D:U���ِD�iag Summ�ary����
CONSLOG��n����ٯ���Console log����	TPACCN��t�%\�����T�P Accoun�tin;���FR�6:IPKDMPO.ZIPͿј
��ϥ���Excep�tion"�ӻ��MEMCHECK���������-�Mem�ory Data|����Jn )��RIPE�~ϐ�%���%�� Pa?cket L:����L�$�c���ST�AT��߭� �%A�Stat�us��^�	FTP�����	��/�m�ment TBD�2�^� >I)E?THERNEw�
��d�u�﨡Eth�ernJ�1�fig�uraAϩ��DCSVRF&���7������ veri?fy all:���� 4��DIF�F/��'���;�Q�d�iff��r�d���CHG01������A�����it�2���2 70���fx�3���I ��p�VTRNDIAG.LSu�&8���� O�pe��L� ��no�stic��lϿ)VDEV�D�AT�������Vis�Devisce�+IMG���,/>/�/:�i$I�magu/+UP� ES/�/FR�S:\?Z=��U�pdates L�istZ?��� FLEXEVEN��в/�/�?���1 UIF EvM�M����-vZ)CR?SENSPK�/˞��\!O���CR�_TAOR_PEA�KbOͩPSRBW�LD.CM�O͜�E2�O\?.�PS_R?OBOWELS���:GIG��@_�?d_>��GigE�(O~��N�@�)UQHADOW__D_V_��_��Shado�w Change�����Edt�RRCMERR�_�_�_oo���4`CFG E�rroro tai}lo MA�k�CMSGLIBgo�No`o�o|R�e��z0iyc�o�a�)�`�ZD0_O�os���ZD�Pad�l= �RNOTI�R�d���Noti�fic����,�AG��P�ӟt����� ����Ώ]�����(� ��L�^�폂������ G�ܟk� ����6�ş Z��~������C�د �y����2�D�ӯh� �������¿Q��u� 
�ϫ�@�Ͽd�v�� ��)Ͼ���_��σ�� ��%�N���r�ߖߨ� 7���[�����&�� J�\��߀���3�� ��i����"�4���X� ��|������A����� w���0��=f�� ���O�s �>�bt� '�K���/� :/L/�p/��/�/5/ �/Y/�/ ?�/$?�/H? �/U?~??�?1?�?�? g?�?�? O2O�?VO�? zO�OO�O?O�OcO�O 
_�O._�OR_d_�O�_ _�_�_M_�_q_oo �_<o�_`o�_mo�o%o �oIo�o�oo�o8 J�on�o��3� W�{�"��F�� j�|����/�ď֏e�������0��$FI�LE_FRSPRT  ������?��MDONLY 1�|S�� 
 ��)MD:_V�DAEXTP.Z�ZZ1�⏹�ț�6%NO Ba�ck file <���S�6P��� ��>��K�t�����'� ��ί]�򯁯�(��� L�ۯp������5�ʿ Y�׿ Ϗ�$ϳ�H�Z� �~�Ϣϴ�C���g� ��ߝ�2���V���c� ��߰�?�����u�
� ��.�@���d��߈��~C�VISBCKq�|[���*.VD��|��S�FR:\���ION\DATA�\��v�S�Vision VD� ��Y�k����y�� B�����x���1C ��g���,�P ����?�P u�(��^� �/��M/�q/�/ >/�/6/�/Z/�/?�/ %?�/I?[?�/??�?�2?D?�?9�LUI_�CONFIG �}S����; '$ �3v�{S�;O�MO_OqO�O�O�I#@|x�?�O�O�O__%\ �OH_Z_l_~_�_'_�_ �_�_�_�_o�_2oDo Vohozo�o#o�o�o�o �o�o
�o.@Rd v������ ��*�<�N�`�r��� �����̏ޏ����� &�8�J�\�n������ ��ȟڟ쟃���"�4� F�X�j��������į ֯����0�B�T� f�����������ҿ� {���,�>�P�b��� �ϘϪϼ�����w�� �(�:�L�^��ςߔ� �߸�����s� ��$� 6�H���Y�~���� ��]������ �2�D� ��h�z���������Y� ����
.@��d v����U�� *<�`r� ���Q��// &/8/�\/n/�/�/�/ ;/�/�/�/�/?"?�/ F?X?j?|?�?�?7?�? �?�?�?OO�?BOTO fOxO�O�O3O�O�O�O �O__�O>_P_b_t_ �_�_/_�_�_�_�_o o�_:oLo^opo�o�o>$h  x�o�c��$FLUI_D�ATA ~�����a�(a�dRESULT� 3�ep ��T�/wi�zard/gui�ded/step�s/Expert �o=Oas��������z�C�ontinue �with Gpance�:�L�^�p� ��������ʏ܏� �� �b-�a�e�0 �0`��c�a6?��ps��� ������ҟ����� ,�>�P��0ow����� ����ѯ�����+��=�O�a�?�1�C�U�e�cllbs�ֿ� ����0�B�T�f�x� �Ϝ�[���������� �,�>�P�b�t߆ߘ�@��i�{��ߟ�]�e�rip(pſ-�?�Q� c�u��������� ����)�;�M�_�q� �������������� ������`�e�#p�TimeUS/DST	��������!3E�Enabl(�y� ������	//(-/?/Q/�b�)0�/M_q24|�/ �/??)?;?M?_?q? �?�?Tf�?�?�?O O%O7OIO[OmOO�O �Ob/t/�/�/Z�"q?Region�O5_ G_Y_k_}_�_�_�_�_��_�_�America!�#o5oGoYo ko}o�o�o�o�o�o�o��Ay�O�O3�O_~qEditor�o ����������+�=� � Tou�ch Panel� rs (reco/mmenp�)K��� ����Ə؏���� �2�D�|�%��I|[qacceso ܟ� ��$�6�H�Z��l�~�����Con�nect to Network�� ֯�����0�B�T��f�x�����x��@���}����,!��s I�ntroduct !_4�F�X�j�|ώϠ� �����������0� B�T�f�xߊߜ߮��������� ɿ� �"�i�{���� ����������/�A�  �e�w����������������+=�H�3��+�O� ���� 2D Vhz�K���� ��
//./@/R/d/ v/�/�/Yk}�/� ??*?<?N?`?r?�? �?�?�?�?�?��?O &O8OJO\OnO�O�O�O �O�O�O�O�/_�/1_ �/X_j_|_�_�_�_�_ �_�_�_oo0oBoS_ foxo�o�o�o�o�o�o �o,>�O_!_ �E_������ �(�:�L�^�p����� So��ʏ܏� ��$� 6�H�Z�l�~���O�� s՟���� �2�D� V�h�z�������¯ԯ 毥�
��.�@�R�d� v���������п⿡� �ş'�9���`�rτ� �ϨϺ��������� &�8���\�n߀ߒߤ� �����������"�4� �=��a��Mϲ��� ��������0�B�T� f�x���I߮������� ��,>Pbt �E��i���� (:L^p�� ������ //$/ 6/H/Z/l/~/�/�/�/ �/�/����/?� V?h?z?�?�?�?�?�? �?�?
OO.O�ROdO vO�O�O�O�O�O�O�O __*_<_�/??�_ C?�_�_�_�_�_oo &o8oJo\ono�o?O�o �o�o�o�o�o"4 FXj|�M___q_ ��_���0�B�T� f�x���������ҏ�o ���,�>�P�b�t� ��������Ο���� �%��L�^�p����� ����ʯܯ� ��$� 6�G�Z�l�~������� ƿؿ���� �2�� S��w�9��ϰ����� ����
��.�@�R�d� v߈�G��߾������� ��*�<�N�`�r�� Cϥ�g���ύ��� &�8�J�\�n������� ����������"4 FXj|���� ������-��T fx������ �//,/��P/b/t/ �/�/�/�/�/�/�/? ?(?�1U??A �?�?�?�?�? OO$O 6OHOZOlO~O=/�O�O �O�O�O�O_ _2_D_ V_h_z_9?�?]?�_�_ �?�_
oo.o@oRodo vo�o�o�o�o�o�O�o *<N`r� �����_�_�_�_ #��_J�\�n������� ��ȏڏ����"��o F�X�j�|�������ğ ֟�����0��� �u�7�������ү� ����,�>�P�b�t� 3�������ο��� �(�:�L�^�pς�A� S�e��ω��� ��$� 6�H�Z�l�~ߐߢߴ� �߅������ �2�D� V�h�z�������� ��������@�R�d� v��������������� *;�N`r� ������ &��G	�k-��� �����/"/4/ F/X/j/|/;�/�/�/ �/�/�/??0?B?T? f?x?7�?[�?�? �?OO,O>OPObOtO �O�O�O�O�O�/�O_ _(_:_L_^_p_�_�_ �_�_�_�?�_�?o!o �OHoZolo~o�o�o�o �o�o�o�o �OD Vhz����� ��
���_%o�_I� s�5o������Џ�� ��*�<�N�`�r�1 ������̟ޟ��� &�8�J�\�n�-�w�Q� ��ů������"�4� F�X�j�|�������Ŀ �������0�B�T� f�xϊϜϮ������ �����ٯ>�P�b�t� �ߘߪ߼�������� �տ:�L�^�p��� ��������� ��$� �����i�+ߐ����� �������� 2D Vh'����� ��
.@Rd v5�G�Y��}��� //*/</N/`/r/�/ �/�/�/y�/�/?? &?8?J?\?n?�?�?�? �?�?��?�O�4O FOXOjO|O�O�O�O�O �O�O�O__/OB_T_ f_x_�_�_�_�_�_�_ �_oo�?;o�?_o!O �o�o�o�o�o�o�o (:L^p/_� ����� ��$� 6�H�Z�l�+o��Oo�� sou����� �2�D� V�h�z�������� ���
��.�@�R�d� v���������}�߯�� ��ٟ<�N�`�r��� ������̿޿��� ӟ8�J�\�nπϒϤ� �����������ϯ� �=�g�)��ߠ߲��� ��������0�B�T� f�%ϊ��������� ����,�>�P�b�!� k�Eߏ���{����� (:L^p�� ��w��� $ 6HZl~��� s�������/��2/D/ V/h/z/�/�/�/�/�/ �/�/
?�.?@?R?d? v?�?�?�?�?�?�?�? OO���]O/�O �O�O�O�O�O�O__ &_8_J_\_?�_�_�_ �_�_�_�_�_o"o4o FoXojo)O;OMO�oqO �o�o�o0BT fx���m_�� ���,�>�P�b�t� ��������{oݏ�o� �o(�:�L�^�p����� ����ʟܟ� ��#� 6�H�Z�l�~������� Ưد����͏/�� S��z�������¿Կ ���
��.�@�R�d� #��ϚϬϾ������� ��*�<�N�`���� C���g�i������� &�8�J�\�n���� ��u��������"�4� F�X�j�|�������q� ������	��0BT fx������ ���,>Pbt �������/ ����1/[/�/�/ �/�/�/�/�/ ??$? 6?H?Z?~?�?�?�? �?�?�?�?O O2ODO VO/_/9/�O�Oo/�O �O�O
__._@_R_d_ v_�_�_�_k?�_�_�_ oo*o<oNo`oro�o �o�ogOyO�O�O�o�O &8J\n��� ������_"�4� F�X�j�|�������ď ֏�����o�o�oQ� x���������ҟ� ����,�>�P��t� ��������ί��� �(�:�L�^��/�A� ��e�ʿܿ� ��$� 6�H�Z�l�~ϐϢ�a� ��������� �2�D� V�h�zߌߞ߰�o��� ���߷��.�@�R�d� v����������� ��*�<�N�`�r��� �������������� #��G	�n��� �����"4 FX�|���� ���//0/B/T/ u/7�/[]/�/�/ �/??,?>?P?b?t? �?�?�?i�?�?�?O O(O:OLO^OpO�O�O �Oe/�O�/�O�O�?$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_�? o2oDo Vohozo�o�o�o�o�o �o�o�O_�O%O_ v������� ��*�<�N�or��� ������̏ޏ���� &�8�J�	S-w��� cȟڟ����"�4� F�X�j�|�����_�į ֯�����0�B�T� f�x�����[�m���� 󿵟�,�>�P�b�t� �ϘϪϼ������ϱ� �(�:�L�^�p߂ߔ� �߸������� ￿ѿ �E��l�~���� ��������� �2�D� �h�z����������� ����
.@R� #�5�Y���� *<N`r� �U�����// &/8/J/\/n/�/�/�/ c�/��/�?"?4? F?X?j?|?�?�?�?�? �?�?�??O0OBOTO fOxO�O�O�O�O�O�O �O�/_�/;_�/b_t_ �_�_�_�_�_�_�_o o(o:oLoOpo�o�o �o�o�o�o�o $ 6H_i+_�O_Q ����� �2�D� V�h�z�����]oԏ ���
��.�@�R�d� v�����Y��}ߟ� ���*�<�N�`�r��� ������̯ޯ𯯏� &�8�J�\�n������� ��ȿڿ쿫���ϟ� C��j�|ώϠϲ��� ��������0�B�� f�xߊߜ߮������� ����,�>���G�!� k��Wϼ�������� �(�:�L�^�p����� S߸������� $ 6HZl~�O�a� s����� 2D Vhz����� ���
//./@/R/d/ v/�/�/�/�/�/�/�/ ���9?�`?r?�? �?�?�?�?�?�?OO &O8O�\OnO�O�O�O �O�O�O�O�O_"_4_ F_??)?�_M?�_�_ �_�_�_oo0oBoTo foxo�oIO�o�o�o�o �o,>Pbt ��W_�{_��_� �(�:�L�^�p����� ����ʏ܏���$� 6�H�Z�l�~������� Ɵ؟꟩��/�� V�h�z�������¯ԯ ���
��.�@���d� v���������п��� ��*�<���]���� C�EϺ��������� &�8�J�\�n߀ߒ�Q� �����������"�4� F�X�j�|��Mϯ�q� �������0�B�T� f�x������������� ��,>Pbt ���������� ��7��^p�� ����� //$/ 6/��Z/l/~/�/�/�/ �/�/�/�/? ?2?� ;_?�?K�?�?�? �?�?
OO.O@OROdO vO�OG/�O�O�O�O�O __*_<_N_`_r_�_ C?U?g?y?�_�?oo &o8oJo\ono�o�o�o �o�o�o�O�o"4 FXj|���� ���_�_�_-��_T� f�x���������ҏ� ����,��oP�b�t� ��������Ο���� �(�:�����A� ����ʯܯ� ��$� 6�H�Z�l�~�=����� ƿؿ���� �2�D� V�h�zό�K���o��� ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�� ������������� #���J�\�n������� ����������"4 ��Xj|���� ���0��Q �u7�9���� �//,/>/P/b/t/ �/E�/�/�/�/�/? ?(?:?L?^?p?�?A �?e�?�?�/ OO$O 6OHOZOlO~O�O�O�O �O�O�/�O_ _2_D_ V_h_z_�_�_�_�_�_ �?�?�?o+o�?Rodo vo�o�o�o�o�o�o�o *�ON`r� �������� &��_/o	oS�}�?o�� ��ȏڏ����"�4� F�X�j�|�;����ğ ֟�����0�B�T� f�x�7�I�[�m�ϯ�� ����,�>�P�b�t� ��������ο���� �(�:�L�^�pςϔ� �ϸ����ϛ�����!� �H�Z�l�~ߐߢߴ� ��������� �߿D� V�h�z�������� ����
��.������ s�5ߚ����������� *<N`r1� ������ &8J\n�?�� c������/"/4/ F/X/j/|/�/�/�/�/ �/��/??0?B?T? f?x?�?�?�?�?�?� �?�O�>OPObOtO �O�O�O�O�O�O�O_ _(_�/L_^_p_�_�_ �_�_�_�_�_ oo$o �?EoOio+O-o�o�o �o�o�o�o 2D Vhz9_���� ��
��.�@�R�d� v�5o��Yo��͏�� ��*�<�N�`�r��� ������̟���� &�8�J�\�n������� ��ȯ��я������ F�X�j�|�������Ŀ ֿ�����ݟB�T� f�xϊϜϮ������� ����ٯ#���G�q� 3��ߪ߼�������� �(�:�L�^�p�/ϔ� ��������� ��$� 6�H�Z�l�+�=�O�a� �������� 2D Vhz������ ��
.@Rd v��������� ��/��</N/`/r/�/ �/�/�/�/�/�/?? �8?J?\?n?�?�?�? �?�?�?�?�?O"O� �/gO)/�O�O�O�O �O�O�O__0_B_T_ f_%?w_�_�_�_�_�_ �_oo,o>oPoboto 3O�oWO�o{O�o�o (:L^p�� ����o� ��$� 6�H�Z�l�~������� Ə�o珩o��o2�D� V�h�z�������ԟ ���
���@�R�d� v���������Я��� ��׏9���]��!� ������̿޿��� &�8�J�\�n�-��Ϥ� �����������"�4� F�X�j�)���M����� ��������0�B�T� f�x��������� ����,�>�P�b�t� ��������{��ߟ��� ��:L^p�� ����� �� 6HZl~��� ����/���� ;/e/'�/�/�/�/�/ �/�/
??.?@?R?d? #�?�?�?�?�?�?�? OO*O<ONO`O/1/ C/U/�Oy/�O�O__ &_8_J_\_n_�_�_�_ �_u?�_�_�_o"o4o FoXojo|o�o�o�o�o �O�O�O	�O0BT fx������ ���_,�>�P�b�t� ��������Ώ���� ��o�o�o[����� ����ʟܟ� ��$� 6�H�Z��k������� Ưد���� �2�D� V�h�'���K���o�Կ ���
��.�@�R�d� vψϚϬϾ�Ͽ���� ��*�<�N�`�r߄� �ߨߺ�y��ߝ����� &�8�J�\�n���� �������������4� F�X�j�|��������� ��������-��Q ������� �,>Pb!� �������/ /(/:/L/^//A �/�/y�/�/ ??$? 6?H?Z?l?~?�?�?�? s�?�?�?O O2ODO VOhOzO�O�O�Oo/�/ �/�O_�/._@_R_d_ v_�_�_�_�_�_�_�_ o�?*o<oNo`oro�o �o�o�o�o�o�o�O _�O/Y_��� ������"�4� F�X�o|�������ď ֏�����0�B�T� %7I��mҟ� ����,�>�P�b�t� ������i�ί��� �(�:�L�^�p����� ����w���������$� 6�H�Z�l�~ϐϢϴ� �������ϻ� �2�D� V�h�zߌߞ߰����� ����
�ɿۿ�O�� v����������� ��*�<�N��_��� ������������ &8J\�}?� c�����"4 FXj|���� ���//0/B/T/ f/x/�/�/�/m�/� �/�?,?>?P?b?t? �?�?�?�?�?�?�?O �(O:OLO^OpO�O�O �O�O�O�O�O _�/!_ �/E_?	_~_�_�_�_ �_�_�_�_o o2oDo VoOzo�o�o�o�o�o �o�o
.@R_ s5_��mo��� ��*�<�N�`�r��� ����gȍޏ���� &�8�J�\�n������� c��џ���"�4� F�X�j�|�������į ֯������0�B�T� f�x���������ҿ� ������ٟ#�M��t� �ϘϪϼ�������� �(�:�L��p߂ߔ� �߸������� ��$� 6�H���+�=ϟ�a� ��������� �2�D� V�h�z�����]����� ����
.@Rd v���k�}������$FMR2_�GRP 1���� ��C4  B��	� ��9K6F�@ a@�6G��  �Fg�f�C�8R�y?��  ��66�X����875t���5���5`+=�yA�  /+�BH�w-%@S3	39%�5[/l-6@6!�/xl/�/�/�/ �/?�/&??J?5?G?��?k?�?��_CF/G �TK�?��? OO�9NO �
F0FA �K@�<RM_CHK?TYP  ��p$&� ROMa@�_MINg@������@�R XSS�B�3�� 7�O���C�O��O�5TP_DEF�_OW  ��|$WIRCOMf@�_�$GENOV_RD_DO�F��fE]TH��D dbU�dKT_ENB7_ �KPRAVC�:�G�@ �Y�O�_�?oyo&oI*� �QOU��NAIRI<�@��oGo�o�o,�o��C�p3�P�O:��B�+spL�i�O�PSMTኹY(�@
t�$HoOSTC�21�ε@�5 M5C��R{���  27.00�=1�  e�]� o�������K�ď֏���������	ano?nymous!�O�a�s����� �4��������D�!�3� E�W�i���������ï 柀�.���/�A�S� ��课�П����Ŀ ����+�r�O�a�s� �ϗϺ�������� �'�n��������ϓ� ڿ����������F�#� 5�G�Y�k���υ�� ��������B�T�f�C� z�g��ߋ�������� ����	-P����� u������(� :�<)p�M_q� �������/$ ZlI/[/m//�/� ���//�/D!?3? E?W?/?�?�?�?�? �/�?./OO/OAOSO �/�/�/�/�?�O?�O �O__+_r?O_a_s_ �_�_�O�?O�_�_o�o'o�t�qENT {1�hk P!�_.no  �p\o�o �o�o�o�o�o�o �o:_"�F�j �����%��I� �m�0���T�f�Ǐ�� 돮��ҏ3���,�i� X���P���t�՟��� ��
�/��S��w�:� ��^�������������ܯ=� �QUIC�C0J�&�!19�2.168.1.10c�X�1��v�8���\�2�ƿؿ9�!ROUTER:���!��a��P�CJOG��e�!�* ��0��U�C�AMPRT�϶�!1�����RTS����x� !Sof�tware Op�erator PanelU߇���7kNAME !Kj?!ROBO�����S_CFG 1��Ki ��Auto-sta�rted�DFTP�Oa�O�_���O ����������E_�.� @�R�u�c�	������� ����cN:�L�^�;r� ��R������� �%H�[m ���jO|O�O�O 4!/hE/W/i/{/�/ T�/�/�/�/�//�/ /?A?S?e?w?�?�� ��??�?</O+O=O OO?sO�O�O�O�O�? `O�O__'_9_K_�? �?�?�?�O�_�?�_�_ �_o#o�OGoYoko}o �o�_4o�o�o�o�o f_x_�_g�o��_ �����o��-� ?�Q�tu�������� Ϗ�(:L^`�2� �q�����������ݟ ���%�H�ʟ[�m� ���������� �ί 4�!�h�E�W�i�{��� T���ÿտ�
�Ϟ��/�A�S�e�w����_?ERR ��ڇ����PDUSIZ � �^6�����>��WRD ?�(����  ?guest����+�=�O�a���SC�D_GROUP [3�(� ,�"�wIFT��$PA��wOMP�� �޷_SH��ED�� �$C��COM��T�TP_AUTH �1��� <!iPendanm��x�#�+!KAR�EL:*x����KC������V�ISION SET��(����?�-�W�R���v������������������G�CTR/L ���a��
�FFF9�E3��FRS�:DEFAULT��FANUC� Web Server�
tdG��� �/� 2DV���WR_CONF�IG ���������IDL_CPU_PC� ��B���� BH�MIN����?GNR_IO�������ȰHMI_E�DIT ���
 ($/C/��2/k/ V/�/z/�/�/�/�/�/ ?�/1??U?@?y?d? �?�?./�?�?�?�?O O?OQO<OuO`O�O�O �O�O�O�O�O__;_��NPT_SIM�_DO�*NS�TAL_SCRN�� �\UQTPM?ODNTOL�Wl[�RTYbX�qV�.K�ENB�W�ӭOLNK 1�����o%o7oIo[omo|o�RMASTE���Y%OSLAV�E ��ϮeRA?MCACHE�o�R}OM�O_CFG�o��S�cUO'��bCMT_OP�  "�ʎ5sYCL�ou� _?ASG 1����
 �o���� ���"�4�F�X�j�p|����kwrNUM��5��
�bIP�o�gRTRY_CN@<uQ_UPD��a���� �bp�b���n��M��аP}T?=��k ��._�� ����ɟ۟퟈S��� )�;�M�_�q� ����� ��˯ݯ�~��%�7� I�[�m��������ǿ ٿ�����!�3�E�W� i�{�
ϟϱ������� �ψϚ�/�A�S�e�w� ��߭߿�������� ��+�=�O�a�s��� &������������ 9�K�]�o�����"��� ������������G Yk}��0�� ���CUg y��,>��� 	//-/�Q/c/u/�/ �/�/:/�/�/�/?? )?�/�/_?q?�?�?�? �?H?�?�?OO%O7O �?[OmOO�O�O�ODO VO�O�O_!_3_E_�O i_{_�_�_�_�_R_�_ �_oo/oAo�_�_wo �o�o�o�o�o`o�o +=O�os�� ���\n��'� 9�K�]�����������ɏۏi�c�_MEMBERS 2�:��   u$:� ���v����1���RCA_�ACC 2���   �[~�� T��  � 5�Я 5�`l�l��l��1� (1_������  l����a�BUF001 �2�n�= �n�u0  u0�{������������������J�����T�R��u0Hq�U$R�1R�=R�K���-�  �S�<����X��g���u��������� �@Ȑ@�'��4�ڤBڤOڤ\ڤk�ڤw�� 6H ���
�
�٤�VᤘC
�P
�]
�Ul
�x
��
��
�U�
��
��
��
�VA���
����U��+�8��F�S�b�ߙ2�����u0#�Qx(��0�5�9�5�A��5�I�H�,�P�s�(X�q �`�,�HHp�p�i�x�u0L )���@ H��B�3��j�
h��h�������0������ɠt��Ѡ ҡد���� �2�D� V�h�z�������¿Կ�3���7��7�� 7��7�!�7�)�7���9�G��I�7�Q�   X�h�a�h�i�f�q�h� ��h���h��������� �����婢�����Þ� ���Þ�Ѣ�������� �����������
����  � �"� �*�  ���9� �B� �J� � R� �Z� �b� �j� � r� �z� ��� ��� � �� �S�� ��7��� 7���7���7���7��� 7���7���7�����d��CFG 2�n�� 4��l�l�<�l�47��HIuS钜n� ��� 2025-1�1-3�l� �   # &�f  ' "8珪�  Pl�7 �X���6hl��p�l�$  x {�8w �l�;  ��� 7 ����9 ��  :��7[}�Rq29}	7v����������   % � � � -�R  I*� l��B��a N/`/r/�/�/�/�/�/ �/�/'/9/&?8?J?\? n?�?�?�?�?�?�/? �?O"O4OFOXOjO|O �O�O�?�?�O�O�O_ _0_B_T_f_x_�O�O �O�_�_�_�_oo,o >oPo�O��[m
8 c� 8���o�o�6d� �b���b�� +  X�  2X�  d!qc��,: J!r_0  Q��0p�o;M_���@�����$:�a� 2�a ,*q 1  \�_�_m�� ������Ǐُ���� �_X�E�W�i�{����� ��ß՟��0���/� A�S�e�w��������� ������+�=�O� a�s���������߿ ���'�9�K�]�o�@��J�Ѐo�o

eq� ��������� @��� ��p��� eq� Geq	$"6pMr��po�]o ������������#�5���� �� Z�  �־�п������ ������&�8�o�� n��������������� ��G�Y�FXj| ������1 �0BTfx�� ���	//,/ >/P/b/t/�/�/�Ϙ��I_CFG 2���� H
Cy�cle Time��Busy��Idl�"�mi�n�+1Up|�&�Read�'Dow8?�`� 1�#Count>�	Num �"�����<��b�qaP�ROG�"�������)/sof�tpart/ge�nlink?cu�rrent=me�nupage,1133,1�/OO�/OAO3b5leSDT�_ISOLC  ����p�/J2�3_DSP_EN�BL�vK0�@INCG ��M�ӄ@An��?&p=���<#��
�A�I:�o����N_���O<_�GOB�0C�CF�1�FVQ�G_GROUP �1�vK	r<A��C�٢_D_?���?�_��Q�_o.o�@o�_dovo�o�o���,_NYG_IN_A�UTODԫMPOS�RE^_pVKANJ?I_MASK v�H�qRELMON #��˔?��y_ox������.6r�3��7�C���u�o�D�KCL_L�`NU�ML��EYLOGOGINGDЫ���Q��E�0LANGUA_GE ��~���DEFAUgLT ����LG�!���:2�?��W�80H  ����'��  � 
ɾgҊ�GOUF ;���
��(UTg1:\��  � -�?�Q�h�u������� ��ϟ�����(g4��8i�N_DISP ��O8�_�_��?LOCTOL�����Dz`�A�A��GB�OOK ���d �1
�
�۠#�� ���#�5�G�Y�i���3{�W�	��쉞Q�QJ¿Կ1��_B�UFF 2�vK ���25
�ڢ�VB&�7 Col�laborativ�=�OΗώϠϲ� ��������'��0�]��T�fߓߊߜ��DCS ��9�B�Ax� ��Rh�%�-�?�Q����IO 2��� 1���Q��� �����������*� <�N�b�r��������� ������&:e�ER_ITMsNd �o������� #5GYk}� ��������h�SEV�`�MdTYPsN�c/u/�/�
-�aRST5���S�CRN_FL 2�s��0����/?�?1?C?U?g?�/TP�K�sOR"��NGN�AM�D��~�N�UPS_ACR� �4�DIGI�8+)U�_LOAD[PG �%�:%T_N�OVICEt?��MAXUALRM2�,�a���E
ZB�1_P�5�` ��y�Z@CY��˭�O+���xۡ�D|PP 2�˫ �Uf	R/_
_ C_._g_y_\_�_�_�_ �_�_�_�_oo?oQo 4ouo`o�o|o�o�o�o �o�o)M8q Tf������ �%��I�,�>��j� ����Ǐُ�����!� ��W�B�{�f����� ��՟����ܟ�/�� S�>�w���l�����ѯ ��Ư��+��O�a��D���p���RHDBG?DEF ��E����O��_LDXDI�SA�0�;c�MEM�O_AP�0E ?=�;
 ױ�� 3�E�W�i�{ύϟϱ��Z@FRQ_CFG� ��G۳A ���@��Ô�<��dA%�� ������B��K���*zi�/k� **:t� ��g�y�ߔ��߱��� �������J�E�s�J d�����,(H���[�����@� '�Q�v�]��������� ������*NPJ?ISC 1��9Z� ������ܿ������	Zl_MS�TR �#-,S_CD 1�"͠ {������� �//A/,/e/P/�/ t/�/�/�/�/�/?�/ +??O?:?L?�?p?�? �?�?�?�?�?O'OO KO6OoOZO�O~O�O�O �O�O�O_�O5_ _Y_ D_i_�_z_�_�_�_�_ �_�_o
ooUo@oyo do�o�o�o�o�o�o�o ?*cN�MK���;љ$MLTARM����N��r ��հ��İMETsPU��zr��C�NDSP_ADC�OL%�ٰ0�CMNmTF� 9�FNb�|f�7�FSTLI��x�4 �;ڎ�s�����9�POSC�F��q�PRPMle��STD�1�;w 4�#�
v� �qv�����r������� �̟ޟ ���V�8� J���n���¯��������9�SING_C�HK  ��$M7ODA���t�{��~2�DEV 	��	MC:f�HOSIZE��zp�2�TASK %��%$123456�789 ӿ�0�T�RIG 1�; lĵ�2ϻ�!�bό��YP����H��1�EM_INF �1�N�`)�AT&FV0E0�g���)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ��2��H6�^���Rφ��A�߶�q�������� ��5����� �ߏ�B߳������� �����1�C�*�g�� ,��P�b�t������ R�?���u0� ������������ ��M q���Z ���/�%/�� [/ 2�/�/h�/ /�/�/�3?�/W?>? {?�?@/�?d/v/�/�/ O�//OAOx?eO?�O�DO�O�O�O�O_�NIwTORÀG ?z��   	EX�EC1~s&R2,X3�,X4,X5,X��.V7*,X8,X9~s'R�2 �T+R�T7R�TCR�TOR �T[R�TgR�TsR�TR��T�R�S2�X2�X2��X2�X2�X2�X2��X2�X2�X2h3ʘX3�X37R2�R_�GRP_SV 1ݺ�� (�>�;�>y��m��B<H�
�������c����_D�B���cION�_DB<��@�zq�  �$��$�ϬY�1t�2p�>w��$�?$�ޡ
��@No   Qp�>{���p9p[�-u�d1�����8�P�G_JOG ��ʏ�{
�2�:��o�=���?����0�B��~\�n��������H�?��C�@�ŏ׏�N��  �����q�L_NAME �!ĵ8��!D�efault P�ersonali�ty (from� FD)qp0�RM�K_ENONLY��_�R2�a 1��L�XL�<8�gpl d���� şן�����1�C� U�g�y���������ӯ ���	����
�<�N� `�r���������̿޿� :��)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+��<�Sew�� �������/A�a��B�Bw��Pf��� ���/!/3/E/W/ i/{/�/�/�/���/ �/??/?A?S?e?w? �?�?�?�?�?�?�?�/ �/+O=OOOaOsO�O�O �O�O�O�O�O__'_`9_&O�S���x_�]�rdtS���_�]�_ �_�W�����S"oe_oXoa ��qogo yo�o�o�o�o�ouP�ph"|����	`[o Ugy8qK�A\��8��s� A ��y�@h�Q�Q��"����Tk\$�� W ��P�PE�x?C�  �I�@o a�<o��p�������ߏ 
f�Q*�����0��P�Cr� � �3r �.� @D��  A�?�G�-�?x.I�.@I�A�����  ;�	l�Y�	 �X?  ������� �, ǀ �����uPK��o�����]K���K]�K	�.��w�r_	����@
�)�b�1������I�Y������T;fY�{{S���3�����I�>J���;Î?v߮>��=@�����E��RѯעZ����wp��u�� D�!�3��7pg  �  �9��͏W���	'� �� u�I� ��  ��u��:��È��È=�s�ͱ���@��@ǰ�3��\�3�E��&���N�pC�  'AY�&�Z�i�b�@f��i�n�C����I�Ch����b��r0����ڟ.�B�p����q���}ر�.Dz Ə<ߛ�`�K�pߖ���w������А 4P�����.z��d  ��Pؠ?�ff0�_��	�� 2p>��P���8.f�t�>L����U���(.��P ���٨�����É���{ x��;e�m����KZ;�=g;�4�<<����%�G��3����p�?fff?ذ?&�S���@=0e�?��q�+�rN�Z� ��I���G���7���(� ����!E0iT�����+��F �p���#��D�� w����� ��//=/(/a/L/ �/p/��/�p�6�/ Z#?�/ ?Y?k?}?� �?�?>?�?�?�?�?�?�1O�����KD�y^KC�O�OO�O����`�O�O�O�Oai���1J��}�DD1���.B�D��@�AmQa��9N�,ȴA;�^@���T@|j@�$�?�V�>��z�ý��=�#�
>\)?��
=�G�-]��{=���,���C+��B�p���P��6���C98R����?N@��(��5�-]G�p�G�sb�F�}�G��>.E�VD��Kn���I��� F�W�E���'E���D���;n���I���`E�G���cE�vmD���-_�oQ_�o�o �o �o$H3X ~i������ ���D�/�h�S��� w��������я
��� .��R�=�v�a�s��� ��П����ߟ��(� N�9�r�]��������� ޯɯۯ���8�#�\� G���k�������ڿſ ���"��F�1�C�|� gϠϋ��ϯ����������P(�Q34�] �����Q�	�9�O��53~�mm��a�ǀ5Q�߫�aғ�����ߵ1��� ����1��U�C�y�g�J�%P�P���!�/���'���
���.������4�;�t�_��� ������������ :%��/�/d�������� 7%[Im���027�  B��S@J@�CH#PzS@�0@ZO/1/C/U/g/y/�-�#��/�/0�/�/�/�3?�3�� @�3��0ĵ0�13��5
 ?f?x?�?�?�?�? �?�?�?OO,O>OPO��Z@1 ���ۯ��c/�$MR_CABLE 2ƕ� ��TT �����ڰO���O�)�@ ���C_���_O_u_ 7_I__�_�_�_�_�_ o�_�_oKoqo3oEo {o�o�o�o�o�o�o�o �oGm/�K!�"���O����ذp�$�6���*Y��** �COM }ȖI���#��1 8u%% �2345678901���� ��Ï��R� � !� �!�
���Mnot sent b���W��TE�STFECSAL?GR  eg�*!�d[�41�
k�������$pB����������� 9UD1�:\mainte�nances.xsmlğ�  C:��DEFAU�LT�,�BGRP {2�z�  �� ���%  �%!�1st clea�ning of cont. v��ilation +56��ڧ�!0�����+B��*������+��"%��me�ch��cal c�heck1�  ��k�0u�|�� ԯ����Ϳ߿�@���?rollerS�e�w�ū��m�ϑϣ����@�Basic� quarterCly�*�<�ƪ,\��)�;�M�_�q�8�MXJ��ߓ "8��� ���ߕ �����+�=��C�g�ߋ�ʦ�߹���������@�Overha�u�ߔ��?� x� I�P����}���������� $n���� ���)l�ASew� ����� � +=O�s��� ����/R�9/ �(/��/�/�/�/�/ /�/�/N/#?r/G?Y? k?}?�?�/�???�? 8?OO1OCOUO�?yO �?�?�O�?�O�O�O	_ _jO?_�O�Ou_�O�_ �_�_�_�_0_oT_f_ ;o�__oqo�o�o�o�_ �oo,oPo%7I [m�o��o�o� ���!�3��W�� ������ÏՏ�6� ���l����e�w��� ������џ�2��V� +�=�O�a�s���� ��ͯ����'�9� ��]�������⯷�ɿ ۿ���N�#�r���Y� ��}Ϗϡϳ������ 8�J��n�C�U�g�y� ���ϯ������4�	� �-�?�Q��u����� �ߞ���������f� ;������������ �����P���t�I [m����� �:!3EW� {��� ��� //lA/��w/���/�/�/�/�/X*�"	� X�/?.?@?�)B a/o?m/o%w?�?�? }?�?�?OO�?�?OO aOsO1OCO�O�O�O�O �O__'_�O�O]_o_ �_?_Q_�_�_�_�_�_��\ Џ!?� ; @�! M?Ho Zolo�&4o�o�o�o�(�*�o** F�@ �Q�V�`o�'9�o]o�����/^&�o��� ��/�A�S�e��� #�����я����� +�q�����7������� k�͟ߟ��I�[��� K�]�o���C�����ɯ���o$�!�$M�R_HIST 2���U#�� 
 �\7"$ 2345?6789013�;���b2�90/���� [���./����ǿٿ F�X�j�!�3ρϲ��� {��ϟ�����B��� f�x�/ߜ�S����߉� �߭��,���P��t����=��$�SKCFMAP  �U�&��b
�� ����ONREL  �$#�������EXCFENB��
����&�FNC�-��JOGOVL�IM�d#�v���K�EY�y���_�PAN������R�UNi�y���SFSPDTYPM�<���SIGN���T1MOTk�����_CE_GRP7 1��U��+� 0�ow�#d�� ����&�6 \�7y�m� ��/�4/F/-/j/ !/t/�/�/�/{/�/�/�/?�+��QZ_E�DIT
����TC�OM_CFG 1����0�}?�?�? }
^1SI �NB����?�?���?�$O����?XO78T__ARC_*��X�T_MN_MO�DE
�U:_S�PL{O;�UAP_�CPL�O<�NOCHECK ?��/ �� _#_ 5_G_Y_k_}_�_�_�_��_�_�_�_oo��N�O_WAIT_L�	S7> NTf1�����%��qa_ERMRH2������� ?o�o�o�o��O�Gj�@O�cӦm| �T�GA�����A����<7G��(j3/@����<���?���)��n�b_PARAM�b����vHO��w
�.�@� = n�]�o� w�Q�����������`Ϗ�)���w�[��m� �����ODRD�SP�C8�OFFSET_CARI0��OǖDISԟœS;_A�@ARK
T9�OPEN_FIL�E��1T6�0OPTION_IO�����K�M_PRG ;%��%$*�����'�WO��N�s�ǥ�# ��5����G	 ������>d����RG_DS�BL  �����jN���RIENTkTO���C������A ��U�@IM�_DS���r��V~��LCT �{m�P2ڢ�3̹��d��<%���_PEX�@��n�RAT�G d8���̐UP ���:����S�e�KϬ�ϗ��$�r2G��L�XL���l㰂����� ��'�9�K�]�o߁� �ߥ߷����������#�5�G���2��v�� ������������e�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?�q1� ~?�?�?�?�?�?�?�?�O O2ODO�yA�a�m?~N��~O�O�P�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�O�Oo$o6o HoZolo~o�o�o�o�o �o�o�o �_oV hz������ �
��.�@�R�d�QO�ES������B�d�ӏ�ʏ����@����Y�D�}�0�� r���������ԟڟ��@�p���=�M��q��	`��������c�:�o�¯ԯ���>�A�  �k�TC�C�ڰ"ڰ����O��  ����-���)�C�  �t�k��� g�����Կ��ѿ
�5����_:�ĳ�OU����F��F�H���n�� �� ^�\� @oD�  p�?�v�b\�?:px�:qC4r��p�(��  ;�	�l��	 �X  ������� �,� � �������H�ʪ����H����Hw�zH���ϝ�8�<B���B�  Xѐ�x`�o�*��3����t�>u���fC{ߍ���:pB\�
�Ѵ=9:qK�t�� ����$���*���� DP�^���b�g  � � �h�����)�	�'� � ���I� �  y��'�=�������t�@����!�b��^;b�t�U�(�yN��r�  '��"E�C�И�t�C�И�`�ߗ���jA�@�����%�B�� ��,0���H:qDz�k��ߏz���݀������ 4P���:u�z:���	f��?�ff'�&8�� ]�m�8:p��>L�����$�(:p�P��	��`����:� x��;e�m"�KZ�;�=g;�4�<<���E/Tv���b���?ff�f?�?&� )�@�=0�%?�� �%_9��}!��$�x��/ v��/f'��W,??P? ;?t?_?�?�?�?�?�? �?O�?(OOLO�/�/ �/EO�OAO�O�O�O�O _�O_H_3_l_W_�_ {_�_�_1��_A���eO +o�ORooOo�o�o�o K/�o�omo�o*'`+�,�zt����CL�H��}?Ƀ����
�������u����D1��/n�t��p�q��@�I�h~,ȴA�;�^@��T@�|j@$�?��V�n�z������=#�
>�\)?��
=��G����{�=��,��C+��Bp�����6��C98R����?}p���(��5��G��p�Gsb�F��}�G�>.E�VD�KL�����I�� F��W�E��'E���D��;L�����I��`E��G��cE�vmD���\� ՟��ҟ���/��S� >�w�b�������ѯ�� �����=�(�:�s� ^���������߿ʿ� � �9�$�]�Hρ�l� �ϐϢ���������#� �G�2�W�}�hߡߌ� �߰��������
�C� .�g�R��v���� ����	���-��Q�<� u�`�r�����������@��'M�(��34�]O!����8h~�%3~�qm����5Q�������!���  `N��r��	eP@"P��Q�_/V/9/x$/]/H)����c/ j/�/�/�/�/�/�/�/ !??E?0?i?T?"&�_0�_�?�?�8��?�? O�?OBO0OfOTO�O@xO�O�O�O�O2f?_  B��pyp$QKCHR�z�p@� N_`_r_�_�_�_�]c�O�_�_oo+o�?�Bc� @Jd4�QJc�D
 2o�o�o �o�o�o�o%7�I[m��oa ������c/�$�PARAM_ME�NU ? ��  �DEFPULS�E��	WAIT�TMOUT�{R�CV� SH�ELL_WRK.�$CUR_STY�L�p"�OPT�8Q8�PTBM�G�C��R_DECSN �p������������ ��-�(�:�L�u�p���������qSSREL_ID  ���̕USE_P�ROG %�z%8���͓CCR�pޒ���s1�_HOST7 !�z!6�s��+�T�=���V�h����˯*�_TIME��rޖF��pGDE�BUGܐ�{͓GI�NP_FLMSK���#�TR2�#�PG�AP� ��_b�CyH1�"�TYPE�|�P������� �0�Y�T�f�xϡϜ� �����������1�,� >�P�y�t߆ߘ��߼� ����	���(�Q�L��^�p��%�WORD� ?	�{
 	�PR�p#MA9I��q"SUd���cTE��p#��	1���COLn%��!����L�� !���F�d�TRACE�CTL 1� ��q � #����_�_DT Q� ���z�D � � K`��c`�� _`������������@M`��k`���� $6�������� ����#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_8�^��� oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�.�o P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv���� ���*<N `r������ �//&/8/J/\/n/ Dϒ/�/�/�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z�����������$PGTR�ACELEN  ���  ������Ά_U�P ����2������΁_CFG ���S烸�
���*��:�D�O���O� � �O��DEF�SPD ��췁���΀H_C�ONFIG �\��� ����5dĔ�݂ ��ǑaP^�a�㑹��΀�IN�TRL ���=�8^���PEv��೗���p*�ÑO�΀LID����	T�LLB �1ⳙ ���BӐB4��O�� 䘼����Q�� << ��?�������M�3� U���i���������ӿ ��	�7�T�Ϣk� b�tϡ�诚���������S�GRP 1�������@A!�ߚ�4I���A ��Cu�C��OCjVF�/��Ȕa�zي�ÑÐ��t��ޯs������ӿߨ�B������������A�S�&�B34�_�������j������ ���	�B�-���Q����M�������  Dz ����.�����&L 7p[���� ���6!Zh�)w
V7.1�0beta1*��Ɛ@�*�@��) @�+A �Ē?��
?f�ff>����B_33A�Q�0��B(��A���AK��h���@�//'/9/P�p*��W�ӑ�n/�/�%����R�fh����*���P2�L R��/�/�/�/�/H?�Ĕ�I�u�&:�� �?��x?�?A���P!6\3 Bu�B��?�5SBH�3[4��o�L�4��[45��/B
\3x3Dx�?YO�?aOkO}O�<<�R@��O �C�O�O�O�O�DA�X��KNOW_M  �Z�%�X�SV 賚ڒ]��_ �_�_?�_�_�_o��Ԃ�W�M+�鳛 ���	@�3#����_�o�\A��o
]bV4�@u���u��e�o�l,�X�MR+��JmT3?��W��1C{�OADBA�NFWDL_V�ST^+�1 1����P4C���[��i/ �����?�1�C� ��g�y��������ӏ �*�	��`�?�Q�c�w2�|Va�up�<ʟ���p3��Ɵ؟Ꟃw4��+�=��wA5Z�l�~����w6����ѯ㯂w7 ��$�6��w8S�e�w����w+MAmp������OVLD  ���yo߄rPARNUM  �{+þ��?υqSCH�� ��
��X���{s��U�PDX�)ź��Ϧ�_CMP_@`���p|P�'yu�ER_C;HK���yqbb3��.�RSpp?Q'_MOm��_}ߥ��_RES_G�p���
�e�����0�#� T�G�x�k�}��������������׳��� ������:�Y�^��� Y�y������Ӭ����� ����������R� 6UZ�ӥ�u����V 1�FvpVa�@k�p��THR_INRp��(bzyudMASS� Z)MNGM�ON_QUEUE� �uyvup\!*��N�UZ�NW���END��߶EcXE����BE�|��OPTIO���ۚPROGRAoM %z%���~ϘTASK_�I��.OCFG ��z+�n/� DAkTACc�+�1}�-b2 �?�?/?A?S?]51  s?�?�?�?�?�6p1�?��?�?O"O,F�!IN+FOCc��-��bd lO~O�O�O�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_�_�_�/A@FD���, 	��!��K�_�!�)fN!fECNB��0m��Pf2Yo�khG�!2�0k �X,		d�=���·o���e�a$��pd��i�i�g_E?DIT ��/%�7����*SYS�TEM*upV9.�40107 cr7�/23/2021� A0Pw���PRGADJ_�p  h $X|[�p $Y�xZ�xW�xқtZқt?SPEED_�p�p�$NEXT_C�YCLE�p���q�FG�p ���pALGO_V� �pNYQ_F�REQ�WIN_�TYP�q)�SIuZ1�O�LAP�r�!�[��M+����qC?REATED�r��IFY�r@!NAM��p%h�_GJ�S�TATU��J�DE�BUG�rMAIL�TI����EVE<U��LAST������tELEM� �� $ENAB<�rN�EASI򁼁�AXIS�p$P�߄�����qROT�_RA" �rMAX� ��qE��LC�A�B
���C D_L9VՁ`�BAS��`��1�{���_� ��Y$x���RM� RB��;�DIS����X_cSPo�΁�� �u|�P� | 	�� 2 \�AN�� �;����8�Ӓ�� �0�PAYLO��3�V�_DOU�qS���p��tPREF� �( $GRID*�E
���R����Y� �pOTO|ƀ�q  �p℄!�p��k�OXY�� � $L��_PO|�נVa.�SRV��)����DIRECT_1T� �2(�3(�4(�U5(�6(�7(�8���qF��A�� �$VALu�GRgOUP���  ����� !���@!�������R#AN泲���R��/���TOTA��F���PW�I=!%�REGEN#�8���@����/���ڶnTz�����#�_S����8��(�V[�'���4���G#RE��w���H��D�܅���V_H��DAuY3�V��S_Y��Œ;�SUMMAR���2 $CONFIG_SEȃ8���ʅ_RUN�m��C�С�$CMPR:��P�DEV���_�I�ZP�*��q���ENHANCE*�	�
���1�N��INT��qM)b��q�2K����OVmRo�PGu�IX��;���OVCT�����>v�
 4 ����|a˟��PSLG"�>� \ �;��?�1���SƁϕc�U�����Ò��4�U�q]�Tp�G (`�-��rJ<��O� CK�IL_M�J���VN�+��TQ�n{�N5���C�U�LȀD�V(�C6�P�_�຀@�MW�V1VV�V1d�2s�2d�U3s�3d�4s�4d� �'�	�������p	�{IN	VIB1qp�1� 2!pq/,3* 3,4 4,�p ?��;��A���N��������PL��TO�Rr3�	��[�S{AV��d�MC_FOLD ?	$SL�����M,�I��L�� �pL�b��KE�EP_HNADD�	!Ke�UCCOMc�k��
�lOP���pl\��lREM�k���΢���U��enkHPW� K�SBM��ŠCOLLAB|�Ӱn��n��+�IT�O���$NOL�FCALX� �DON�r����� ,��FL|���$SYN�y,M�C=����U_P_DLY�qs"�DELA� ����Y�(�AD��$TA�BTP_R�# ��QSKIPj% ����OR� �E�� P_��� �)�� �p7��%9��%9A�$: N�$:[�$:h�$:u�$:t��$:9�q�RA��� X�����M}B�NFLIC]���0"�U!�o���NO�_H� �\�< _S�WITCHk�RA_PARAMG�O ��p��U���WJ��:Cӣ�NGRLT� OO�U���p��X�<A��T_Ja1�F�rAPS�WEI{GH]�J4CH��aDOR��aD��OO��)�2�_FJװ���saA�AV��C�HOB.��.�`�J2�0�q�$�EX��T$�'QIT��'Q�p�"'Q-�!η�RDC�m" G� ��<��
R]���
H���RGEAp��4��U�FLG`�g��H��ER	�SsPC6R�rUM_'P>��2TH2No��@�Q 1 ����0����  �D �وIi�2_P�25cS�ᰁ+�_L10_CI�Ad� �pk�� ��UՖD��zaxT�p�Q(�;a��c���޲+�i���e��`� P`DESIG\Rb$�VL1:i1Gf��c�g10�_DS���D��w�POS11�q l�pr��x1C/#AT�Br��U
WusIND�Ѐ}�mqCp�mq`B	�HGOME�r|�?t2GrM_q���`!
@s3Gr��� �(�$�6�4GrG�Y�0k�}����� `a�q5Grď֏����(��!@s6GrA�S�0e�w����� �0Ar7Gr��П�����0�8Gr;�M�_��q�����0�S �q    �@sM��P�B�K@��! T0`M��M�IO��m��I��2�OK _OPPy��� »Q)�R�p{WE" 7��x EQ�b � #�s%Ȳ$DSBo�G#NA�b� C�P2н��S232S�$� �iP��xc�I3CE<@%�PE`2�� @IT��P�OPB�7 1�FLOW�T�Ra@2��U$�CU8N��`�AUXT��2�>��ERFAC3İmUU��CH��'% t<_9�E���A$FREEF'ROMЦ�A�PX q�UPD"YbA�3PT.�pEEX0����!�FA%bҲ���RV�aG� &�  ��E�" 1�AL�  �+�jc�'��D�  2& ��S\PcP(
 ' �$7P�%�R�24� ��T�`AXU���DSP���@�W���:`$��RNP�%�@��z��K��_MIR������MT��AP����P"�qD�QSY�z������QPG7�B�RKH���ƅ AXI�  ^��i�����1 ����BSO�C���N��DUM�MY16�1$S�V�DE��I�FS�PD_OVR7d9� D����OR��֠N"`��F_����@�OV��SF�RU�N��"F0�����U�F"@G�TOd�LC�H�"�%RECOV��9@�@W�`&�ӂ�H��:`_0�  }@�RTINVE��.8AOFS��CK�KbFWD������1B,��TR�a�B �FD� ��1= B1pBL� �6� A1L�V��Kb����#��@+<�AM:��0��j��_M@ ~�@h���T$X`x ��T$HBK���F���AS����PPA�
��	����~��DVC_DB�3�@pA�A"��X1`�X3`��Se@��`�0��Uꣳ�h�CABPP
R�S #���c�B�@���GUBCPU�"��S�P�` R��11)ARŲ�!?$HW_CGpl�11� F&A1Ԡ@8p��$UNITr�|l e ATTRIr@�y"��CYC5B�C�A��FLTR_2_FI������z2bP��CHK_���SCT��F_e'F1_o,�"�*FS�Jj"CHA�Q�'91Is�82RSD����1���_Tg�`�L i�EM�NPMf�T&2 8p&2- �6�DIAGpERAI�LACNTBMw�L�O@�Q��7��PSı�� � ��PRRBSZ`�`BC4�&�	��FUN5s��RIN�PZaߠ�0�7Dh�RAH@���`�� `C�@�`C�Q�C�BLCURuH�DA0�K�!�H�HDAp�aA�H�C�ELD�������C��jA�1�CTI�BUu�8p$CE�_RIA�QJ�AF� P��>S�`DUT�2�0C��};OI<0DF_LC�H���k�LMLF�aH�RDYO���RG��@HZ0��ߠ�@�UM�ULSE�P�'3.iB$J��J�����FAN_ALM��dbWRNeHA#RD��ƽ�P��k@!2aN�r�J�_}��AUJ R+4�TO_SBR��~b�Іj�e 6?A�cMPIN�F��{!�d�A�cREG�NV��ɣZ�5D��NFLW%6r$M�@� ��f� ��0 h'uCM4NF�!�ON	 e!e�#�(b*r3F�3 �h	 ���q)5�$�g$Y�r��u�|_��p*$ �/��EG������qAR��i���2�3�u�@<�wAXE��ROB��7RED��WR��c�_���SY`��q� :?�SI�WRI���vE STհ�ӭ d���%Eg!���t8��^a"��B����9�3� �OTO�a���ARY��ǂ�1�����FIE���$LI�NK�QGTH���T_������390���XYZ����!*�OFF������ˀB��,B`l������m�FI� ���C@Iû�,B��_J$�F�����S`����3-!$1�w0��d�R��C��,�DU��r��3�P�3TUR`!XS.�Ձ�bXX�� ݗFL�d���pL��0���34���� +1)�K��M��5�5%B'��ORQ�6��fC㘴��0B�O;�D�,������aN�OVE��rM�� ���s2��s2��r1���`0���0�g /�AN=! �2�DQ�q���q�} R�*��6����s��V����ER��jA	�2E���.�C��A���0���XE�2Ӈ�A��AAX��F��A�N!�S� �1_��Q_Ɇ�^ʬ�^� ��^��0^ʙ�^ʷ�^�1&�^ƒP[ɒPkɒP {ɒP�ɒP�ɒP�ɒP �ɒP�ɒP�����ɪ ��R>�DEBU=#�$8ADc�2����
�A!B�7����V� <" 
��i�q��-! ��%��׆��׬��״� ���1�י��׷�JT���DR�m�LAB��8ݥ9 FGRO� ݒ=l� B_�1�u� ��}��`����ޥ��qa��AND�����qa� �Eq��`1��A@�� �NT$`��c�VEL�1��m���1u���QP��m�NA[w�(�CN1� ��3�줙��SERsVEc�p+ $@@�d@��!��PO�
�� _�0T !� �򗱬p, w $TRQ�b�
(� -DR2�,+"P�0_ .� l"@!�&ERR���"I� q���~TOQ����L�p]�e����0G��%��� �RE�@ / �,��/I -��RA~� 2. d�r&�"  0�p�$&��2tPM����OC�A8 1 � pCOUNT��� �qFZN_wCFG2 4B �f�"T�:#��Ӝ�ƞ ��`�s3 ���M:0�R�qC@0��/�:0�FA1P��?V�X�����r$���� �P:b.�HELpe4� 5��B_BA�S�cRSR�f @"�S�!QY 1�Y U2|*3|*4|*5|*�6|*7|*8�L!RaO�����NL�q� �AB���0Z ACmK��INT_u�US`�Pta9_PUX�>b%ROU��PH@��h9#�u`w�9�TPFWD_KAR�L�ar RE���PP��A]@QUE�i&��	�f�>`QaI`��9#��j3r��f�SEM�E��6��PA�ST�Y4SO�0�DI�'1�`���18�rQ_T}M�cMANRQXF��END�$K�EYSWITCH�j31:A�4HE	�BoEATM�3PE�pCLE��1��HU~3�F�42S?DDO_�HOMBPO:a0EF��PRr��*�v��uC�@O�Qo �O�V_Mϒ��Eq�O#CM���7��p8%;HK�q5 D��g�Uj�2M�p�4R���FORC�cWAeR��	:#OM�p 6 @�Ԣ�v`U|�P�p1�V'p�TE3�V4��*#O�0�L�R7��hUNLiOE0hdEDVa�  ���@d8 <�pAQ9�l1MSU�PG�UaCALC__PLANcc1���AYS1�@�9 '� X`��P � q;a�թ�w��2��j�M$P�㣒�fyt$��rSC�M�pm�q ����aq��0�tYzZ�zEU�Q�b�� T�!�Hr�pPvNPXw_ASf: 0g �ADD��$S{IZ%a$VA��~�MULTIP�"�]pq�PA�Q; � $T9op�B����rS��j!C~ �vF'RIF�2S�0�Y�T�pNF[DODB�UX�B��u&�!���CMtA�Е����������\Z ��< �3 �p�TEg���^��$SGL��T���X�&{���㰀��S�TMTe�ЃPSE�G�2��BW���S�HOW؅�1BAN�`TPO���gᣥ��Ԣ���.V�_Gv�= ��$PC��X�O�FB�QP\��SP�0A&0^���V�DG��>� �cA00�����P����P���P���P��5���6��7��8��9��A��b`���P��w���S`��F����h����1��v�h�י1�1��1��1�1�1�%�12�1?�1L�1�Y�1f�2��2��2���2ʙ2י2�2��2��2�2�2�%�22�2?�2L�2�Y�2f�3��3��3���3ʙ3י3�3P�����3�3%�U32�3߹3L�3Y�U3f�4��4��4��U4ʙ4י4�4�U4��4�4�4%�U42�4߹4L�4Y�U4f�5��5��5��U5ʙ5י5�5�U5��5�5�5%�U52�5߹5L�5Y�U5f�6��6��6��U6ʙ6י6��6�U6��6�6(�6%�U62�6߹6L�6Y�U6f�7��7��7��U7ʙ7י7��7�U7��7�7(�7%�U72�7߹7L�7Y��7f�ORV�`_UP�D��? �c� 
�PV���@ x $TOR�1T�  �cOP �, 6ZQ_7RE^��(� J��SsC�A���_U�p�Y�SLOA"A � �u$�v��w�@��x�@��bVALUv�10�6�F�ID�_L[C:HI5I~�R$FILE_X3�eu4$�C�SA�V��B hM �E_BLCK�3�ȁ>�D_CPU��p@��p5hz�pY���R3R C � �PW��� 	�!LAށSR�#.!.'$RUN�`G@%$ D!'$�@G%e!$e!'%�HR03$� '$��T2�Pa_LI�RD � � G_O�2>�0P_EDI�R@��T2SPD�#E��"i0ȁ�p�Q�D�CS9@G)F � 
$JPC71Tq�� S:C;C9�$MDL7$�5P>9TC�`@7UF�@?8S� ?8COBDu �@��"|�L�G�PE;;� 9:;����TAB'UI_�!L�HGb�%r�0FB3G$�3�A�sR�LLB_A�VAI�B�7�!��I� $� SEL� N�Ẽ�@RG_D N���TaOQ�3SC�P�J �1/AB�PT��RsD_M]`L�K 1\M f/QL_��F)Mj��PGi�U9R�]6��PS_�P\�� �p�EE7B�TB;C2�eL ���``l�`b$�!FT�Pp'T�`TDCg��� BPLp�sNU;WTHD��qhTgtWR�2{$�pERVE.S��T;S�Tw�R_AC�kP MX -$�Q�`.S�T;S�PU@r�`IC�`LOW�GF1�QR2g�`���p�S�ERTIA��d^0iP�PEkDE|Ue�LACEMzCC#c�V�BrpTf8�edg�aTCV�l�adgTRQ�l�e�j|� Scu��edcu�J7_ D4J!��Se@q
de�Q2�0���1�PlRcuPJKlvVK<� ~qcQ~qw�spJ0��q��sJJ�sJJ�sAAL�s�p�s�p�v��2�r5sS�`N1�l�p�k�`5dXA_́��vQCF�BN `M GROU ��bh��NPC0sD�REQ�UIR�R� EBU��C�Q�6g0 2aMz��Pd�QSGU�O�@�)APPR�0C7@� 
$� NN��CLO� ǉS^U�܉Se
Q�@A�"P �$PM]P�`�`sRN�_MGa!�C����+��0�@,�BRK�*�NOLD*�SHORTMO�!m�Z��JWA�SP�tp`�s p`�sp`�sp`�sp`�A
��7��8sQ!�QTQ� m��R.Q��cQ�PATH �*� �*��X&���-P�NT|@A�"p�l�� �IN�RUC4`�a��C�`UM��Y
`�)p��>�Q���cP���p��PAYL�OAh�J2L& R_Am@�L ������+�R_F2LgSHR�T/�LO����0���>���ACR@L0z�p�y�ޤsRH�5b$H+���FL[EX��_PJVR P��_._�_�_�QJ�US :�_�Vd`0�G��_tQ0d`�_�_lF1G��� ��o0oBoTofoxo��E�o�o�o�o�o�o�o  ����wz3lt��@��3EWF�^zT!��X�'qju��uu ~�W؁���p�u�u��u�u���� 	��(�T �P5�G�Y�' AT��l�pCEL0�_B��s�J��Sz�JEW�CTR�7B`NA��d�HA_ND_VB����TUO@`+�`TSW�tA�A�V� $$M� �e G�AV�Qs�De�oAA��@�	�$�A5�G�AU�A�d�� 6��G�DU�D�d�PD�G/ -ST�I�5V�5Ng�DY F ��+�x����P&� G�&�A��lw�o�Q�k�P������ʕӕܕ��RJUW 7 �� ��3%遞?!ASYMT���m�T�V�o�A�t�_SH�~������$ ����Ưد�J񬢐��#39"���_VI���`8�q0V_UCNIrS�4��.�Jmu �2��2A��4X��4�6 a�pt�������&E_�������E��CH~( X ̱l���TOc�PPСVsSvD�US�RU�P������z@�D�A}@_�5�U��P�EyAa��RP�ROG_NA��}$�$LAST����CANs�ISz@XYZ_SPu�DW]R@Ͱ,VSV@�E1QsENc��DCUR�H�' ��HR_T��YtQ9S�d���O�T%uP?�Z ��I�!A�D���Q ���#�S����3�vP [ � ME�O��R#B�!T�PPT0F@1�a��̰� h1a%i�T0� $D�UMMY1��$7PS_��RF��% �$lfװFLA�*�YP�bc$GLB_TI �U�e�`ձ��LIF(!\c����g`OW�P\��eVOL#qb &�a_2��[d2�[`�����b�P�cZ`TC~��$BAUDv���cST��B�2g`A�RITY0sD_W-AItAIyCJ2��OU6�ZqyyTL�ANS�`�{S�SZ<c��BUF_�r��fиx�PyyCHK_��@CES��� JO`E�aA�x�bUBYT����� r�.�.� ��aA��M��������Q] XXʰ����ST�����SBR@M21_�@��T$SV_E1R�b����CL�`��eA1�O�BpPGLh0�EW(!^ 4 m$a$Uq$�q$W�9�A�@]R�� �ӃUم�_ "��D$G�I��}$ف p��Ӄ�(!` L�\.��"}$F�"E6��NEAR��B$�F}��TQL�ic� �J�@R� �a7�$JOIN�Ta�o� ӃMS�ET(!b  +�E(c�2�^�ST�
H�_�(!c�  ��U��?���LOCK�_FO@� �PBG�LV��GL'�TE��@XM���EMPĹ���K��b�$1U�؂a�2_���Bq�`<� �q�^���CE/�?��� $K�ARb�M�STPD�RA܀����VECXX�����IUq�av�{HE�TOOL����V��REǠIS�3��6��ACH4̐m b^QONe[d�3���IdB�`@$�RAIL_BOXuEa���ROB�@�D�?���HOWW�AR0Aa�i`-�ROLMtb��$�*���T��`����O_FU�!}��HTML58Q S�� e�%Հ�(!d����@�(!!e���������@Ӄ�}p(!f t��m�^`a��t��B�PO�%�AIPE�N����O����q��AOR�DED�m �z�XIT`��A)mSP�O�P g D �`OB�����ǯ�Ucp�`��� ��SYS��ADR��pP`U@^ � h ,"��f$A��E��E�Q�PVWVA�Qi� � �@ق�UP�R�B�$EDI|�Ad�VSHWRU�z���IS�Uq�p�ND�P7���G�HECAD�! @���!i�3KEUqO`CP)P�֗JMP��L�U R�ACE�Tj����IL�S��C��N�E���TICK4!MKQC$���{HNr�k @���HWC��PHVF��`gSTYeB+�LO�a�g���[�C�l3�
L�@�F%$A��D=��S�!$�1�p aȌe�q�ePv HVSQ�U��#LO�b_1TGERC`! S?�m 5���R�m@3���ܡ��O`	c #IZ�d�A�eha�q�tb}�hA}pP~r��_SDO�B�X�pSSQN�SAXI�q��v��bS�U�@TL���RgEQ_ܠ��ET��(�`�CY%��FY'��YAf\!\d9x��P �RSR$$nl-�w �����c
�uV
Qh(��A���dC`�A���	�Y��D ��p�E"�	CC�AC��/�/�/	4 ���SSC�` o �h5�DSmడ[`S�P�@�AT� 
R���L��XbADDRf�s$Hp� IF�C�h�_2CH���pO�����- �TUk�Inr p�CUCpT#�V��I�Rq�P4���c��
K�
�RqV*���Pr \z��D����|,K� P�"C�N��*CƮ��!�TXSCREE��qs�Pp@�INA˃<�4�D�Q����`t Tᫀ�b�����O Y6���º�U4h�R�R�������R1�T����UE��u ��j �qz`Ś��RSML��U����V�1tPS_��6\��1�9G\���C��2@4� 2��0Ov�R��&F�AMTN_FL*�`Q��W���� �BBL_/�W�B`�Pw ����BO ��BLE"�Cg��R"�DRIGHtRyD��!CKGRB`��ET���G�AWIDTHs���RB��a�ro�UI��EYհRx d�ʰ����z�`y�BACK��h��>U���PFO��nQWLAB�?(�PyI��$URm��~P:�P�PHy1 �y 8 $�PT!_��,"�R�PRUp� s5�da�`�QO%!t�%zV�ȇ�pU�@�S9R ���LUM�S��� ERVJ���PP|��T{ � " �GE�Rh� �¯�LIPAeE��)^g@�lh�lh�ki5ik6ik7ikpP`�Z�x����$u1��p�Q� zQUSR�ل| <z��PU�2�a#2�FOO 2�P�RI*m9�[�@pT�RIPK�m�U�NDO��})� ��Yp��y����0i�����p ~�Rp�qG ��T���-!�rOS2��vR��2�s�CA�����r`�$��h�UIaCA���p�3Ib_�sOFFA�*D@���Ob�r�a5�L�t��GU���Ps������+QS�UB`� ��E_�EXE��VeуsW]O� �#��wF��WAl�p΁fP=
 V_DB��$�pT�pO�V░̷��3OR/�5�RA�U@6�TK���_<_���� |j ��OWNj�34$S#RC�0`���DA���_MPFI����ESP��T�$0��c���g�n�z�E!�# `%�ۂ34J���7COP��$`��p�_���/�+�6���C�T�Cہ�ہ�#�D�CS��P4��COMp�@ �;��O`�=����K�^�/�VT�q*'���Y٤Z��2�`��@p�w#SB��P��2�\0˰_��M�Ü%!]�DIC#��A�Y�3G�PEE�@T��QS�VR1���eQL�� a��P�D �� f�z��f�> ���6�p1A�t�b# �L2?SHADOW��#~ʱ_UNSCAd��׳OWD�˰DGD}E#LEGAC)�^q'��VC\ C��� v�������m�RF07���7d`yC2`7�DRIVo�	��ϠC�A]�(�` ����MY_UBY �d?Ĳ��s��1��$0�����_ఆ���mL��BM�A$�7DEY	�EXp@C�/�MU��X��,��0cUS����;p_R"1��0p#�2�GP�ACIN*���RG ��c�y�:�y��sy�C�/�RE�R"!�q8�y�D@� L !��G�P�"�Й �R�pD@�&P�Px1Q���	.���RE��SW&q�_Ar�u@+�{��Oq�AA/�3�hErZ�U���� �PV�HK���PJ���_/�Q0{�EAN���ۀ2�2�p�MR�CVCA� �:`O#RG��Q�dR	��L�����REFoG���� ��!�+`	�p���@�����<���q�_����r��� S�`C���Κ� �@D� ��0�!��#q�š��OU����?� ��Վ2�J@0� 1�*p����0� UL�@��C�O�0)��� NT�[��Z�Qf�af% L飏��Q|��a�VIAچ7� �ÀHD7 6P�$JO�`oB?�$Z_UPo��2Z_LOW��$�QiBn��1$EP �s�y�� 1!f� ��0æ4� m5�PA�A �oCACH&�LO�w�ВQB���CJn�I#F^��Tm�����$HO2�32{��Uÿ2O�@����Ro��=a��ƐVPx���@A"_SIZ&�K$Z$�F(�G'���C�MPk*FAIo�G���AD�)/�McRE���"P'GP�0�е�9�ASYNB;UFǧRTD�%�$�P!�COLE_2D�_4�5W�sw�~�U�ӍQO��%ECCU��VEM��v]2�VIRC�!5�#�2�!_>�*&�pWp���AG	9R�XYZ@�3�W���8��4d+Qz0T"��IM�1�6�2P�GRABqB�q��;�LERD�9C ;�F_D��F��f50MH�PE�R�[�����JRLAS��@��[_GEb�� �H൑~23�ET@����"���b��I�D��ҙ6m�BG_LEVnQ{�PK|Л6\q��GI�@N\P4���B��!g�dr�S$� �NRT�Lʁc��Ų��#a��c"!D�qDE����Xа�X��t6Q�1��d��pzZ���d�c����D4q�	  ��2pT��U&�� -$�ITPr9p[Q8��ՓV�VSF$�d��  fp/�f�U�R&���R`MZu9�dr��ADJ`C�v� ZDVf� D�X�AL� � 4 P�ERIKB$MS7G_Q3$Q!o%����p'��dr:g�qxQ� �XVR\t���B�pT_\��R _�ZABC"���ҨSr���
R���aA�CTVS' � � $|u�0�c�CTIV�Q!IO0u¥s&D�IT�x�DVϐ
x�P��i�!���pPS���� �#��!���q!LSTD�!�  �_ST���aq�;CHx�� L-�@���u�Ɛ*���P G�NA#�C�!q�_�FUN�� ��ZI�Pu��HR�$L���XZMPCF"��`bƀ�rX�فn��LNK��
Ł��0#�� $x !��ބCMCMk�EC8�C"����P{q? $J8�2�D6!>�O�H���T���`2�����M���UX�1݅UXE1Ѡ��1C� ��Y���������˗7�FTFG>�����Qp��� �k������YD'@ �� 8n�R� Uӱ?$HEIGHd�:h�?(! 'v��|���� � Gd��qp$B% � E���SHIF��hRVBn�F�`�HpC�  3�(�8H`O�ѡ�Cd��+%D	�"�CE�p�V�1�SPHE}Rs� � ,! �M�c�u��$PO?WERFL 4P|�e���|�p�RG�`  �������A� E ��?�p���pd���NSb ����?�  �Bz|� l�  <k@�|��%�涀�˃����ŵ�� �2ӷ�� 	H���l&���>ߪ��A |��t]$��*��/�� **:���p�ϥ�d�͘���������ɘ��|�����5� ������%ߟ�I�[� ��ߑ��������� ��w�!�3�a�W�i��� ���������O���� 9�/�A���e�w����� ��'����� =O}s���� ���k'UK ]������C/ ��-/#/5/�/Y/k/ �/�/�/?�/�/?�/ ?�?1?C?q?g?y?�? �?�?�?�?�?_O	OO IO?OQO����O�O �O_�E��3_���O`_��O�_�_÷PREF� Ӻ�p�p
���IORITY �4�|����p����pSaPL`z����WUT�V�qÈ�ODU~��e���_?�OG���Gx��R��,fHIB�qOy�|kTOEN�T 1��yP(!AF_t�`�o�g?!tcp�o}�!ud�o)~!icm�0b�XY̳�k �|�)� �����p����u��� ���N�5�r�Y���@����̏�����*/c̳ӹ���E�W�|��>�~F�F��/���4���|��,�7�A~��,  ��P�����%�|�'���Z��h�z�����|���ENHANCOE 	#�7�A9��d�����  �D,f�T
�_�S����OPORTe�rb�@��U��_CAR�TREP�Pr|brS�KSTAg�kSL�GS�`�k�����@Unothing�������Ϳ>�P�b�To��TEMP ?isϨE�/�_a_seibanm_��i_��� ��0��T�?�x�cߜ� �ߙ��߽������� >�)�N�t�_���� ����������:�%� ^�I���m��������� �� ��$H3l Wi������ �D/hS��w���uϪ�VE�RSI�P=g  �disabl�e��SAVE �?j	267_0H705���k/!�m//*�/ !	�(%b�O�+�/�S�e?6?H?Z?l?z:�%<�/�?4�*'_j` +1�kX �0ub�uE�?OqG�PURG�E��Bp`�ncqWF <@�a�TӒ*fW�`]D�aa�WRUP_DELAY z��f�B_HOT �%?e'b��OnER_?NORMAL�HGbx�O%_�GSEMI_�*_i_�QQSKIP�3.��3x��_� �_�_�_�]?eo+go Ko]ooo5o�o�o�o�o �o�o�o�o5GY i�}���� ���1�C�U��y� g���������я�����-�?�7%�$RA?CFG �[ќ��3�]�_PAR�AM�Q3y��S �@И@`�G�42�C۠��2��C�bFB�B]�BTI�F���J]�CVTMkOU�����]��DCR�3�Y ���Q<����B�w�BԢ�@���@H��;�+��]����$x�o������;e��m���KZ;��=g;�4�<�<���f@����� �5�G�Y�k�}� ������ſ׿���xU�RDIO_TYP�E  �V�5��E�DPROT_a��&>��4BHbbCEސSǆQ2c�7 ��B�ꐪ� ����ϐ����&�� ��W�V_~�o����� ����������A�O� m�r���9����� ���������=�_�d� �������������� ��'I�Nm�� ������� #EJi+k� �����//4/ F//g//�/y/�/�/ �/�/�/	?+/0?O/? c?Q?�?u?�?�?�?�?��??;?,O��S�INOT 2�I���l�G;� jO|K���<�O�f�0 �O�K �?�O�?___N_<_ r_X_�_�_�_�_�_�_ �_�_&ooJo8ono�o fo�o�o�o�o�o�o�o "F4j|b� ���������B�O�EFPOS1� 1"�  xO��o×O���� ݏ鈃���Ϗ0��T� �x����7���ҟm� �������>�P���� 7�������W��{�� ���:�կ^������ ����S�e��� ��$� ��H��l��iϢ�=� ��a��υ�� ߻��� �h�Sߌ�'߰�K��� o���
��.���R��� v��#�5�o������ �����<���9�r�� ��1���U��������� ��8#\���� ?��u��"� FX�?��� _��/�	/B/� f//�/%/�/�/[/m/ �/?�/,?�/P?�/t? ?q?�?E?�?i?�?�? O(O�?�?OpO[O�O /O�OSO�OwO�O_�O 6_�OZ_�O~_�_+_=_ w_�_�_�_�_ o�_Do��_Aozocf�2 1r�o.oho�o�o
 o.�oR�oO�# �G�k���� �N�9�r����1��� U����������8�ӏ \���	��U�����ڟ u�����"����X�� |����;�į_�q��� ���	�B�ݯf���� %�����[���ϣ� ,�ǿٿ�%φ�qϪ� E���i��ύ���(��� L���p�ߔ�/�A�S� ��������6���Z� ��W��+��O���s� �������V�A�z� ���9���]������� ��@��d��# ]���}�* �'`���C �gy��&//J/ �n/	/�/-/�/�/c/ �/�/?�/4?�/�/�/ -?�?y?�?M?�?q?�? �?�?0O�?TO�?xOOx�O�o�d3 1�o IO[O�O_�O7_=O[_ �O__|_�_P_�_t_ �_�_!o�_�_�_o{o fo�o:o�o^o�o�o�o �oA�oe �$ 6H�����+� �O��L��� ���D� ͏h�񏌏�����K� 6�o�
���.���R��� ퟈����5�ПY��� ��R�����ׯr��� ������U��y�� ��8���\�n������ �?�ڿc�����"τ� ��X���|�ߠ�)��� ����"߃�nߧ�B��� f��ߊ���%���I��� m���,�>�P���� �����3���W���T� ��(���L���p����� ������S>w� 6�Z���� =�a� Z� ��z/�'/�$/ ]/��//�/@/�/�O�D4 1�Ov/�/ �/@?+?d?j/�?#?�? G?�?�?}?O�?*O�? NO�?�?OGO�O�O�O gO�O�O_�O_J_�O n_	_�_-_�_Q_c_u_ �_o�_4o�_Xo�_|o oyo�oMo�oqo�o�o �o�o�oxc� 7�[���� >��b����!�3�E� ���ˏ���(�ÏL� �I������A�ʟe� ������H�3�l� ���+���O���ꯅ� ���2�ͯV���� O�����Կo������ ���R��v�Ϛ�5� ��Y�k�}Ϸ���<� ��`��τ�߁ߺ�U� ��y���&������� ��k��?���c��� ����"���F���j�� ��)�;�M������� ��0��T��Q�%��I�m��/�$5 1�/���m X���P�t� /�3/�W/�{// (/:/t/�/�/�/�/? �/A?�/>?w??�?6? �?Z?�?~?�?�?�?=O (OaO�?�O O�ODO�O �OzO_�O'_�OK_�O �O
_D_�_�_�_d_�_ �_o�_oGo�_koo �o*o�oNo`oro�o �o1�oU�oyv �J�n���� ���u�`���4��� X��|�ޏ���;�֏ _������0�B�|�ݟ ȟ���%���I��F� ����>�ǯb�믆� �����E�0�i���� (���L���翂�Ϧ� /�ʿS�� ��Lϭ� ����l��ϐ�ߴ�� O���s�ߗ�2߻�V� h�zߴ�� �9���]� �߁��~��R���v�����#�	6 1&����������� ����}���<�� `����CUg ��&�J�n 	k�?�c�� /���	/j/U/�/ )/�/M/�/q/�/?�/ 0?�/T?�/x??%?7? q?�?�?�?�?O�?>O �?;OtOO�O3O�OWO �O{O�O�O�O:_%_^_ �O�__�_A_�_�_w_  o�_$o�_Ho�_�_o Ao�o�o�oao�o�o �oD�oh�' �K]o�
��.� �R��v��s���G� Џk�􏏏���ŏ׏ �r�]���1���U�ޟ y�۟���8�ӟ\��� ���-�?�y�گů�� ��"���F��C�|�� ��;�Ŀ_�迃����� �B�-�f�ϊ�%Ϯ� Iϫ����ߣ�,���xP�6�H�7 1S� ���I��߲������ ��3���0�i���(� ��L���p�����/� �S���w����6��� ��l�������=�� ����6���V� z� 9�]� ��@Rd�� �#/�G/�k//h/ �/</�/`/�/�/?�/ �/�/?g?R?�?&?�? J?�?n?�?	O�?-O�? QO�?uOO"O4OnO�O �O�O�O_�O;_�O8_ q__�_0_�_T_�_x_ �_�_�_7o"o[o�_o o�o>o�o�oto�o�o !�oE�o�o>� ��^����� A��e� ���$���H� Z�l�����+�ƏO� �s��p���D�͟h� 񟌟���ԟ�o� Z���.���R�ۯv�د ���5�ЯY���}�c�u�8 1��*�<� v���߿��<�׿`� ��]ϖ�1Ϻ�U���y� ߝϯ�����\�G߀� ߤ�?���c����ߙ� "��F���j���)� c����������0� ��-�f����%���I� ��m������,P ��t�3��i ���:��� 3��S�w / ��6/�Z/�~// �/=/O/a/�/�/�/ ? �/D?�/h??e?�?9? �?]?�?�?
O�?�?�? OdOOO�O#O�OGO�O kO�O_�O*_�ON_�O r___1_k_�_�_�_ �_o�_8o�_5ono	o �o-o�oQo�ouo�o�o �o4X�o|� ;��q���� B����;������� [�������>�ُ�b�����!�������M�ASK 1 ��⤒���ΗXNO�  ݟ���MO�TE  ���S�_?CFG !Z����N�����PL_RGANGV�N������OWER "���Ϡ��SM_DRYPRG %����%W��եTAR�T #Ǯ�UME_PRO���q����_EXEC_E�NB  ����G�SPDJ�����Ρ�TDB����RM�п��IA_OPTgION��������NGVERS���`�řI_AIRPUR��� R�+���ÛMTE_֐T X���ΐ�OBOT_ISO�LC��������^��NAME8��H��ĚOB_CATEG�ϣ,��S�[��.�ORD_NUM� ?Ǩ���H705  �N��ߨߺ�ΐPC_TIMEOUT��{ xΐS232s��1$��� L�TEACH PENDAN��o����)��V�T��Maintena�nce Cons�N�&�M�"B�P�?No Use6�r� 8��������̒��GNPO$��Ҏ�"Ž��CH_LM��Q���	a�,�!OUD1:��.�RՐ�VAILw���|��*�SR  t�� ���5�R_I�NTVAL��� ���V_DA�TA_GRP 2�'���� D��P�������	� �����B 0RTf���� ��/�/>/,/b/ P/�/t/�/�/�/�/�/ ?�/(??L?:?p?^? �?�?�?�?�?�?�?O  O"O$O6OlOZO�O~O �O�O�O�O�O_�O2_  _V_D_z_h_�_�_�_ �_�_�_�_o
o@o.o�Povodo�o��$S�AF_DO_PU�LSW�[�S���i�S'CAN��������SCà(F��G���+S�S�
����P��q�q�qN� � L^p���5���� ��$���+��r2M�qqd�Y�P�`�J�	t/� @��������ʋ|�� r ք��_ @N�T ��'��9�K�X�T D��X���������ɟ۟ ����#�5�G�Y�k��}�������䅎������Ǧ  ="�;�oR� ����p"�
�u��Di���q$q�?  � ���u q%�\�������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$�6�H�Z����珈�� �����������g� ;�D�V�h�z�������@��������(�Ӣ0� r�i�y���$�7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/?r�+? =?O?a?s?�?�?�?�? �?8��?OO'O9OKO ]OoO�O��$�r�O �O�O�O	__-_?_Q_ c_u_�_�Y�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|�c�路g����� ��0�B�T�f�x����������ҏ����p��:�Ҧ��y��3�	�	123�45678��h�!B!�� +\��p0�� ��Ο�����(�:� @��c�u��������� ϯ����)�;�M� _�q�����R���ɿۿ ����#�5�G�Y�k� }Ϗϡϳ����ϖ��� ��1�C�U�g�yߋ� �߯���������	�� -���Q�c�u���� ����������)�;� M�_�q���B������ ����%7I[ m������� �!3EWi{ �������/ ///�S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?D/�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O*����O	_�E�?5_�G_Y_�yCz  �A��z   ���x2�r }��)�
�W_�  	�*�2�O �_�_ oo"l�#\��_hozo�o�o�o�o �o�o�o
.@R dv����Mo� ���*�<�N�`�r� ��������̏ޏ��� �&�8�J��X #P$Pt�Q�R<u� k�~�Q  �������S�P���Q�Qt�  �PÙ۟�P(� `,b����]��PFl�$SCR_�GRP 1*G�+G4� �� �,a ��U	 v��~������ d���%���ɯ���h]���P�D1� D7n��3��Fl�
CRX-10�iA/L 234�567890�P�d� r��Pd�L ��,a
1o�����Z���[ ¶~� +fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@��R�d�t���H�~�Ă�m��ϴ�@�����ϼ��,a�Ϡ1���U�[�G�imXh�uP,[~����B�  BƠߞҷ�r��A�P��  @1`��՚�@����� ?	���H����ښ�F@ F�`A� I�@�m�X��|���� ��������������`:�%�7�I�[�B�i� ��������������� -Q<u`��@En�ٯ���W�P�"+f@_�5��1`4b���x����ͣ�O�,dA����$���Fa�,a �#!"/4/E-!�Z(f/x/G/ (�P�!(� �/�/�/��/�/?#9b�����S7س�M�ECLV�L  ,a���ݲ�Q@f1L_D?EFAULTn4b1_�1`�3?HOTSTR�=���2MIPOWER�Fm0pU�5�4W7FDO�6 �5L��ERVENT 1�+u1u1�3 L!�DUM_EIP�#?5H�j!AF�_INE�0SO,d!'FT)O�NIO�O9!���O ��O�O�!RPC_MAIN�O�H��O>_S'VIS_�I�-_�_?!OPCUf�_�Wy_�_!TMP�PPU�_<Id�_�"o!
PMON_�PROXY#o?Fe ono�R<o8Mf]o�o�!RDM_SR�V�o<Ig�o!�R��"=Hh�oR!%
PM�o9LiA��!RLSYNC̟�y8��!gROS(O��4��6�!
CE�PMT'COM7�?Fk%���{!	K�CONS���>Glq�Ώ!K�WOASRC�o?Fm��v�!K�USB��=Hn	�f�!STM�0��;JoU����O�֟�c����CICE�_KL ?%K� (%SVCPGRG1��G�1�2G�DL�6�3o�t�6�4��D��6�5��į6�6��6�7��6���W�R�9_�d�3��� 6�9���6�a�ܿ6��� �6���,�6�ٯT�6� �|�6�)���6�Q��� 6�y���^����^�ʿ D�^��l�^�ϔ�^� Bϼ�^�j���^���� ^���4�^���\�^�
� �2���6��/� ���V��<�'�`�K� ��o����������� ��&J5nY� ������� 4F1jU�y� ����/�0// T/?/x/c/�/�/�/�/ �/�/�/??>?)?P?�t?_?�?
�_DEV� I�M{C:�84���4?GRP 2/E�0�+�bx 	�/ 
 ,@�0	A O!MC8OJO1OnOUO �O�O�O�O�O�O�O�O "_	_F_-_j_|_c_�_ �[O�_�_�_o�_,o oPo7oIo�omo�o�o �o�o�o�o(:!^�_  �t�C �����
��� @�'�d�K�]������� ����ۏ�o�N�"�U���T���� :�ϟ���ڟ�)�� M�4�]���j�����˯ ݯ�_����7��[� B����x�����ٿ� ҿ���3��,�i�P� ��䯂���^����ϴ� �ޙ�'��v�]ߚ� �߾��߷������*� �N��r��;��� ���������&�8�� \�C���g�y������� ����g�4-j Q�u����� B)fx_ ����)��/ ,//P/7/t/[/m/�/ �/�/�/�/?�/(??�L?^?E?�?�7d ��[~
�6 s� 	 A;*�=� 6?�=����D�>�����g�:�0���ī��|@��-�@�5_�e�A5�-�=B�G+h�&����6)AB�m����`x��=��?7O%TELE�OP8OcN[~y���5�o�ʾT�F�����������|��?ҝ����E�1��E@�*��A`�~�n�!���$�A����M�Y<T�������C=��J����Gc��McO��IJO/_��[~��6r �_�1<�׻���y;��	A`��ʛ1bP��N	V��A�&@в�@���@)E��]�1������0ד� x����Q��U?�Q��O�__ _o�DU�NU9��6�>���E��bQ�2]�j_ ���rAS��AT�@���@G$�_ �ߍyC� �Pr}���Q� 2i?�R�_�o�_�_�oDS �I�I�o*N<^�%��o�ho� ����(��L�� s��<���8���܏ʏ  ��$�f�K����~� l�������؟Ɵ��>� #�b��V�D�z�h��� ����ԯ���:�į.� �R�@�v�d���ܯ�� ӿ��������*��N� <�rϴ���ؿb��Ϻ� ������&��Jߌ�q� ��:ߤߒ��߶����� ��"�d�I���|�j� ��������*�P�!� `���T�B�x�f����� �����&�����* P>tb������ ���&L: p���`��� �/ /"/H/�o/� 8/�/�/�/�/�/�/? P/5?G?�/ ?�/h?�? �?�?�?�?(?OL?�? @O.OPOROdO�O�O�O  O�O$O�O__<_*_ L_N_`_�_�O�_�O�_ �_�_oo8o&oHo�_ �_�o�_no�o�o�o�o �o4vo[�o$�  ������N 3�r�f�T���x��� �����&��J�ԏ>� ,�b�P���t������� �"�����:�(�^� L���ğ����r���n� ܯ� �6�$�Z����� ��J�����Ŀƿؿ� ��2�t�YϘ�"ό�z� �Ϟ�������
�L�1� p���d�R߈�v߬ߚ� ���8�	�H���<�*� `�N��r������� ������8�&�\�J� �������p������� ��4"X���� H������
 0rW� �x� ����8///� /�P/�/t/�/�/�/ /�/4/�/(??8?:? L?�?p?�?�/�??�?  O�?$OO4O6OHO~O �?�O�?nO�O�O�O�O  __0_�O�O}_�OV_ �_�_�_�_�_�_o^_ Co�_ovoo�o�o�o �o�o�o6oZo�oN <r`���� �2�&��J�8�n� \�~����ˏ
����� �"��F�4�j����� ��Z�|�V�ğ���� �B���i���2����� ����������\�A� ��
�t�b��������� ���4��X��L�:� p�^ϔςϤ��� ��� 0���$��H�6�l�Z� ���Ϸ��π���|���  ��D�2�h�ߏ��� X�����������
� @���g���0������� ��������Z�?~� r`�����  ���8n \������ /� /"/4/j/X/�/ ��/�~/�/�/?�/ ??0?f?�/�?�/V? �?�?�?�?O�?On? �?eO�?>O�O�O�O�O �O�O_FO+_jO�O^_ �On_�_�_�_�_�__ oB_�_6o$oZoHojo �o~o�o�_�oo�o �o2 VDf��o ��o|��
��.� �R��y���B�d�>� ���Џ��*�l�Q� �����r�������ޟ ̟�D�)�h��\�J� ��n�������گ�� @�ʯ4�"�X�F�|�j� ����ٿ������ 0��T�B�xϺ���޿ h���d������,�� Pߒ�w߶�@ߪߘ��� �������(�j�O�� ��p��������  �B�'�f���Z�H�~� l�������������� ���� VDzh� ������
 R@v���f ����///N/ �u/�>/�/�/�/�/ �/�/ ?V/|/M?�/&? �?n?�?�?�?�?�?.? OR?�?FO�?VO|OjO �O�O�OO�O*O�O_ _B_0_R_x_f_�_�O �__�_�_�_oo>o ,oNoto�_�o�_do�o �o�o�o:|oa s*L&���� ��T9�x�l�Z� |�~���Ə���,�� P�ڏD�2�h�V�x�z� ����(����
� @�.�d�R�t�ʟ���  ��������<�*� `�����ƯP���L�ʿ �޿��8�z�_Ϟ� (ϒπ϶Ϥ������� �R�7�v� �j�Xߎ� |߲ߠ�����*��N� ��B�0�f�T��x�� �����������>� ,�b�P��������v� ��������:(^ �����N���� �� 6x]�& �~�����> d5/t/h/V/�/z/ �/�/�//�/:/�/.? �/>?d?R?�?v?�?�/ �??�?O�?*OO:O `ONO�O�?�O�?tO�O �O_�O&__6_\_�O �_�OL_�_�_�_�_�_��_"od_Io[ob  ��$SERV_MAIL  �U��`��QvdOUT�PUT�h��P@vdRV 2�0f  �` (�a\o�ovdSAVE��l�iTOP10 �21�i d �6 s�P6r _>q2oXj|� �������� 0�B�T�f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�gu�YP�cFZN_�CFG 2e��c�T�a�e|�G�RP 23��q ,B   AƠ~�QD;� BǠ��  B4�S�RB21�fHELL�4ev�`�o���/�>�%RSR>�?�Q���u����� ҿ������,��PϠ;�t�_Ϙϩ����  �¼���(�Ϸͻ��P�&Ҧ'�ސW��2�Pd���g��HK 15�� ,ߡ߫� ����������@�;� M�_���������������OMM �6��?��FTOV_ENB�d�au��OW_REG_U�I_��bIMIOFWDL*�7.�ɥ��/WAIT\�`ٞ�ȼ��`���d��TI�M������VA��`����_UNIT�[�*yLCy�TR�Y��uv`ME�8���aw֑d ���9� ���j��<��X�Pxڠ6p`?�  � �o+=IpVL�l�fMON_�ALIAS ?e.��`heGo�� ����/)/;/M/ �q/�/�/�/�/d/�/ �/??%?�/I?[?m? ?�?<?�?�?�?�?�? �?!O3OEOWOO{O�O �O�O�OnO�O�O__ /_�OS_e_w_�_�_F_ �_�_�_�_�_o+o=o Ooaoo�o�o�o�o�o xo�o'9�o] o��>���� ��#�5�G�Y�k�� ������ŏ׏����� �1�C��g�y����� H���ӟ���	���-� ?�Q�c�u� ������� ϯᯌ���)�;�� L�q�������R�˿ݿ ��Ͼ�7�I�[�m� �*ϣϵ������ϖ� �!�3�E���i�{ߍ� �߱�\��������� ��A�S�e�w��4�� ����������+�=� O���s���������f� ����'��K] o��>���� �#5GY}�����l�$S�MON_DEFP�ROG &����� �&*SYSTE�M*���REC�ALL ?}�� ( �}8co�py frs:o�rderfil.�dat virt�:\tmpbac�k\=>192.�168.56.1?:15124/�/�/�-}/K"mdb:*.*`/r/{/?�?0?�$3xK$:\ �/U0�/0�/�?�?�?
� 4K5aS?e?�%�?�O#O5O }
xy�zrate 11 �?�?�?�O�O�O�%9KGkL880� jO�|O__1_�#tp�disc 0�O4� �O�O�_�_�_�&�tpconn 0 T_f_x_	oo-o@O RA�_�_�_�o�o�o�%y�Ow&716 jo |o1�#K_�h �o�o����_Tf x	��-�@oRm�� �������o�o�or�� �'��-J/\/�/恃� �����/�/g�߈{�� �0�C?ԟhO����� �����?X�j�瀀�� #�5�HOگ�������x���O�4772ho@z���/�B_ֿ � ���ϜϮ���\b�t���)߼�7K�]�S�!27ߓߥ�8�.˟f�@޸z���/�2K� ^�ڼ�ߏ���F�ӯ d����"�4�G�Y� ���ߎ�������`��� {�0C�����y� �������d�� ,?�Q���u��� �����j��//(/ ;M�q�/�/�/� �\/��/?$?6?I� �/�/�/�?�?�?Ǐ�344�z?OO/O B�?ea�?�?�O�O�O ��VOhOzO__/_B� T��9�_�_�_����g_�8{_oo0oCS��$SNPX_AS�G 2:����Va� � 0DQ%�7o~o � ?�GfPARAoM ;Ve`a� �	lkP>T�DP>X�d� ���I`OFT_K�B_CFG  �CS\eFcOPIN_�SIM  Vk��b+=OYsI`R�VNORDY_DOO  �eukr�QSTP_DSB�~�b�>kSR �<Vi � & TELEO�e��{v>TW`I`TOP_ON_ERRx�Gb�PTN zVeP��D:��RING_PRM�'��rVCNT_GOP 2=Ve�ac`x 	���DP��яؼ���BgVD�RP' 1>�i�`�Vq ؏0�B�T�f�x����� ����ҟ�����,� >�e�b�t��������� ί���+�(�:�L� ^�p���������ʿ� � ��$�6�H�Z�l� ~ϐϷϴ��������� � �2�D�V�}�zߌ� �߰���������
�� C�@�R�d�v���� ������	���*�<� N�`�r����������� ����&8J\ n������� �"4[Xj| �������!/ /0/B/T/f/x/�/�/ �/�/�/�/�/??,? >?P?b?t?�?�?�?�?��?�?�?O�PRG�_COUNT�f9�P�)IENBe�+E�MUC�dbO_UPD� 1?�{T  
ODR�O�O�O�O�O __A_<_N_`_�_�_ �_�_�_�_�_�_oo &o8oao\ono�o�o�o �o�o�o�o�o94 FX�|���� �����0�Y�T� f�x����������� ���1�,�>�P�y�t� ��������Ο��	�� �(�Q�L�^�p����� �����ܯ� �)�$� 6�H�q�l�~������� ƿؿ���� �I�D��V�"L_INFO {1@�E�@��	 yϽϨ������?��?w~�>B|<����� A��A_�e�T���?3�L��������j`� >�` =U�<�@ =����� D58o�G���C˃]�3�����n����bp߂�-@YSDOEBUG:@�@�o��d�I��SP_PA�SS:EB?��L_OG A���A�  o�i�v� � �Ao�UD�1:\��}���_M�PC�ݚEk�}�A�&�� �AK�SAV B��IA���*�i�1�SVB�T�EM_TIME �1C���@ 0o  n��i��f��*���MEMBOK  �EA��������X|΀@� @��n��@��������h�9
�� ��@�`r �������� �@Rd�v�����
Le �//(/:/L/^/p/ �/�/�/�/�/�/�/ ?�?$?6?H?Z?��SK V�[�EAj��?�?�?��+(�@]2���?>i�  0�o�^ 
:O.@R�O�O�O8}N�mҀ ��OB �C__,_ P_G2Dt_�_�_�_�_�]$�_�_�o'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk�_?T1SVGUNwSPD�� '�����p2MODE_?LIM D���2�t2�p�qE�݉u�ABUI_DCS' H}5���0�G�n��D��|-�X��>���*���� !
��e��i���r��i�����uED�IT I��xS�CRN J��<�rS�G K�.��(�0߅SK_OPTION��^�����_DI��ENB � -����BC2_GRP 2L�a��MPC�ʓ^�|BCCF/�N����� ����` �>�W�B�g���x��� ��կ�������� S�>�w�b��������� Ͽ�����=�(�a� Lυϗ�Ň�϶����� ��v��
�/�U�@�y� ���`�iМ��߰��� ��
���.��>�@�R� ��v���������� �*��N�<�r�`��� ������������̀ 4FX��|j� ������ B0fTvx�� ���/�,//</ b/P/�/t/�/�/�/�/ �/�/�/(??L?d? v?�?�?�?6?�?�?�? O O6OHOZO(O~OlO �O�O�O�O�O�O�O _ _D_2_h_V_�_z_�_ �_�_�_�_
o�_.oo >o@oRo�ovo�ob?�o �o�o�o<*L r`������ ��&��6�8�J��� n�����ȏ���ڏ�� "��F�4�j�X���|� �������֟��o$� 6�T�f�x��������� ү�������>�,� b�P���t�������� ο��(��L�:�\� ��pϦϔ��ϸ����� �� ��H�6�l�"��� �ߴ�����V������ 2� �V�h�z�H��� �����������
�@� .�d�R���v������� ������*N< ^`r������ �&8�\Jl �������� "//F/4/V/X/j/�/ �/�/�/�/�/?�/? B?0?f?T?�?x?�?�? �?�?�?O�?,O�DO VOtO�O�OO�O�O�O��O�O_ V4P�$T�BCSG_GRP� 2O U��  �4Q 
? ?�  __q_ [_�__�_�_�_�_�_�o%k8R?SQF\d��HTa?4Q	� HA���#e>�>$a�\~#eAT��A WR��o�hdjma�G�?�Lfg�bp�o�n�ffhf��ͼb4P|jy��o*}@��Rhf�ff>�33pa�#e<qB�o+=xr�Rp�qUy�rt~���H�y rIpTv�pB� �t~	xf	x(�;�� �f���N�`���ˏڋ�����	V3.�00WR	crxlڃ	*��3R�~t��HH��� �\�.�]�  cCa.�����8QJ2?S�RF]����CFG� T UPQ �SPܚ��r�ܟ1��1�W�e� 	Pe���v�����ӯ�� ������Q�<�u� `���������Ϳ�޿ ��;�&�_�Jσ�n� �ϹϤ�������WR q@�0�B���u�`߅� �ߖ��ߺ������)� ;�M��q�\���� ��4Q _���O ��� J�8�n�\��������� ��������4"X Fhj|���� ��.TBx f��nO���� //>/,/b/P/�/t/ �/�/�/�/�/�/�/? :?(?^?p?�?�?N?�? �?�?�?�?�? O6O$O ZOHO~OlO�O�O�O�O �O�O�O __D_2_T_ V_h_�_�_�_�_�_�_ 
o�_o@o�Xojo|o &o�o�o�o�o�o�o *N`r�B� ������&�� 6�\�J���n�����ȏ ��؏ڏ�"��F�4� j�X���|���ğ��� ֟���0��@�B�T� ��x�����ү䯎o�� �̯ʯP�>�t�b��� �����������Կ &�L�:�p�^ϔϦϸ� �τ������ �"�H� 6�l�Zߐ�~ߴߢ��� �������2� �V�D� z�h���������� ���
�,�.�@�v�� ������\������� <*`N��� �x���8 J\(���� ����/4/"/X/ F/|/j/�/�/�/�/�/ �/�/??B?0?f?T? v?�?�?�?�?�?�?O O��2ODO�� O�OtO �O�O�O�O�O_�O(_ :_L_
__�_p_�_�_ �_�_�_ o�_$oo4o 6oHo~olo�o�o�o�o �o�o�o D2h V�z����� 
��.��R�@�b��� v���&OXO֏菒��� ��N�<�r�`����� ��̟ޟ🮟��$� &�8�n�������^�ȯ ���گ��� �"�4� j�X���|�����ֿĿ ����0��T�B�x� fψϊϜ��������� ��>�P���h�zߌ� 6߼ߪ���������� :�(�^�p���R�������� ���  &�*� *�>�*���$TBJOP_�GRP 2U����  �?���C*�	�V�]�Wd������X  �*��� �, � ���^*� @&�?��	 �A�����?C�  DD������>v�>\?� ��aG�:��o��;ߴAgT������A�<���MX����>��\)?���8�Q�����L��>y�0 &�;iG.��Ap< � F�A�ff�v��� x):VM�.��� S>o*�@�;�R�Cр	���������ff��:�6/�?�{33�B   � �/������^>):�S����x �/�/@��H�%�&/�/��=� <�#�
*��v�;/��ڪ!?���4B�3?'?2	��2?h Z?D?R?�?�?�?F?�? �?�?�?OAOO�?`O�zOdOrO�O�O*�C��*���A��	V3�.00{�crxl��*P��%�%�c5Z F�� JZH F6�� F^ F��� F�f F�� G� G5� G<
 G^]� G� G����G�*�G�S� G�; G���ERDu�\E[�� E� F(� F-� FU`� F}  F�N� F� F��� Fͺ F�� F�V G�� Gz Ga� 9ѷ�Q�LHDefJ4�o,b*��0c1���OH�ED_TCH Xd�,+X2S�&�&��d$'X�o�o*�1�F�TESTPAR�S  ��cV�H�RpABLE 1Yd� N`*������g$j�g�hP�h)�1��g	�h
�hQ�hHu*��h�hu�h%vRDI0n�GYk}��u	�O�#�-�?�Q�c�$u�)rS�l� �z6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z���I���m�Fw ͩ��ȏڏ쏘������x)r��NUM�  ��n����2� Ep�)r_?CFG Z��I����@V�IMEBFG_TTqD��e޶GVER�����޳�R 1[8{ 8I�o*�%�Q� ��د  9�K�]�oρ� �ϥϷ���������� #�5�G�Y�k�}��ߡ� ������������1� ��E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oĩ_���@��`L�IF \���D`����DR�(�FP
�!p�!p�� d� ��MI_CWHAN� � �DBGLVL���fETHERAOD ?u��0`�1�_}�RO�UT�!�j!���SNMAS�KY�j255.%S///A/S�`�OOLOFS_D�Ip�CORQCTRL ]8{��1o�-T�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OL�/�6O%OZOcPE_D�ETAI7�*PG�L_CONFIG� c�������/cell/$C�ID$/grp1�^O�O�O�O
__|�� �G_Y_k_}_�_�_0_ �_�_�_�_oo�_Co Uogoyo�o�o,o>o�o �o�o	-�oQc u���:��� ��)���_�q���������׮}N��� �%�7�I�a�KOq�P��M�����ʟܟ� � G�$�6�H�Z�l�~�� ����Ưد������ 2�D�V�h�z������ ¿Կ���
ϙ�.�@� R�d�vψϚ�)Ͼ��� �����ߧ�<�N�`� r߄ߖ�%ߺ������� ��&��J�\�n�� ���3���������� "���F�X�j�|���������@�User View �I�}}1234567890�����+=Ex �e����2��B����� �`r��3�O as����x4>//'/9/K/]/�~/x5��/�/�/@�/�/?p/2?x6�/ k?}?�?�?�?�?$?�?x7Z?O1OCOUOgOyO�?�Ox8O�O�O��O	__-_�ON_TR �lCamera���O�_�_�_�_�_�_˂E�_o)o ;n��Uogoyo�o�o�o�)  mV�	�_�o #5GY o}�� �o������F_�mV=�k�}����� ��ŏl����X�1� C�U�g�y���2�D�� "�ן�����1�؏ U�g�y�ğ������ӯ �����D��k��E�W� i�{�����F�ÿտ� 2���/�A�S�e�� nUY9������������ 	߰�-�?�Qߜ�u߇� �߽߫���v�D�If� �-�?�Q�c�u�ߙ� ����������)� ;���D��I������� ��������)t� M_q���N�`�93��0B ��Sx�1������//�J	oU0 �U/g/y/�/�/�/V �/�/�/�?-???Q? c?u?/./tPv[?�? �?�?OO(O�/LO^O pO�?�O�O�O�O�O�O �?oU�k�O:_L_^_p_ �_�_;O�_�_�_'_ o o$o6oHoZo_;%N� �_�o�o�o�o�o �_ $6H�ol~�� ��moe��]�$� 6�H�Z�l������� �؏���� �2�� e&�ɏ~�������Ɵ ؟���� �k�D�V� h�z�����E�e��5� ���� �2�D��h� z���ׯ��¿Կ���<
ϱ�  ��9� K�]�oρϓϥϷ���x������   � �5�G�Y�k�}ߏߡ� ������������1� C�U�g�y������ ������	��-�?�Q� c�u������������� ��);M_q��  
��(  ��-�( 	  �������# 35G}k��t��
� �Y� 
//./��R/d/v/�/ �/�/����/�/�/A/ ?0?B?T?f?x?�/�? �?�??�?�?OO,O >O�?bOtO�O�?�O�O �O�O�O_KO]O:_L_ ^_�O�_�_�_�_�_�_ #_ oo$ok_HoZolo ~o�o�o�_�o�o�o1o  2DVh�o�o ���	��
�� .�@��d�v������ ��Џ���M�*�<� N���r���������̟ �%���&�m�J�\� n��������ȯگ� 3��"�4�F�X�j��� ��������ֿ���� �0�w���f�xϊ�ѿ �����������O�,� >�Pߗ�t߆ߘߪ߼� �������]�:�L��^�p����߻@ A������������� ��"frh:�\tpgl\ro�bots\crx�!�10ia_l.xml��D�V�h�z��������������������0BTfx ��������� ,>Pbt�� ������/(/ :/L/^/p/�/�/�/�/ �/�/��/?$?6?H? Z?l?~?�?�?�?�?�? �/�?O O2ODOVOhO zO�O�O�O�O�O�?�O 
__._@_R_d_v_�_ �_�_�_�_�O�_oo *o<oNo`oro�o�o�oкo�o�n �6� ����<< 	� ?��k!�o ;iOq���� �����%�S�9��k���o�����я�����(�$TPGL�_OUTPUT sf������ �&�8�J�\� n���������ȟڟ� ���"�4�F�X�j�|�@������į�p�ր�2345678901�����1�C� K����r��������� ̿d�п��&�8�J��}T�|ώϠϲ��� \�n�����0�B�T� ��bߊߜ߮�����j� ����,�>�P����� ���������x��� �(�:�L�^���l��� ��������t���$ 6HZlz�� ����� 2D Vh ���� ���/./@/R/d/ v//�/�/�/�/�/�/��/ۂ $$ ��ί<7*?\?N?�?r? �?�?�?�?�?�?OO 4O&OXOJO|OnO�O�O �O�O�O�O_�O0_"_T_}�an_�_�_�_�_��_�]@�_o	z? ( 	 V_Do 2ohoVo�ozo�o�o�o �o�o
�o.R@ vd������ ���(�*�<�r�`����ܦ�  <<I_ˏݏ���� ���:�L�֪��}��� )���ş�������k� �C�ݟ/�y���e��� ����������-�?� �c�u�ӯ]�����W� ��Ϳ��)χ���_� q��yϧρϓ����� M��%߿��[�5�G� �ߣ�߫���s���� !���E�W��?��� 9���������i��� A�S���w���c�u��� �/�����= )s�����U� ��'9�!o 	[�����K �#/5/�Y/k/E/w/ �/�/�/�/�/�/? �/?U?g?�/�?�?7?��?�?�?�?	OO��)�WGL1.XM�L�_PM�$TPOFF_LIM ��|�P���^F�N_SVf@  ��TxJP_MON7 g��zD�P��P2ZISTRT?CHK h��xF�k_aBVTCOM�PAT�HQ|FVW�VAR i�M\:X�D �O R_��P�BbA_DE�FPROG %��I%TELE�OPi_�O_DIS�PLAYm@�N�RI�NST_MSK � �\ �ZIN�USER_�TLC�Kl�[QUICK�MEN:o�TSCR�EY`��Rtpsc�Tat`yi4xB�`_�iSTZxI�RACE_CFGW j�I:T�@�	[T
?��hHNL 2k�Z���aA[ gR-?Qcu����z�eITEM� 2l{ �%�$1234567�890 ��  =�<
�0�B�J�  !P�X�dP���[S ���"���X�
�|� ��W���r�֏����.� �0�B�\�f�����6� \�n�ҟ�������� >���"���.����� ίR����Ŀֿ:�� ^�p�9ϔ�Tϸ�xϊ� ��d���H��l� �>�Pߴ�\������� v� ������h�(�� �߰�4�L��ߦ��� ��@�R��v�6���Z� l���������*��� N��� ���������� ��X���J
 n���b�� ��"4F�/| </N/�Z/���// �/0/�/?f/?�/�/ e?�/�?�/�?�?�?,? �?P?b?t?�?�?DOjO |O�?�OOO(O�O�O ^O_0_�O<_�O�O�_ �O�__�_�_H_�_l_(~_Go�dS�bm�oLj��  �rLjq �a�o�Y
 �o��o�o�o{jUD1�:\|��^aR_�GRP 1n�{� 	 @�P Rd{N�r����~��p���q+�x�O�:�?�  j� |�f����������ҏ ����>�,�b�P���`t���������	e����\cSCB 2ohk U�R�d� v���������Я�Rl�UTORIAL �phk�o-�WgV_�CONFIG �qhm�a�o�o��<�O�UTPUT r<hi}�����ܿ � ��$�6�H�Z�l� ~ϐϢϴ�z�ɿ����  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������� �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/��/�/?? 0?B?T?f?x?�?�?�? �?�/�?�?OO,O>O PObOtO�O�O�O�O�? �O�O__(_:_L_^_ p_�_�_�_�_�_f�x� ǿoo,o>oPoboto �o�o�o�o�o�o�O (:L^p�� �����o ��$� 6�H�Z�l�~������� Ə؏��� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я�� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� ���������������X���# ��N�_r���� ���&8J ��n������ ��/"/4/F/X/i |/�/�/�/�/�/�/�/ ??0?B?T?e/x?�? �?�?�?�?�?�?OO ,O>OPOa?tO�O�O�O �O�O�O�O__(_:_ L_^_oO�_�_�_�_�_ �_�_ oo$o6oHoZo k_~o�o�o�o�o�o�o �o 2DVgoz �������
� �.�@�R�d�u���� ����Џ����*� <�N�`�q��������� ̟ޟ���&�8�J��\�k��$TX_S�CREEN 1s�% �}�k�����ӯ���	���Z��I�[�m� ������,�ٿ��� �!�3Ϫ�W�ο{ύ� �ϱ�����L���p�� /�A�S�e�w��� ߭� ���������~�+�� O�a�s���� ��� D�����'�9�K��� �������������R� ��v�#5GYk}�����$UALR�M_MSG ?����� �n�� �	:-^Qc ������ /��SEV  ��2&�ECFG �u����  }n�@�  Ab!�   B�n�
 /u����/�/�/�/ �/�/??%?7?I?W7~>!GRP 2vH+w 0n�	 /��?� I_BBL_NOTE wH*�T��l�u���w�T �2DE�FPRO� %� (%�Ow�	OBO -OfOQO�OuO�O�O�O��O�O_�O,_�<FK�EYDATA 1yx���0p W'n��?�_�_z_�_�_ưZ,(�_on�(�POINTo>o �POOK ,ojoQa?NDIRECYomo�  CHOICE�]�onTOUCHUP�o�o�o�o 8\nU�y� �����"�	�F���Y��/frh�/gui/whi�tehome.pngQ�������ŏ׏��h�point�z���/�A�S�� = i�look�����������ɟ۟j�indirec���'��9�K�]�h�choicy�������ͯ߯��h�touchup���/�A�S�e��}h�arwrg� ����ÿտ�n��� (�:�L�^�p����Ϧ� ��������}��$�6� H�Z�l��ϐߢߴ��� �����ߋ� �2�D�V� h�z�	��������� ����.�@�R�d�v� ��_������������� �2DVhz� �����
� @Rdv��) ����//�</ N/`/r/�/�/%/�/�/ �/�/??&?�/J?\? n?�?�?�?3?�?�?�? �?O"O�?4OXOjO|O �O�O�OAO�O�O�O_ _0_�OT_f_x_�_�_ �_=_�_�_�_oo,o >o�_boto�o�o�o�o�W��k�b�����o}�o8J$v,6�{.��� ������/�� S�:�w���p�����я �ʏ��+��O�a� H���l�������ߟ� ��'�9�Ho]�o��� ������ɯX����� #�5�G�֯k�}����� ��ſT������1� C�U��yϋϝϯ��� ��b���	��-�?�Q� ��u߇ߙ߽߫����� p���)�;�M�_��� ���������l�� �%�7�I�[�m���� ����������z�! 3EWi����� ����П/A Sew~���� ��/�+/=/O/a/ s/�//�/�/�/�/�/ ?�/'?9?K?]?o?�? �?"?�?�?�?�?�?O �?5OGOYOkO}O�OO �O�O�O�O�O__�O C_U_g_y_�_�_,_�_ �_�_�_	oo�_?oQo couo�o�o�o:o�o�o �o)�oM_q ���6������%�7�9��>���b�t� ��^�������,��� �����3�E�,�i�P� ������ß������� ��A�S�:�w�^��� ����ѯ����ܯ�+� 
O�a�s�������� Ϳ߿���'�9�ȿ ]�oρϓϥϷ�F��� �����#�5���Y�k� }ߏߡ߳���T����� ��1�C���g�y�� �����P�����	�� -�?�Q���u������� ����^���); M��q����� �l%7I[ ������h �/!/3/E/W/i/@� �/�/�/�/�/�/�? ?/?A?S?e?w??�? �?�?�?�?�?�?O+O =OOOaOsOO�O�O�O �O�O�O_�O'_9_K_ ]_o_�__�_�_�_�_ �_�_�_#o5oGoYoko }o�oo�o�o�o�o�o �o1CUgy� �����	�� �?�Q�c�u�����(� ��Ϗ������;��M�_�q�������~ ����~ ���ҟ���Ο�*��,�[���f����� ��ٯ�������3�� W�i�P���t���ÿ�� �ο��/�A�(�e� Lωϛ�z/�������� ��(�=�O�a�s߅� �ߩ�8��������� '��K�]�o���� 4����������#�5� ��Y�k�}�������B� ������1��U gy����P� �	-?�cu ����L��/ /)/;/M/�q/�/�/ �/�/�/Z/�/??%? 7?I?�/m??�?�?�? �?�?���?O!O3OEO WO^?{O�O�O�O�O�O �OvO__/_A_S_e_ �O�_�_�_�_�_�_r_ oo+o=oOoaosoo �o�o�o�o�o�o�o '9K]o�o�� ������#�5� G�Y�k�}������ŏ ׏������1�C�U� g�y��������ӟ� ��	���-�?�Q�c�u� �������ϯ������0���0���B�T�f�>�����t�,��˿~�� ֿ�%��I�0�m�� fϣϊ����������� !�3��W�>�{�bߟ� �ߘ��߼�����?/� A�S�e�w���� ����������=�O� a�s�����&������� ����9K]o ���4���� #�GYk}� �0����// 1/�U/g/y/�/�/�/ >/�/�/�/	??-?�/ Q?c?u?�?�?�?�?L? �?�?OO)O;O�?_O qO�O�O�O�OHO�O�O __%_7_I_ �m__ �_�_�_�_�O�_�_o !o3oEoWo�_{o�o�o �o�o�odo�o/ AS�ow���� ��r��+�=�O� a����������͏ߏ n���'�9�K�]�o� ��������ɟ۟�|� �#�5�G�Y�k����� ����ůׯ������ 1�C�U�g�y������ ��ӿ������-�?ϠQ�c�uχ�^P��}�^P�����@���ͮ���
���,�� ;���_�F߃ߕ�|߹� �����������7�I� 0�m�T������� �����!��E�,�i� {�Z_������������ �/ASew� ������ +=Oas�� ����//�9/ K/]/o/�/�/"/�/�/ �/�/�/?�/5?G?Y? k?}?�?�?0?�?�?�? �?OO�?COUOgOyO �O�O,O�O�O�O�O	_ _-_�OQ_c_u_�_�_ �_:_�_�_�_oo)o �_Mo_oqo�o�o�o�o ���o�o%7>o [m����V ���!�3�E��i� {�������ÏR���� ��/�A�S��w��� ������џ`����� +�=�O�ޟs������� ��ͯ߯n���'�9� K�]�쯁�������ɿ ۿj����#�5�G�Y� k����ϡϳ������� x���1�C�U�g��� �ߝ߯����������`�����`���"�4�F��h�z�T�,f���^������ ���)��M�_�F��� j����������� ��7[B�x �����o!3 EWixߍ��� ����///A/S/ e/w//�/�/�/�/�/ �/�/?+?=?O?a?s? �??�?�?�?�?�?O �?'O9OKO]OoO�OO �O�O�O�O�O�O_�O 5_G_Y_k_}_�__�_ �_�_�_�_o�_1oCo Uogoyo�o�o,o�o�o �o�o	�o?Qc u��(���� ��)� M�_�q��� �����ˏݏ��� %�7�Ə[�m������ ��D�ٟ����!�3� W�i�{�������ï R������/�A�Я e�w���������N�� ����+�=�O�޿s� �ϗϩϻ���\���� �'�9�K���o߁ߓ� �߷�����j����#� 5�G�Y���}���� ����f�����1�C�hU�g�>�i��>������������������,�� ?&cu\��� ����)M 4q�j���� �/�%//I/[/:� /�/�/�/�/�/���/ ?!?3?E?W?i?�/�? �?�?�?�?�?v?OO /OAOSOeO�?�O�O�O �O�O�O�O�O_+_=_ O_a_s__�_�_�_�_ �_�_�_o'o9oKo]o oo�oo�o�o�o�o�o �o�o#5GYk} ������� �1�C�U�g�y���� ����ӏ���	���-� ?�Q�c�u�����p/�� ϟ�����;�M� _�q�������6�˯ݯ ���%���I�[�m� �����2�ǿٿ��� �!�3�¿W�i�{ύ� �ϱ�@��������� /߾�S�e�w߉ߛ߭� ��N�������+�=� ��a�s�����J� ������'�9�K��� o�����������X��� ��#5G��k}@����������������&�HZ4, F/�>/����� 	/�-/?/&/c/J/�/ �/�/�/�/�/�/�/? �/;?"?_?q?X?�?|? �?�?���?OO%O7O IOXmOO�O�O�O�O �OhO�O_!_3_E_W_ �O{_�_�_�_�_�_d_ �_oo/oAoSoeo�_ �o�o�o�o�o�oro +=Oa�o�� �������'� 9�K�]�o�������� ɏۏ�|��#�5�G� Y�k�}������şן ������1�C�U�g� y��������ӯ��� 	��?-�?�Q�c�u��� ������Ͽ���� ��;�M�_�qσϕ�$� ���������ߢ�7� I�[�m�ߑߣ�2��� �������!��E�W� i�{���.������� ����/���S�e�w� ������<������� +��Oas�� ��J��' 9�]o���� F���/#/5/G/��$UI_INU�SER  ����h!��  H/L/_M�ENHIST 1�yh%  �( u ���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1�/�/??0?�)�/�/13�/|?�?�?$�?�'E?W>2k?�?�O"O4O��/�?148,29O�O�O�O�O�?]O,71�?__�+_=_�+�O_Eed�it�"TELEOAP�O�_�_�_B_��_ �_�_o o2oDo�_ho@zo�o�o�o�o��\a �!\o�o/AS Vow�����` ���+�=�O��� ��������͏ߏn�� �'�9�K�]�쏁��� ����ɟ۟j�|��#� 5�G�Y�k��������� ůׯ��o�o�1�C� U�g�y�|�������ӿ ������-�?�Q�c� uχ�ϫϽ������� ߔ�)�;�M�_�q߃� ߧ߹��������� ��7�I�[�m��� � �������������� E�W�i�{��������� ��������AS ew���<�� �+�Oas ���8���/ /'/9/�]/o/�/�/ �/�/F/�/�/�/?#? 5? �2�k?}?�?�?�? �?�/�?�?OO1OCO �?�?yO�O�O�O�O�O bO�O	__-_?_Q_�O u_�_�_�_�_�_^_p_ oo)o;oMo_o�_�o �o�o�o�o�olo�%7I[F?��$�UI_PANED�ATA 1{�����q � 	�}  f�rh/cgtp/�flexdev.�stm?_wid�th=0&_height=10�p��pice=TP&�_lines=1�5&_colum�ns=4�pfon�t=24&_pa�ge=whole��pmI6)  rim�9�  �pP�b� t������������Ǐ ��(�:�!�^�E��� ��{�����ܟ�՟��I6� �  �   }�J�O�a�s������� ��ͯ@����'�9� K���o���h�����ɿ ۿ¿���#�5��Y�@@�}Ϗ�vϳ�&��� �s�����)�;�M� ��q�䯕ߧ߹����� ��V��%��I�0�m� �f���������� ��!��E�W����ύ� ����������:�~� /ASew�� ���� = $asZ�~�� ��d�v�'/9/K/]/ o/�/��/�/*�/�/ �/?#?5?�/Y?@?}? �?v?�?�?�?�?�?O �?1OCO*OgONO�O� /�/�O�O�O	__-_ �OQ_�/u_�_�_�_�_ �_6_�_o�_)ooMo _oFo�ojo�o�o�o�o �o�o%7�O�Om �����^_ �!�3�E�W�i�{�� ����Ï�������� �A�S�:�w�^����� ��џDV��+�=� O�a�������
���ͯ ߯���|�9� �]� o�V���z���ɿ��� Կ�#�
�G�.�k�ޟ�}�|ϵ����������)��4ߧ�#�`� r߄ߖߨߺ�!����� �����8��\�C�� ��y������������������$UI_�POSTYPE � ���� 	 �s�B�Q�UICKMEN � Q�`�v�D�R�ESTORE 1�|��  O������������mASe w�,����� �+=Oan �����// �9/K/]/o/�/�/6/ �/�/�/�/�/�?? 0?�/k?}?�?�?�?V? �?�?�?OO�?COUO gOyO�O6?@O�O�O.O �O	__-_?_Q_�Ou_ �_�_�_�_`_�_�_o o)o�O6oHoZo�_�o �o�o�o�o�o% 7I[�o�������SCRE��?���u1s]c��u2�3�U4�5�6�7��8��sTATM��� ����:�USE�R�p��rT�p�k�s���4��5��6ʝ�7��8��B�ND�O_CFG }�Q�����B�PDE����Non�e��v�_INFOW 2~��)���0%�D���2�s�V� ������͟ߟ�� '�9��]�o�R���z���OFFSET �Q�-���hs�� p�����G�>�P� }�t���Я��׿ο� ���C�:�L�^Ϩ����͘���
����av���WORK �!�����.�@ߢ��u�UFRAME � ���RTO?L_ABRT���Ω�ENB�ߣ�GR�P 1�����Cz  A���� ��*�<�N�`�r��ĥ֐�U�����MS�K  �)���N6��%!��%z�����_EVN������+�ׂ3�«
 }h�UEV���!td:\ev�ent_user\�u�C7z���jpYF��n�SPs�x��spotweld��!C6��������!���G|' ��5kY���� �>���1 �Ug���/� �	/^/M/�/-/?/�/ c/�/�/�/�/$?�/H?h�/:J�W�3���F��8C?�?�? �? �?�?�?O+OOOOaO <O�O�OrO�O�O�O�O _�O'_9__]_o_J_��_�_�_�$VAL�D_CPC 2�« �_�_� w��qd�R�*oP_oqo��hsNbd�j �`��i�da{�oav�_ �ooo3BoWi{ �o�o�o�o��o� PA�0�e�w��� �������(� =�L�a�s�
������� ʏ�����$�ޟH� :�o���������ڟ؟ ����� �2�G�V�k� }�������¯ԯ��� ��.��R�S�yϋ� �����������	�� *�<�Q�`�u߇ߖϨ� ����������&�8� M�\�q���߶��� n������"�4�F�[� j������������� ���!0�B�Wf�{ ����������� ,>teT�� �����/+/ :La/p�/�/./� ����//'?6/H/ ?l/^?�?�?�/�/�/ �/�/?#O�?D?V?kO z?�O�O�?�?�?�?�? _O1_@ORO9_vOw_ �_�_�O�O�O_�__ -o<_N_`_uo�_�o�o �_�_�_�_o&o; Jo\oq�o����o �o�o� �"7�FX j��������� ��!�0�E�T�f�{� ������ßҏ���� 
�,�A�P�b�����x� ����Ο�����(� *�O�^�p��������� R�ܯ� ��Ϳ6�K� Z�l�&ϐ��Ϸ���ؿ ���"� �2�G���h� zϏߞϳ��������� 
��1�@�U�d�v�]� �ߛ����������,� �<�Q�`�r����� ����������&�; J�_n�������� ������$F[ j|������ �0E/Ti/x ��/��/�/�/�/ /,/.?P/e?t/�/�/ �?�?�?�?�/??(? :?L?NOsO�?�?�O�? �O�OvO OO$O6O�O ZOo_~O�OJ_�O�_�_��_�O_ _F_D_V[��$VARS_CO�NFIG ���Pxa � FP]S�\lC�MR_GRP 2��xk ha	�`�`  %1:� SC130EFG2 *�o�`]T�VU��P�h`�5_P~a?�  A@%pup*`�Vn No9xCVXdv��a8��<uA�%p�q��_R��_R B���#�_Q'� �H��l�;���{��� ��؏ÏՏ�e��D��/�A�z�-�����ddI�A_WORK ��xeܐ�Pf,�		�Qxe���G��P ���YǑR�TSYNCSET�  xi�xa-�W�INURL ?=�`����������ȯگSIONOTMOU9�]Sd�� ��_CFG� �S۳�S�۵P�` �FR:\��\DA�TA\� ��� MC3�LOG�@�   UD1�3�EXd�_Q' B@ �����x�e_ſx�ɿ�VW� � n6  ���VV��l��q  =����?�]T<�y�Y�TR�AIN���N� 
�gp?�CȞ��T�K���b�xk ( g�����_�������� �U�C�y�g߁ߋߝ�p�������_GE�ݑxk�`_P�
��P�RꋰRE���xe*�`hLEX��xl`1-e�VM�PHASE  �xec�ecRTD�_FILTER �2�xk �u� 0����0�B�T�f� x�����VW��������  $6HZl_i�SHIFTMEN�U 1�xk
 <��\%������ ����=& sJ\��������'/�	LI�VE/SNA�c%vsfliv��9/��� 7�U<�`\"menur/w/@/�/�/�����]�V�MO��y��5`�h`ZD4�V�_Q<���0��$WAIT?DINEND��a|2p6OK  �iȋ<���?S�?�9TI]M�����<Gw? M�?*K�?
J�?
J�?�8RELE��:G6�p3���r1_ACT�O 9Hܑ�8_<� �ԙ�%�/:_af�B�RDIS�`�N�o$XVR��y��$ZABC�b1��S; ,��j��I�2B_ZmI1�@VSPT �y��eG�
�*�/o�*�!o7o�WDCSCHG �ԛ(��P\g�@�PIPL2�S?i��o�o�o�Z�MPCF_G 1	��ii�0'¯S;M�s�S��i��p'���g��e2�� �Z� ����	=������곿�  ��Z�q�5�g���pD5�8o�G��C��]I�1�q>;��>y��m��B<H�
�����N��� ����+�Z�~����Ï�>��3�����n����b ڏ�ӈ*���*�@�@N�x��$�6�H�0N��`��Tp���o�_�CYLIND��� { Х� ,(  *=�N�G�:�0w�^����� ��ѯ ���7����<�#�5� r�����������޿y� _����8�ύ�nπ��㜻ã wQ � 5�����S�����(��ٻ�X�זr�A���SPHERE 2���ҿ��"ϧ� �����P�c�>�P�̿ t���ߪ�����'� ��]�o�L���p�W��i������������PZZ�F �6