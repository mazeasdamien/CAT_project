��   8��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����DCSS_I�OC_T   �P $OPER�ATION  $L_TYPB7IDXBR1H[ �S2]2R��$�$CLASS  �������Pz��P� VERS?��  �XK�IRTUAqL��' 2 ��P @ �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt����������_C_CCL ?���  	All param���
Base!��Pos./Sp�eed chec�kF�Safe I�/O connect�}R��,�>�XP�b�t�SI��@���� �,�>�g�b� t���������Ο��� ��?�:�L�^����� ����ϯʯܯ��� $�6�_�Z�l�~����� ��ƿ�����7�2� D�V��zόϞ����� �����
��.�W�R� d�vߟߚ߬߾����� ���/�*�<�N�w�r� ������������O����C�l�g�y� ��������������	 D?Qc��� �����) ;d_q���� ���//</7/I/ [/�//�/�/�/�/�/ �/??!?3?\?W?i? {?�?�?�?�?�?�?�? O4O/OAOSO|OwO�O �O�O�O�O�O__�}N�  7�_b_�_ �_�_�_�_�_�_�_o o(o:oco^opo�o�o �o�o�o�o�o ; 6HZ�~��� ����� �+_�SI��6�7������� ��ȏ�����9�4� F�X���|�����ɟğ ֟����0�Y�T� f�x����������� ���1�,�>�P�y�t� ��������ο�	�� �(�Q�L�^�pϙϔ� �ϸ������� �)�$� 6�H�q�l�~ߐ߹ߴ� �������� �I�D��O�PC_�u�SF'DI1N��2���I3���4���5��6���7���8 -�`�Q�c�u������� ��������); M_q����� ��%7I[ m������ �/!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy� ������	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q���������˟ ݟ���%�7�I�[�$f�x�O���O�ﵣ �ﵣ�ﵣ�ﵣ�ﵣ ���,���D�~�o��� ������ɿ����� :�5�G�Yς�}Ϗϡ� �����������1� Z�U�g�yߢߝ߯��� ������	�2�-�?�Q� z�u���������� 
���)�R�M�_�q� �������������� *%7Irm� �����! JEWi���� ����"////A/ j/e/w/�/�/�/�/�/ �/�/??B?=?O?a? �?�?�?�?�?�?�?�? OO'O9ObO]OoO�O �O�O�O�O�O�O�O_ :_5_G_Y_�_}_�_�_ �_�_�_�_ooo1o�ZoUogoyo�o��SIz����VOFF�o�FENCE�oEXEMG�o�os�NTED"�OP2qAUTO:T��ysӯq�MCC�3pCS�BP�
POSSPD_ENBz�CONF_OK��~F_IPAR_�CR�z�g�������o�q_�oY�p�E�DIS�|C_6�r_~��� 