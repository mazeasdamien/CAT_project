��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1�TU4QQ���AR�x1R� � /$TIT91� �� � �Td�T0�ThP�TU5�V6�V7�V8�V9�W0�W�WOQ�U�W�gQ�U�W1�W1�W1��W1�W2�R�SBoN_CF�!@$<!J� ; ;2�1�_CMNT�$�FLAGS]�C�HEK"$�b_O�PTJB � ELL�SETUP � `@HO8@9 P�R�1%�c#�aREPR�hu0D+�@���b{uHM9 MN�B;16 UTOB�J U�0 }49DEVIC�STI/@�� �@b3�4pB�d�"VAL��#ISP_UNI�tp_DOcv7�yFR_F�@|%u13���A0s�C_WAx�t,q�zOFF_T@]N�DEL�Lw0pdq�1�Vr?^q��#S?�o`Q"U��t#*�QTB��bMyO� �E � �[M�����RE�V�BIL���!X�I� v�R  �!D�`��$NOc`M�|����ɂ/#ǆ� �ԅ��ނ�@Ded �p E RD_E���h�$FSSB�6�`KBD_SEV�uAG� G�2Q"!_��2b�� V!�k5�p`(��C�00q_ED|� � � t2d�$!S�p-D%$� ��#�B�ʀ_�OK1��0] P_C�� ʑ0t��U �`LACI�!�a�Y�� ��qCOMM� # $D
� ��@���J_�\R BIGALL;OW� (Ku2:-B�@VAR���!|�AB   �BL�@� � ,K�q��r�`S�p�@M_O]�˥��CCFS'_UT��0 "�A�Cp'��+pXG��b�0� 4� IMCM ��#S�p�9���i �_�"t\b���M�1 h$�IMPEE_F�s���s��� t����D_(�����D��F��� �_����0 aT@L��L�DI�xs@G�� �P�$I�'�����CFed XF@GRU@��Mb��NFLI�\Ì@U�IRE�i42� SgWITn$`0_N�`�S 2CF�0M�' �#u�D��!���v`����`J�tV��[ E��.p�`��>�ELBOF� � շ�p`0���3����� F�2T��A`��rq1J1��z _To!��p��g����G� �r0WARNM�p#tC�v`�ø�` � COR-�UrFLTR��TR�AT9 T%p� $ACCVq��� ��r$ORI�_&��RT��S<��HG*�0I���TW��A��I'�T���H9K�� �2028�a1��HDR�2��2�2J; S���3���4��5��6��7
��8��9��׀
 �2� @� TRQB�$vf��'�1�<�c_U<�G� COec  <� P�b�t�x53>B_�LLEC��}!~�MULTI�4��"u�Q;2�CHI�LD��;1ذO�@T�� "'�STY 92	r��=��)2��������ec# |@r056$J ђ��`����uTO���E^	EXTt����2��22"����$`@D	�`&��p������(p�"��`% �ak�����s�����A&'�E�Au��Mw��9 �% ��TR>�� ' L@�U#9 ���At�$J�OB����P��}IG��( dp��� ���^'#j�~�L��pOR�) tf$�FL�
RNG%Q@�TBAΰ �v&r� *`1t(��0 �x!�0«+P�p�%4��*��͐U��q�!�;2MJ�_R��>�C<QJ�8&<J D`5CF9���x"�@J���P_p�7p+ \�@RO"pF�0��I9T�s�0NOM��>Ҡ�4s�2�� @U<PPTgў�P8,|Pn�ć0�P�9�͗ RA����l�?C�� �
$�TͰtMD3�0TD��pU�`�΀+AYHlr>�T1�JE�1 \�J���PQ��\Q��hQ�CYNT�P��PD'BGD̰�0-���PU6$$Po�|�u��AX����TAI�sBUF,�O!�A�1�. ����F�`PIV|�-@PvWMuX�M�Y�@�VFvWSI�MQSTO�q$7KEE�SPA��  @?B�B>C�B�2��/�`=��MARG�u2��FACq�>�SLEW*1!0����
�4ذs�CW$0'����pJB�Ї�qDE�Cj�e��s�V%w1 Ħ�CHNR�;MPs�$G_@�g�D�_�@s��1_FP�5�@TC�fFӓC@�Й���qC��+�VK��*��"*�JRx���SoEGFR$`IOh!v�0STN�LIN>�csPVZ�z�Ц@�D2����r 2��hr�r��1��3` + ^?���եq�`��q|`������t��|aSI!Z#�!� �T�_@%�I��qRS�*s���2y{�Ip{�pTpLpF�@�`��CRC����CCTѲ�Ipڈ�a8���bL�MIN��aP1순���D<iC �C/���!uc�OP4�n �j�EVj���F��_
!uF��N����|a�֔=h?KNLA�C=2�AVSCA�@�A�WQ�a�4�  cSF�$�;�Ir�Kঠ'��05��	 D-Oo%g��,,m�����ޟ��RC�6� n���sυ��U��R�0HANC���$LG��ɑDQ�$t�NDɖ��AR۰N��aqg��ѫ�X��ME��^�Y�[PS�RAg�X�AZ�П���:rEOB�FCT��A���`�2t!Sh`0ADI��O��y�s"y�n!@�������~#C�G3�t!��BMPmt@�Y8�3�afAES$���v��W_;�BAS#?XYZWPR��*��m!��	y�U�87/  ƀI@d��2�8\�p_C:T����#��_L
 � 9K ���C�/�(z�J�LB�$�3�xD��5�FORC��b�_AV;�MOM$*�q�SaԫBP`Ր� y�HBP�ɀE�F�����AYLOAD&$�ER�t&3�2�X�rp�!ҁ�QR_FD��� : T`IH�Y3��E�&��Ct���MS�PU
$0(kpD��9 �b��;�B�	EVId�y
�!_IDXY�$���B@X�X�<&�SY5� � �HOPe�<��AL�ARM��2W�r}rR9_�0= hb P�nq�`M\qJ@$PiL`A&�M#�$�` ��� 8�	���V�]�0�U�qU�PM{�U���>�TITu�b
%�![q�BZ_;�.��? �B pQk���6NO_HEADE^az��}ѯ��`� �����dF�ق�tc`����@�@��uCIGRTR�`��ڈL���D�CB@4�RJ�� 1�[Q���A�2>�&��OR�r��O����T`UN_OO�Ҁ�$����T������I�VaCnp�DBP�XWOY���B��$SKADR��DB]T�TRL��C���րfpbDs��~�DIJj4 _�DQ}���PL�qwbWA���WcD�A��A�=�2�UMMY�9��10�VIȾ ����D;[QPR�� 
M�Z���gE O�Y1$�a{$8��L)�F!/��
����0G�G/��9�PC�1H�f/3#PENEA@T�f�I�/���RE�COR`"JH y@ �E$L�#F$#PR���+jp���nq�_D$�qPROSS]�
���R�r�` >u�$TRIG96�PAUS73ltETgURN72�MR:�eU 0Ł0EW$�~�SIGNALA��QR$LA�З5�1�G$PD�H$PDİ�AI�0�A�C�4�C��DO�D�2�!��6GO_AWA�Y2MOZq�Z��,CS��CSCB�g�K Իa#���E+RI�0Nn�T�`$�����FCBPL�@QBGAGE���P��ED`|BD�wA[CD�OF�q�[F0�FoC��MPM�AB0XoC�$FRCIN��2Dk��@��O$NE�@�FD�L8�� L� �����=��Rw�_��P>� OVR10����lҠ�$ESC_|�`uDSBIO��p��pTe�E�VIB�� `s��Z��V��p�SSW��$�VLY�:�Lk��X���ѣ�0bQ����USC�P��qA=�	Q��MP1%e@&S*`�(bt`'c5۳ESUd��-cWg&S Wg?cWd����Wd��Wd<.���AUTO$�Ya҃�ac�SB����-d���&SwB[��GB�f_$VOLT�g ���  �GAOD!��q���@:�ORQ�ҀKra�$DH_THE&0�Rgp� <qtnwALPHnt��o��w0 Vp]�$�.�Ra�[��s�5�`r�CQ�#BUD�S� F1M���sV
��;��L�b�tk���BRTHR��L��T`�Z���Vɖ��D)E  �1��2�⋅ ��������kѯ�a� �Tt0V�ꆸ������@̈Я�-�"�N~���sS2����INHB��ILTG0ɡ�T?� �3$�w��E��PqQxQ��TqPe��0Y�AF}�O�ນ��ڗ ��qPڳē����bPܙ���PL?���3���TMOU��ēS��� � ��s�/�S18���O��Aܙ��I����CDqIƑ˩o�STI��գ�O:ҋ�,0���AN��Qg�S��+r�#x$�����w�1_����PRA�P`�vC����MCN�eQe�����VER�S��r�oPIw�F�PåǲШ۷G.�DEN��G>�����F�2H�Ƿ�M�7�F��_�MN�D̠,���@�d�{ƭa����OB����U˱z���DI ���#���3�����A��w�Fx���3�O�N�5��Q��VAL��CR[�_SIZp��b�;Qn�REQ�R�b��]2b���CH q�΂�ڃ�Ռ�����:�n�S_U��X��wW�FLG���wU$CV�iMGP�QδFLXP�923R�u�L��EAL�P-�C	�F+rT��W��� �R��c���NDMS�7� ��K>S�P_M'0h�STWv������AL�P���Q����U���U�IAG@,�o��d�U�-�T"	A-`� ���A��� ��H`��Q`��6��Pq_D&��1s��.�P��F�"2�T�� ?7 1A>���#�#L��?`_=i @@>LD�pc�F�0�FRI�0 `Ѐ��1}Ѳ�IV\1�*�^1�U�P`��a��C�L!W��
`L=S&-c&&S�C.w��  L���!����d�Q$w!�҇��$w��p��
�P�5RSM��P���V0h � r�l�d^2AW�a_TRp�}�8@NS_PE�A����< ��$�SAVG�8�6G]%���CAR �`�!�$���"CRa���$ d�#qE�@��"STD���!Fpo��'QOF0��%��"RC���&RC۠�(F�2A�R#7����%, gMA�Q_�a��
QQ��al2��%u4Ib�r7I�R�9�wQ�7�8M/��!C:pR�  �p�2F<�SDN�a0 � W2QM P $Mi��s$cA �$C�cm�9���4���AT�0CY_ �N LS!IG1@x'yB��y@@H2Y��NO����SDE�VI�@ O@�$�RBT:VSP0�3�CuT�DBY|�A�	W`3CHNDGD�AP H@GRP�HE iXL�U��VSЌFx2� DL1p aQ6ROp��FB�\]�FEN�@��S���ChAR d�@DyOd�PMCSb���P薇P�R��HOT�SWz42�DMpEL�E�1/ex\8`�RS T�@���r� hf��`OL�GHA�Fk�Fs�����C�A@�T � $MD�LUb 2S@�E ���q�6�q	0�i�c�e
�cJ��	uݢ�#~X5t+w�PTO��� x�byU DSLAVS�� U  ��INAP �	V�ЊyA_;�wENUAV $R��PC_�q�2 1bLp�wpp B�pSHO+� W ���A�a�qB�2�r�v�u�v�b�_CF� X�` ,f��r�OG� gE��%D�h��p2C�Iߣi�MA��D��x AY?�W� p�N3TV	�D�VE�0@�SKI��T�`g?Ň2�� JZs�! �Cꆻ��f�_SV</ �`XCLU��H����ONL��'�Y��T��OT:eHI_�V,11 APPLY���HI4`;�U�_M�L�� $VR�FY8�	�U�M{IGOC_I���J 1/d��߃O�@X�LSw"�`@$DUMMY�4���ڑ�Cd L_TP���kC��^1CNFf���E��@HT�y� D_#UQ_��ݥ�YPCP��=�� ������uJ �ҟ Y +�
0R�T_;P��uNO�CCb Z�r�TAE���=�פ�DG��@[ D�P_B�Ae`kc�!I��_��H�t~T��E \�pyAb=cARGI�!�$���`[��SGNA] ��`U���IGN�Տ��� ���V������ANNUN��&�˳�EU�<J'�ATCH���J��B��u^ <`@g�����:c$Va������ᑴaE�F] I�� _ �@@FͲITb�	$TOTi �C�O��c� @EM�@NIF�a`tB��c��ùA>���DAY@CLOAD�D\�n���� �EF7�X�I�Ra��K���O�%��a�ADJ_)R�!@b��>�H2��"[�
 c�%��`a�͠MPI�J��D��qA��?�Ac 0� �х�� ��Z�ϡ��Ui ��CTRLܖ Yp d��TR�A8 ?3IDLE_�PW  �Ѡ��Q��V��GV_���`c ��o�;Q@e� �1$��6`<cTAC�-3��P�LQ�Z�Rdz\ A-u:ɰSW;�A\���/Jղ�`b�K�OH�(OsPP; �#IRO� ��"BRK��#AB  �������� _ ���F���`d͠, j@�S�RQDW��MS��P6X�'z��IF�ECAL�� 10^tN��V��豊�V�(0}f�CP
��Nr� Yb�0FLA_#f�OVL ��HE��>�"SUPPO��ޑ�\�L�p��&2XT�$Y-
Z-
W-
���/��0GR�XZl�q�$Y2�CO�PJ�SA�X2R��*r�!���:��"�rI�0)��f `�@CACH�E��c��0�s0L}AZ SUFFI, C��q\��哹6��QMSW�g� 8�KEYIM[AG#TM�@S���n
2j�r���ROC�VIE��~�h ��aBGL����`�?G� 	Q���i��m!`STπ!� �����n����/EMAI�`N��`A��`Z�FAU� �jH�"�qa��U�3�qq� }�k< �$I#�US�� �IT'�BUF`�r�DNB���SUBu$��DC_���J"��"SAV�%�"k�������';��P�$�UOR	D��UP_u �%��8OTT��_B`��8@�LMl�F4��C7AX�@Cv���Xu 	��#_uG��
 @YN_��R�l6���D�E��UM����T��F���caC�DI`BED%T)@C��~�m�rI��G�!c�&��l`���-�P��FZP n (�pSV� )d\��ρ���2ΰ��o�� ����>"$3C_R�IK��kB���hD{pRfgE.(AD�SP~KBP�`�II�M�#�C�Aa�A��UЂG���iCM! IP`��KC��� �DTH� ȷS�B*�T��CHS�3�CBSC��� ���V�dYVSP�#[T_D^rcCONV�Grc�[T� �Fu F�ቐd0�C�0j1��SC5�e�]CMER;dAFBgCMP;c@ETBc� p\FU D�Ui ��+�~�CAD�I%P702#@O��B�qWӏ�SQ��QǀSU��MSS�1ju�4`��TB�Aa��A�1r�� "�Й��4�$ZO@s���l�U�6�&��eP���eCN�c�l��l�l�iGRO�U�W)��S c�MN�kNu�eNu�eNpR|b|�i�cH�pi��z
 �0CYC���s�w�c���zDEL�_D��RO�a���qVf���v{�O�2���1���t��:R�ua�.#�� ���AL� �1s@ˢI1¡�J0�PB��,렒�ER^�T�Gbt ,!@��5��aGzI1LcR1s 
�0&ԠNO��1u����H�����P����Cڠ	�����!���J0��0vH *	�L U�1#J�Q��V
�[�7A z���z��z�n�z�Ѩz�Fz�7w�8w�9Pw���y���1��1��U1��1��1Ě1њU1ޚ1�2��2�����2��2��2��2�Ě2њ2ޚ2�3J��3��3����3��U3��3Ě3њ3ޚ�3�4���EXTF��1w6�.(�0�f�0��U�0ŷ�e.�FD�R5�xTU V�E��?1���SR��R�E�F���OVM�~C)�A2�TROVf2�DT� R�MXa��IN2���Q�2�IN	Dp�r�
���0�0�0�Gu1��[�G`��{�D_�[�RIV�P��oGEAR~AIOr�	K"N�0�y�p��5`@�a�Z_MC�M� ���F��U�R�Ryǀ��!?3 ��p?nЋ�?n�ER�v�Gme��!�P��zIj:�PXqB�RI0%�>`�#ETUP2_� { ���#TDPR�%TBp�������K�"BAC�2| QT��"�4)�:%	`t^B��p�IFI���� Mc���.�PT|��I �FLUI��} � ��K UR�c!���B�1SPx NE�EMP�p�2$��]S^�?x��Jق�0
3VRT���0x/$SHO��Lq�6 ASScP=1��PӴBG_�������FORC�3" �i�d~)"F%UY�1�2\�2
A�h� p� |��N�AV�a��������S!"��$VI�SI��#�SCM4S�E����:0E�V�O���$���M����$��I��@��FMR2��� �5`�r�@ �� �2�I�9 F�"��_���LIMI�T_1�dC_LM�������DGCLFl����DY�LD����5������F  ���D u	 T�sFS0Ed� P���QC�0$EX_QhQ1i0�P�aQ53�5��GoQ��g� ����RSW�%�ON�PX�EBUG���'�GRBp�@U��SBK)qO1L� ��POY 
)�(�P��M��OXta`KSM��E�"�0�����`_E � x
@F���TERMZ%9�c%�aORI�1_ Y�c%d�SMepO��B_ �|&.�`�(�c%��e:�UP>� ?�� -���b����q#� ���G<�*� ELTO��p�0�PFIrc�1Y���P�$�$�$UFR�$��1L0e&� OTY7�PT4q��k3NST�pPATz�q4PTHJ�a�`EG`*C�p1AR�T� !5� y2$2R�EL�:)ASHFTPR1�1�8_��R�P�c�& � $�'@�@� ��s�1 @I�0�U�R G�PAY�LO�@�qDYN_�k���.b�1|��'PERV��RA��H��g7��p�2�J�E-�J�R�C���ASYMFgLTR�1WJ*7����E�ӱ1�I��aUT�pbA�5�F�5aP�PlC�Q1FOR�p�M��GRI!����W��/&�0F0�a H��Ed� �m2N���5`OC1!?�$OP����c��c���bRE�P�R.3�1a�F��3e���R�5e�X�1(�e$PWR��_���@�R_�S�4��et$3U�D��.�Q72 ����$H'�!�`AWDDR�fHL!G�2(�a�a�aT��R��U�w� H��SSC����e-��e���e��S�EE��HSCD���� $���P_"�_ B!rP����}T!HTTP_���HU�� (�OB�J��b(�$�fL�Ex3pWq�� �� ���ะ_��T�?#�rS�P��z�KRN�LgHIT܇5��P ���P�r������PL���PSS<�ҴJQUERY_FLA 1��qB_WEBSOC���HW�1U����`6PINCP	U���Oh��q�����d���d���� �I�HMI_ED� T� �RH�?$��FAV� d�Ł��wOLN
� 8��yR�@$SLiR�$INPUT_�($
`��P�� �؁SLA� ����5�1��C���B��IO6pF_AuS7��$L%�}w%�A��\b.1��0���T@HYķ������Qh�UOP4� `y�ґ�f�¤�������`PCC
`���#���aIP_M�E�񵁗 Xy�I�P�`�U�_NET�9���Rĳs�)��DSP(�Op=��BG�����M��A��� lp:CTiAjB�pAF TI�`-U��Y ޥ�0PSݦBUY IDI�rF ���P�q�� �y0��,����Ҥ�N�Q�Y R��IRCA|�i� � ěym0�CY�`EA������񘼀�CC����R�0�A�7QDAY_<���NTVA�����$��5 ���SCA�d@��CL���� ���𵁛8�Y��2,e�o�N_�PCP�q��ⱶ��,�N�����
�xr���:p�N� �2��Ы�(ᵁ�p���xr۠LABy1���Y ��UNIR��Ë ITY듭��e�ւR#�5���R�_URL���$AL0 EN��ҭ� �;�T��T_U��A�BKY_z��2DI�SԐ�kSJg�����P�$���E��g�R���З A�/���J����FLs��7 Ȁ|���
�UJR� ���F{0G��E7��J7 O^ R$J8I�7�H�R�d�7��E�8{��H�APHIQ�S��DeJ7J8�B��L_KE*� � �K��LM�[� � <X�X�Rl�u���WATCH_VA��o@D�tvOFIELc��cy��L��4� � o1Vx@��-�CT[�9�m�� ��LGH���� $��LG_SIZ�t�z�2y�p�y�FD��Ix���+!�� w�\ ����v��S��� 2��p�������\ ��h�A�0_gCM]3NzU
RFQ\v�v�d(u�"B ��2�p����I��+ �\ ��fv�RS���0  ��ZIPDUƣp�L)N=��ސ�p��z6���f�>sD�PL�MCDAUiEA`Fp���TuGH�R�.OGBOO�a��� C��I�IaT+���`��RE����SCR� �s��D�I��SF0�`RGIO"$D�����T("$�t|�S�s{�W$|��X��JGM^'MN3CH;�|�FN��a&1K�'uЅ)UF�(1@n�(FWD�(HL�)STP�*V�(%Г(,��(RS9HIP�+��C[T�# R��&p:'^9U=q�$9'�H%C�d���"Gw)�0PO�7��*��#W}$���)E]X��TUI�%I�� �Ï���rCO#C� N*�$S��	)���B@�NOFAN1A|��Q
�AI|�t:��EDCS��c�CT�c�BO�HO�GS����B�HS�H(IGN������!O���DDEV<7LL�ѩ�|��­Ц(�;�T��$��2�p������#A
���(�`�{�Y���POS1�U2�U3��Q	��2�@�Ш ��{�PtD�����&q)��0�d��VST�ӐR�Y��B@ ` _�$E.fC.k��p<p=fPf���4�ѩ LRТ� ��x�c �p��<�Fp�d��?"�/_ �����Kqx&���c �MC7�� ���CLD�PӐ��TRQLI0#ѽ�ytFL��,r��5s8�D�5wS�LqD5ut5uORG���91HrCRESERAV���t���t���c~�� � 	u095t5u��PTp���	xq�t�vRCLMC�������q�q�M��k�������$DEBUGMA�S��ް��?U8$T�@��Ee�g���MF�RQՔ� � �j�HRS_RU�7��a��A��k5FgREQ� �$/@x�OVER��n�t�V#�P�!EFI�%�a��g��d���tǯ \R�ԁd�$9U�P��?A��SPS�P��	߃C���͢a��U\�l��?( 	�MI;SC� d@�QkRQ��	��TB �� Ȗ0A՘AX����ؗ�EXCE�SjҔЪ�M��\���W����ԝ���SC>�P � H��̔�_��Ƙǰ]���
�MKHԳK�J� �m�B_K�FLIC��dB�QUIREG3MO��O˫3���ML�`MGմ @�`��T���a#NDU�]��>���k�G�Df��INAsUT���RSM>�a��@N�r]3-��p�5�PSTL\�� �4X�LOC�VRI�%��UEXɶANG�uBu�R�ODA��ŷ�������MF O����Y�b@�e4Ŝ2k�SUP�e��F�X��IGG� � �A��c���c Q6�dD�%�b|�!`�Ȁ!`��|��3w�ZWa�T!I��p�a M��[��� t��MD��I��)֟@���H8ݰM��DIA��ӂ��W,!�wQ�1�D��)��O���]��[ 0�CU��VPА�p���!_V��ѻ� ��P�S�X�5�	�����P��0N��ЍP��KES2���-�$B� ����ND2x����2_TX�d�XTRA�C?�/��qM�|q�`�Pv�`�XҰ�Pt SBq`^�USWCS��T��<	���PULS��A��NSޔ��R��JOIN��H��~`j�=��b��b�����P�=��$��b$���TA����S���S�HS�ME��SCF�aPJ���R��PLQ� 
M��LO��н.�L��^����8��Ҹ����0�RR2���O 1��eA�q/ d$��Iΐ+��G�A2+/� ;�PRIN�w<$R SW0"��a/�ABC�D_�J%�¡u��_J3:�
�1SPܠe�u�P��3��р`
u��J/���r�q�O8QIF��CSKAP"z{�{�J���QL2LBҰ�_AZ�r�~ELxQ��OCMP���T���RT�����c1�+���P1��t>@�Z�SMG0���=�JG�`SCL<�͵SPH_�@���%V�u� RT�ER`  �< A_�@G1"�A�@c���\$DI�
"23U�DF�}!LWn�(VELqIN�b)@� _BL�@u��$ G�q�$�'�'�%`<��� ECHZR/�TS�A_`����E�}`<����5�Bu�Ht1}`_�� �)5 D2d%��A4I��N9t&FR�DH�A���ÀP�$V `�#>Aa$��Ͳ�$Q���R}ӆ��H? �$BELvᵆ><!_ACCE�!c�x�7/��0IRC_] ���pNTT��S'$PS�rL�d� /Es��F{�@F
��9gGCgG36B���_�Q�2�@�A���17_MGăDD�A]"ͲFW�`���3�EC��2�HDE�KPPA�BN>G��SPEE �B�Q%_pB�QY�Y�|�11$USE_��,`Pk�CTReTYhP�0�q P�YN��AAe�V)хQM����ѷ��@O� YA�TINCo�ڱ�B�DՒ�WG֑ENC����u��.A�2Ӕ+@INPO�Q�I6Be��$NT|�#�%NT23_�"ͲIcLO� Ͳ_`��I�_�if� _�k�? ȼ` ej�C400fMOSI�A���ОA䃔�PERCH  �c��B" �g��c��lb =�����oUu@�@		A6B(uLeT	~��1eT�ljgv�fTRK@%�AY��"sY��q 6B�u�s۰�]��RU��MOMq�ՒY�MP�^��C�s�CJR���DUF �BS_BCKLSH_C6B )����f���St�H��R�R��QDCLALM�-d���pm0��CHK����GLRTY ���d��Y��)Üd'_UM]�ԉC��A�!�=PLMT� _AL�0��9��E� .� ��#E)�#H� =�0�Q3po�xPC�ax�HW�頿EׅCMC�E��@�GCN_,N�D�Ζ�SF�1�iV oR��g<!��0r���7CATގSH)�, �DfY��f��7A����܀PAބ�R_P݅�s_ �v��X�s����JG�T]��Y�����TORQ�UaP��c�yPOU`��b��P%�_W�u �t��1D��3C��3C�UIK�IY�I�3F�`6�����@VC�00RQ�t��1���@ӿ��ȳJRK������UpDB M��UpM�C� DL�1BrGR�VJ�Cĭ3Cĳ3$�H�_��"�j@q�COS~˱~�LN���µ �ĭ0�����u�����ē��Z���f$�MY���؊���>�TH�ET0reNK23��3hҧ3��CBm�C5B�3C! AS� ��`u��ѭ3��m�SB�3���x�GTS$=QC������������$DU��Kw�B�%(��%Qq_��a��x�{�K���b(��\сA`Չ��p�{�{�LCPH~�g�Aeg�Sµ ��������g������֚�V��V��0��UV��V��V��V��UV	�V�V%�H��@������G�����H��UH��H	�H�H%��O��O��OV	��O���O��O��O��O*	�O�O�Fg����	�����SPBA?LANCE_-��LE��H_`�SP�!1��A��A��PFULCElTl���.:1��UTO_<����T1T2��22N���29`�!�q�nL�=B�3�qTXpO�v 
A4�INSEG�2�aREV��`agDIF�uS91�8'6t"1�`OB.!t��M��w2�9`��,�L�CHWARRCBA	B�� ��#�`-ФQ 5�X�qPR��&���2�� 
�""��1neROB͠CR0r|5�����C�1�_��T � x� $WEIGH��P`$��?3àI̡Qg`IFYQ�@LA�G�Rq�S�R �RBILx5OD�p�`V2ST�0V2P!t�W0P�11�&1/0�30
�Px�2�QA  2řd^[6DEBUg3L_@z�2�MMY9&E� Nz�D`$D�_A�a$�0��O� � �DO_:@A.1� <B0�6��m�Q�B�2�0N�-cdH_p`�P��2O��� �� %"��T`"a��T/!�4�)@TICKh3| TE11@%�C ��@N͠�XC͠R?��Q�"�E��"�E8@PROMP��SE~� $I�R��Q��R;pZRMCAI)��Q�R4U_r0C2S; �q�PR8�7COD�3FU�Pd6ID_[�vU R!�G_SUFFu� �l3�Q;Q�BD�O�G �E�0�FGR r3�"�T�C�T�"�U�"��Uׁ�T8D�0�B0Hnb _FI�19*c7ORD�1 50�2�36V�+b�Q1@$�ZDT}U 1�0;E��4 *:!L_N�AmA�@�b�EDEF_I�h�b�F�d�E�2��F�4�F�c�E�e�FISP��PAKp�Ds�C�d��44בi��2�D�"�It�3D�O|#OBLOCKEz���S�O�O�Gq�R�PUM�U�b�T�c�T�e�T !r�R�s�U�c�T�d�R �6�q�S� ���U�b��U�c�S�Z��X�@P@` t�@qe�)@W�x4���s 1TE�<D��( l1LO�MB_��ɇ0V2V�IS;�ITYV2A���O�3A_FRI��a SIq�Q!R�@��@�3�3V2�W��W�4����_e��QEAS^3�Rϡ���_�[p:R�4�5��6_3ORMUL�A_Iz���TH]R^2 �Gtg�30�f��<8�5COEFF_O�A	 ��A���GR�^3Sg0BCAnO/C$��]30�1�GRP� � �G $�p�YBX�@TM~w���u�B�s��bCER, Tttsd$`7�  �LL�TSpS~�_SVNt�ߐĸ�$`�@��$`� ���SETUsMEA*P�P��W0�1+b>/0� � h��  @ڐo�l�o�cqDz��b�@cqq`t�P�G��R�� Q\p�*q[p��>�c NPR�EC>at��ASKy_$|�� PB1?1_USER�e"��{ ���VEL@���{ 0�$Ō!I]`���MT�ACFG>���  �@@ =O�"NORE-0l@,o�V�SI.1�d��6��"UXK�fP!��D�E�� $KE�Y_�3�$J3OG��0SV���0���!��}�SW�"�ah\aS�ՐT|�GI����| ^�� 4 �h��'d2�!XYZ�c���31�_ERR#�� 8Ԡ�A�fPV�d��1����/$BUF��X�����MOR|�� HB0CUd�lA�!��GQ�\aB�,"!a$� ���a��u��?��G~�� � $cSIՐ���VO��<T�0OBJE_���ADJU)B��EL�AY���%�DR�O�U.`=ղВQ0b=��T���0���;BDIR���; I�"�0DYNW�2��T���"R���@�0�"��OPWORK����,%@SYSBUy�SOP��ޑ�U�; P�pN�<��PA�t�>�"��OP�PUd!0�`!�Ľl�IMAGw��B0y�2IM�Õ�I�Ne�d��RGOVCRD��-��o�Pq����0��J�Os���"L�pBa���o�PMC�_Ee`���1Ny M� A�21�2T���S�L_��� � $OVSL�ǫ�?qD�`��2�" -�_�� k�P��k�Pu���2�C� �`�Ź�^��_ZER�D��$G�� 82=���� @*����%Oh`RI��� 
 JP8+��=!/��L��ح�T� �0A�TUS��TRC_T���sB��}f�s�9s�1Re`��� !DFAm����L���"`��0a� ޱ��XEw {�����C0�vUP��+p	qPX�P�j�43 � ��PG\���$SUBe�%�qe9JMPWAIT ,z}%LO��F�A�RCVFBQ�@x"�!qR�� �x"ACC� �R&�B�'IGNR�_PL9DBTB2�0Pqy!BWbP�$2w�Uy@�%IGT�P=I��TNLN�&2�R��rL�NP��P�EED \HADCOW�06�w��E[pq4jO!�`SPDV!� LbAz�`�07�3UNIr��02"!R��LYZ`� �o/PH_PK���e�RETRIE9{�q���0'P;FI"�� �G`�0�D 2�g�DB�GLV�#LOGS�IZ��EqKT�!Ud��VDD�#$0_T�
G�MՐCݱ��|@eM�RvC}�3�CHECAK0���0O�V!�kЙI��LE(!��P�ArpT�2K�W��0I�P2V!� h $ARIBiR� c�a�/�O�P8�ӐATT ��2�IF|@z�Aq4S��3UX����PL9I2V!� $g���OITCHx"[�W ��AS9�wSLL�BV!�� $�BA�DYs��BA�M!���Y9�PJ�5��Q��R6�V�Q_�KNOW�Cb��UF��AD�XV��0D�~+iPAYLOAt���Ic_��Rg�RgZ�OcL�q��PLCL=_�� !7��bP�QB��d���fF�iAC֠�js��d�I�h!Rؠ�g�ҢdB���љJ��q_J�a#���AND��Ĳ.t�bؤaL!q�PL0AL_ �P�0���QTրC��DNcE����J3CpWv� TPPDCK������>P�_ALPHgs�s�BE��gy|��K�1�� � �\��HoD_1Oj2ydDP�AR�*��;��&���TIA4U�5:U�6��MOM��a����n���{�Y�B� A�Da���n���{�PUB��R��҅n�҅{��/2�Wp��W � � PMsbT� �BxQ���� e$PI��81���TgJ��niJ�IV�Id�Ir��[��3!��>!��r�Ӫ�U3HIG�SU3�%�4� �4�%� ���"����!x
��!�%SAMP����^��_��%�P4s ю���[ 	ӝ� 3 ���0���&�C��� ��^��Sp��H&0	�IN�SpB�������"��6��6�V�GA�MM�SyI�� E�Tْ��;�D�tA�
�$ZpIBR!62I.T�$HIِ_���$C�˶E��ظAҾ���LWͽ�
���7Ơ��rЖ,0�qC�%C�HK��" �~I_A�����Rr� Rqܥ�Ǚ��ԥ���Ws� �$�x �1���I7RCHk_D�!� RN{��#�LE��ǒ!,���x���90MSWF�L�$�SCR((1#00��R@��3]B�րç��a����َ0��P�I3A9�METHaO����%��AXH��XX0԰62ER)I��^�3��R�0$u�	��pF{�_���$?ⲣ1�L�L�_�a�OOP����wᲡN��APP:���F��`�@{���أRT�V�OBp�0T����;��� 1�I��� ��lr���RA�@MGA1o���SSV-�w�P_@CURg��;�GRO[0S_�SA�Q��Y�#NO�pC!"�tY�� Zolox�������!b��,��&�DO�1A���A ����Х��A���A"�0WS�c L"h�*�� � ��YQLH�qܧ��SrZ�]B�o�=�q�Ô�q_�C1��M_W���g���c�M� �`Vq�$Ap�x1o�3"�PMJ�,�� �'A� 9�!YWi:�$�LWQ |ai�tg�tg�tg{t� �N`���S��JSpX�0O�sRqZ���P� *�� ���M��������������PX��� ��5L�q_~R� |�q#(Y����& n��&{�Y�Z��'�&t���Q��D�#0��@�}`�$PQ�PMO�N_QUc� �{ 8�@QCOU��n%PQTH��HO�n^0HYS:PES�RF^0UEI0O��0O|T�  �0PGõz�RUN_TO�r@Oْ.�� PE`�5C��A<�IND}E�ROGRA�nP� 2g�NE_NO�4�5IT��0�0�INFO�1� p�Q�:A��$PA�B� (��SLE�QݖFAѕF@�6� OySy�T� 4�@�ENAB��0PT�ION.S%0ERV�E���G���1{BGC]F�A� @R0J$�Rq�2���R�H�O�G "�EDITN�1� �v�K�jޓʱE�NU0W�*XAUTu�-UCO�PY�ِN\����M�ѱNXP\[q�PRU�T9� _RN�@OUC�$G�2�T����$$CL`?0[��&������Г �P�S�@�X��PXK�QIGRTU��_�PA� _WRK 2 e��@ 0 � �5�QMoYh\Jo|m |l	�`�m�o��`��o�o�f�e�l}�aI�[ct'`BS�*� �1�Y� <7����� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P��b�t���������srC�C��LMT?0����s  dѴIN�ڿ�дPRE_EXE��)�Ƅ0jP���za'`DV��S��@e)�%s�elect_macro����kϤ�qt�IOCNVVB�� 5��P��USňw����0V 14kP $$p��a�|�`?���߰>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ ���$�ѰLARMRE?COV ^������LMDG ��Ь�LM_�IF ��d���IF-157 �Menu can�not be d�isplayed�  (TCP) �) O���� ���)�;�M�_�q��, 
 ���#��>TELEOP ~ǘLINE 0Ǒ�AUTO ABO�RTEDǘJOI�NT 100 %�����$���1���A�����������ȯ��ANGTO�L  @� 	 A   ��Ѱ�PPINFO �� f�L�^�p����  ������ k���ۿſ�����5���Y�C�iϏ�%��� ٯ����������'߀9�K�]�o߁ߓߙ�P�PLICATIO�N ?t���|�Ha�ndlingTo�olǖ 
V9.40P/17�~��
8834ؒ���F0�	�549���������7DF�5�О�ǓNone���FRA�� �69��_ACoTIVE1�  ��� �  ��ސMO�D��������CH�GAPONL�� ��OUPL[�1	��� >�B�T��f���CUREQ �1
��  Tp�
p�p�	�������� l�������������xi3l�p�g���^H���A�t
HTTHKY�FXv|�� *<N`�� ������// &/8/J/\/�/�/�/�/ �/�/�/�/�/?"?4? F?X?�?|?�?�?�?�? �?�?�?OO0OBOTO �OxO�O�O�O�O�O�O �O__,_>_P_�_t_ �_�_�_�_�_�_�_o o(o:oLo�opo�o�o �o�o�o�o�o $ 6H�l~��� ����� �2�D� ��h�z�������ԏ ���
��.�@���d��v�����������TO������DO_CL�EAN���E�NMw  �� p��������ɯۯv�DS�PDRYRL���H	I��o�@��G�Y�k� }�������ſ׿���8�ϻ�MAX��,�呿��=�X,�<�9�|<���PLUGG,�-�9���PRC��B�m�q�6�(ϗ�Ox����SEGF�K���� �m��G�Y��k�}ߏ�����LAP $�7ޡ������+� =�O�a�s�����> �TOTAL_ƈɾ �USENU$��1� ������RGDISPMMC�ed�C�O�@@��1�O"�D��-�_�STRING 1���
�M���S��
��_I�TEM1��  n ��������� $ 6HZl~��������I�/O SIGNA�L��Tryout Mode���InpNSim�ulated���Out`OV�ERR!� = 1�00��In c�yclT��Prog Aborj���JStatu�s��	Heart�beat��MH� Faul��Aler�!/!/3/�E/W/i/{/�/�/�/ (���(����/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O84OFO�/WORИ� ~A�/XO�O�O�O�O�O  __$_6_H_Z_l_~_��_�_�_�_�_�_�^PO���"`�KoEo Woio{o�o�o�o�o�o �o�o/ASepw��bDEV%n �p9o����#�5� G�Y�k�}�������ŏ�׏�����1�C�PALT�-j��OD� ������ȟڟ���� "�4�F�X�j�|�����p��į֯X�GRIB� ������6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�z�����R�-��&������� ���"�4�F�X�j�|� �ߠ߲����������<��PREGn�W� ��0�~�������� ����� �2�D�V�h��z���������$�$�ARG_~@D ?�	�����  	�$$	[]��$:	��SBN_CONFIG��XWqRC�II_SAVE � $zm��TC�ELLSETUP� 
%  O�ME_IO$$%?MOV_H� ���REP��#��U�TOBACK� �	tFRA;:\D� .D�z '`�D�w� �s  �25/11/2�9 20:26:16D�;D���#//h��C/j/|/ �/�/�/�/D�X/�/ ??(?:?L?�/p?�? �?�?�?�?�?g? OO $O6OHOZO�?~O�O�O�O�O�O�O���  �c_F_\ATB�CKCTL.TM��)_;_M___q_8INIm��j~C?MESSAG� �Q�z �[ODE_D(� �j�XO�p�_�@PAUS6` !�� ,,		�; :oHg.oho Rotovo�o�o�o�o�o��o@*<v���d`TSK  �mw}_CUPD�T�P�Wd�p�VXWZD_ENB�Tf
�vSTA�U�u���XISX UNT� 2�vwy � �	 ������g1���i0gK5h�D�R�����D�z������F�� �jc �D�� ', Q� �Ir��������,�/�MET��2�@��y PQ�?��fU??�?W��P>�f�?U�~?�N�>�caA=��=��<��d<z��>i5��SCRDCFG �1Y ��� ���@�%�7�I�pD�Q�	 ܟ������ϯ��Z� �~�;�M�_�q�����0��6���FGR9��pX�_ԳPNA� s	FѶ_ED�P�1��� 
 ��%-PEDT-`¿ R�v���Es�� -FE�D�;�9/�>���  ����2�����B� ��ˀ�{�����j�����3 ��#� �G�Y���G����6�����4����� �Yި��Z�l������5K������Y�t�@��&�8���\���6 ��d��Y�@����(��7�S0w Y�w��f���!8�W��{�IZ��@C/��2/���9{/��//LZݤ/?V/0h/�/�/��CR�� �?�?Tn?�? ?2?�?�V?԰!�NO_DE�L�ҲGE_UN�USE޿дIGALLOW 1��   (*SYSTEM*
��	$SERV_�GR[�@`REGƜE$�C
��@NU�M�J�C�MPMU|?@
�LAYK��
�PMPA�L�PUCYC10� N3^P!^YSUL�SU_�M5Ra�C�Lo_�TBOXOR=I�ECUR_�P�M�PMCNVV��P10I^�PT4�DLI�p�_�I	*�PROGRA�D?PG_MI!^KoF]`AL+ejoTe]`�B�o�N$FLU?I_RESU9W�o�O�o�dMR�N�@�<�?�;M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3��E�W�2BLAL_OUT �K���WD_ABOR:P�cO��ITR_RT/N  �$�빸�?NONSTO��� lHCCFS_UTIL ��̷CC_AUXA�XIS 3$� h}�j�|�����ƽ�CE_RIA_IL`@�נ��FCFG $��/�#��_LIMv�B2+� �� 7� 	��B\���$�� 
Ԡ��)�Z��%�/�����[����� ���!�����L��(
5������PA�`GP 1H�����A�SϨe�w�6�CC� CU7��J��]��p��}����� C���U������������Ué�̩�ձ�ߩ�U�������;����PCk���������������������Ա��������� D� D!��!�!�!� ���&?��HE@O�NFIpC�G_�P�P1H�  +EH��ߟ߱�����������C�KPAUSf�Q1H�ף b �S�H�A��e��� ������������E��+�i�{�a���A�?Iץ�MؐNFO� 1���� �3��$4�@k��?��@i�*:�]/H�ȿr��
=q�*� D�C�����D
�1���@�G����Y�Pb�O�� � ��LLECT_�!������EN+`�ʒ���N[DE�#�/��1234567890�"�A��H/ҵHw��#)j ��<i{��;�� /��/`/+/=/O/ �/s/�/�/�/�/�/�/ 8???'?�?K?]?o? �?�?�?�?O�?���$� ��I�O &��"S�▒O�O�O�O`GTR�2'DM(��^�?�NN�(oM Z��o_MOR)q3)H��7ىU3��Y�_�_�_@�_�_�[bR�kQ*H�%,S�?<�<Ѡ<cz�QKFd���P,��;ϒo�o�o˿�oP�oœh�UY@E��oS �s�ja�PDB.����4cpmid�bg3��Рs:���>uqpz��v  ��>x��}�.��}�`��|�<�mgP���t��~f�������@ud�1:�?��XqDE�F -��zC)�*�cO�buf.t�xtJ��|K�[`�/zDM��>���Rl�A��MCiR20_{bRCd���hS21�1���G���CzA�d�4�A"R�A��A=.�?���A<� A%�B��\B���GBԖ�A����B�OB����D]^Dc���D���C@��jD��Db��ӭ��Ufg23FDLD�	>z�!� Y2��}��yc
�@�x9� C�Ĵ�  D4G�E����  E%q��F�� E�p��u�F�P E���fF3H ?��GM��Ъ>5�>�33��?��xn9�q@�Q5�����RpA?a��=�L��<#�QU��@,�Cϒ���RS�MOFST +xi�����P_T1Ɠ�4DMA =ք�M?ODE 5dm�@c��	Q�M;���%��?���<�M>��Ͷ�/TESTc�2i�`�ER�6�O�K�CN�QAB���n� 8��\�n�CdB���C�pp�����p:;d�QS ��ՠ ������4�I7R>���>B8m5�$�RT_c�PRO/G %j%��d�|1�h@NUSER���x�KEY_TBL�  e�����	�
�� !�"#$%&'()�*+,-./(:�;<=>?@AB�Cc�GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������>���͓���������������������������������耇��������������������4A8�LCK��F�y��OSTAT��2�X��_ALM�����_AUTO_DO��E�FDR 3]:i�2hi�US�x��i�$g� �A������ T*g�2� bf ��/�/9/;�*p m�P/z/�~/h/�/�/ �/�/�/?"=�G?Y? k?/|?�?L/�?�?�/ �?�?OO�?*O@OvO �O6?�O�O�O~?�O	_ �?*_$_BOD_6_p_~_ T_�_�_�_�_�Oo)o ;o�OLoqo_�o�o�_ �o�o�o�o�o�oF Xo��No�� �o����@�N� $�b�x�����n��� ���A��b�\�z� |�n�������ʟ��� (�֏O�a�s������ T�ʯį��֯�� ��2�H�~���>���ɿ ۿ���ϼ�2�,�J� L�>�xφ�\Ϛϰ��� �Ϧ��1�C��T�y� $Ϛߔ߲ϴߦ����� ����N�`�߇�� ��V߼�������� ��H�V�,�j����� ��v�����$I ��jd���v�� ���0��Wi {&��\��� ��/&/�:/P/�/ �/F�/�/�/��/? �:?4?R/T?F?�?�? d?�?�?�? O�/'O9O KO�/\O�O,?�O�O�? �O�O�O�O�O
_ _V_ h_O�_�_�_^O�_�_ �O
oo"_$ooPo^o 4oro�o�o�o~_�o	 �_,Q�_rl�o �~�����&� 8��o_�q���.���� dڏԏ��� �.� �B�X�����N�ǟٟ 럖���!�̏B�<�Z� \�N�����l������� ���/�A�S���d��� 4�����¯Ŀ����� Կ�(�^�p���ϩ� ��f����Ϝ���*� ,��X�f�<�zߐ��� �߆����#���4�Y� �z�t�ߔ������ ������.�@���g�y� ��6����l������� ����(6J`� �V������) ��JDbdV�� t���/�7/I/ [/l/�/<�/�/� �/�/�/?�/?0?f? x?&/�?�?�?n/�?�? �/OO2?4O&O`OnO DO�O�O�O�O�?__ +_�?<_a_O�_|_�O �_�_�_�_�_�_ o6o Ho�Ooo�o�o>_�o�o t_�o�oo�o0> Rh��^o�� ��o�1��oR�L�j l�^�����|���Џ� ��?�Q�c��t��� D�����ҏԟƟ �� �"�8�n���.����� ˯v�ܯ���"��:� <�.�h�v�L�����ֿ 迖��!�3�ޯD�i� ��τϢ��ϖ����� �����>�P���w߉� ��FϬ���|�����
� ���8�F��Z�p�� ��f���������9� ��Z�T�r�t�f����� ������ ��GY k�|�L����� ���*@v �6���~�	/ �*/$/BD/6/p/~/ T/�/�/�/�/�?)? ;?�L?q?/�?�?�/ �?�?�?�?�?�?OFO XO?O�O�ON?�O�O �?�O�OO__@_N_ $_b_x_�_�_nO�_�_ o�OoAo�Obo\oz_ |ono�o�o�o�o�o (�_Oaso�� To���o���� �2�H�~���>��ɏ ۏ����2�,�J� L�>�x���\������ �����1�C��T�y� $������������� į��N�`������ ��V���ῌ����� ��H�V�,�jπ϶� ��v����߾�$�I� ��j�d߂τ�v߰߾� �������0���W�i� {�&ߌ��\������� �����&���:�P��� ��F���������� ��:4R�TF�� d��� ��'9 K��\�,��� �����
/ /V/ h/�/�/�/^�/�/ �
??"/$??P?^? 4?r?�?�?�?~/�?	O O�/,OQO�/rOlO�? �O~O�O�O�O�O�O&_ 8_�?__q_�_.O�_�_ dO�_�_�O�_�_ o.o�oBoXo�otc�$C�R_FDR_CF�G ;re��Q
UD1�:�W�TJ�d  ��`�\�bHIST �3<rf  �` � ?�RU@tAtBtC�PUpDtEtIt)gqpotw�_���bINDT_EN�6p�T��q�bT1_DO�  �U�u�sT2���wVAR 2=ֹg`qh_r ���R��d4��d�m[��RZ��`STOP��rT�RL_DELET�Np�t ��_SCREEN re~�rkcsc�r�Uw�MMENU �1>��  <�\%�_��T�� R��S/�U���e�w�ğ ������џ�	�B�� +�x�O�a��������� ��ͯ߯,���b�9� K�q�������࿷�ɿ ����%�^�5�Gϔ� k�}��ϡϳ������ ��H��1�~�U�gߍ� �ߝ߯�������2�	� �A�z�Q�c���� �������.���d� ;�M���q�������������YӃ_MAN�UAL{��rZCDƳa?�y�rG +���R�f"
�"
?|(��PK�W�GRP 2@�y�aqB� � s���� �$DBCO��pRIG���v�G�_ERRLOG A��Q�I[�m �NUMLKIM�s��u
��PXWORK 1B�8���/|/�}DBTB_��� C%�ap��S"� �aDB_AW�AY��QGCP� �r=�ןm"_�AL�F�_�Y�z����p�vk  1}D� , 
�`�/"�/%?/(_M�p�qw,@�=5ONT�IM����t��_6�)
�0�'MO�TNENFpF�;R�ECORD 2J�� �-?�SG�O��1�?"x"!O3O EOWO�8_O�O�?�OO �O�O�O�O�O(_�OL_ �Op_�_�_�_A_�_9_ �_]_o$o6oHo�_lo �_�o�_�o�o�o�oYo }o2�oVhz� �o��C�
�� .��R��K������ ��Џ?��ߏ�*��� ��+�b�t�㏘����� Ο=�O�����:�%� ��p�ߟ񟦯��O�ǯ �]������H�Z�� �������#�5�����ϩ�i"TOLER7ENCv$Bȿ"� �L��� CSS_�CCSCB 2K�\0"?"{� �ϟ���7��
���π@�R�d�3߈ߚ�"� x���������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ��1CUgy��� �������R�LL]�L�a�m1T#2 C�C��Fή^ A�C�pC���#�0� 	 gA���B���?�  �$����\0袰�0��B��`#s�K/]/o/�ϓ/�/�/s/��/�/��ʈ����5οRr���o;�&;�'���/��/`?*;�@��O?�?�?�?Ȏ0AF��?{F�A OO�7�1���9M	AB
AZOdB�AE�9$O�O�O�Oi:Pz��`�@0�DJ�CA� @��
�X-.
[#_  	 M?�>O�ڴ�q_@�_�_�_:W�A<o :[<ǲ/o�/�_�+oPoboto�eAC�HC�V�WB$�Dz�cD�`�a=/�o�o o�oW�a.+!���2=t,yD��YqC��I?�-t �s�js�w�yj��������Q��� �@`��$�����A�� ��Bމ�o��'�9� �_]�o�N���r���ɟ ۟_�B�ʄ��YZ�>`��@'BO��Be�@�V�z�RW�:C��l�R�d�v�����  `_м¯���
��� ̯9�,�]�o��� �H� ����ٿ뿊��ƿ3� E�W�iϬ���$ϱ��� �� Ϟ����/�A�S� ��w�V�h߭ߌ��S���ߐ�_�f	�� H�?�Q�~�u���� ���������D�� -�g�q����������� ��
@7Ic�m��߾�   �����)M@ qdv����� ��//I/P�m/� v/�/�/�/�/�/�/�/ ?3?*?<?i?`?r?�? ^/�?�?�?�?�?O/O &O8OJO\O�O�O�O�O�O�O�O�g	 � Q�P�s� �PC4p*�p�p6U6P\Cu9p/p�� ]VT^PM]�6P�:P�>P��VJ_�^P�bP�0fP�Vr]v��Tp Q�
k���_oo�id1Q&oNo ;o_cox�oˏUUA   �o<�k1Q@�  �o�kt�b����逡Up �� 1��6�1C���C�cPfL��?#�c>�{����`�cP�@@��d��r�`B�cP>�s�qC��p�����b�t<�o?��PH�)S�B���tq�q�p�r�`B���eIC�&�Q�4(� �oz�UU�5��=��Bd�=�^��RT�:C�H�Q�-R�?�����C���B��F��b��`ځ`  ?�p���U�[?���}t��$����$DCSS_CLLB2 2M��p�P�^?��NSTCY 2N����  �������ʟ؟ ���� �2�D�Z�h� z�������¯ԯ��S�A�DEVICE K2O��!�$�� 4&V�h�������˿¿ Կ���
�7�.�[�R� ϑϣϵ�����4(A��HNDGD P̅�*�Cz�A�LS 2Q��_�Q�c߀u߇ߙ߽߫���?�PARAM RP���1�`�&�RBT �2T�� 8r�P<C�'p �qdi�l��s@"�R��4(qI�X��0�pB oCW  ��B\x�`N��`Z����%��)���X�j��p����$zq�����B �(s,�F�p�V��q���Xb��B ��4&c � S�e�l�4+����Hx1~����D��C�$Z��b����A,� 4�u@��X@��^@�w���]B����B�cP%��C4��C3:^C4���nЬ ��p8��-B{B?��A���� �l��C�C�3�JC4jC�3��yn+�3 �Dff 2�A PB W4+@:�]o �W�����/ �/P/'/9/K/]/o/ �/�/�/�/?�/�/�/ ?#?5?�?Y?k?�?�? �o�?�?O�?6O!OZO lOWO�O�Es�?�?�? �O�O_�O�OL_#_5_ G_Y_k_}_�_�_�_ o �_�_�_oo1o~oUo go�o�o�o�o�owO  D/Aze�� ��O�o�o
��o�� R�)�;���_�q����� �����ݏ�<��%� r�I�[�m�������� ǟٟ&�8��\�G��� k�������گů��� ��F��/�A�S�e� w�Ŀ������ѿ��� ��+�x�O�aϮυ� �ϩϻ�����,��� b�t�ﯘ߃߼ߧ��� ������:��C�U� ��Y�k������� ����6���l�C�U� g�y�����������  ��	-?Q�� �����@ +dvQ���� ����*///%/ r/I/[/�//�/�/�/ �/�/&?�/?\?3?E? �?i?{?�?�?U�?�? "O4OOXOCO|OgO�O {��?�O�?�O�O0_ __f_=_O_a_s_�_ �_�_�_�_o�_oo 'o9oKo�ooo�o�o�o �o�o�O:%^I�������H��$DCSS_SL�AVE U����	��~�z_4D  	���AR_MENU V	� �j�|� ������ď�BY��� ��~?�SHOW �2W	� �  �b�aG�Q�X�v����������П֏����  @�:�d�a�s������� ���߯��*�$�N� K�]�o�������̯ɿ ۿ���8�5�G�Y� k�}Ϗ϶��������� ��"��1�C�U�g�y� �ϝ߯��������	� �-�?�Q�c��s�� ������������)� ;�M�t���������� ������%7I p�m�������� ��!3ZWi ���J���� //DA/S/e/��/ ��/�/�/�/�/?./ +?=?O?v/p?�/�?�? �?�?�?�??O'O9O `?ZO�?�O�O�O�O�O �OO�O_#_JOD_nO k_}_�_�_�_�_�O�_ �_o4_.oX_Uogoyo �o�o�o�_�o�o�oo Bo?Qcu����o:���CFG7 X)�3�3q�5p�FRA�:\!�L+�%04_d.CSV|	pm}� �qA g�CHo�zv�	����3q�����́܏�� ���4��JPQ����qp1�� �RC_OUT [Y��C���_C_FSI �?i� .�������͟��� ��>�9�K�]����� ����ίɯۯ��� #�5�^�Y�k�}����� ��ſ�����6�1� C�U�~�yϋϝ����� �����	��-�V�Q� c�uߞߙ߽߫����� ���.�)�;�M�v�q� ����������� �%�N�I�[�m����� ������������&! 3Eni{��� ����FA Se������ ��//+/=/f/a/ s/�/�/�/�/�/�/�/ ??>?9?K?]?�?�? �?�?�?�?�?�?OO #O5O^OYOkO}O�O�O �O�O�O�O�O_6_1_ C_U_~_y_�_�_�_�_ �_�_o	oo-oVoQo couo�o�o�o�o�o�o �o.);Mvq �������� �%�N�I�[�m����� ����ޏُ���&�!� 3�E�n�i�{������� ß՟������F�A� S�e���������֯ѯ �����+�=�f�a� s���������Ϳ��� ��>�9�K�]φρ� �ϥ����������� #�5�^�Y�k�}ߦߡ� �����������6�1� C�U�~�y������� �����	��-�V�Q� c�u������������� ��.);Mvq ������ %NI[m�� ������&/!/ 3/E/n/i/{/�/�/�/��/�/�/�/3�$D�CS_C_FSO ?���71� P ??T?}?x?�?�? �?�?�?�?OOO,O UOPObOtO�O�O�O�O �O�O�O_-_(_:_L_ u_p_�_�_�_�_�_�_ o oo$oMoHoZolo �o�o�o�o�o�o�o�o % 2Dmhz� ������
�� E�@�R�d��������� ՏЏ����*�<� e�`�r���������̟ �����=�8�J�\��������?C_RPI4>F?����� ��3?�&�o����� >SLү@d����� �%�7�`�[�m�Ϩ� �ϵ����������8� 3�E�W߀�{ߍߟ��� ���������/�X� S�e�w������� �����0�+�=�O�x� s������������� 'PK]o� �������( #5Gpk}�� ���Q���/6/1/ C/U/~/y/�/�/�/�/ �/�/?	??-?V?Q? c?u?�?�?�?�?�?�? �?O.O)O;OMOvOqO �O�O�O�O�O�O__ _%_N_I_[_m_�_�_ �_�_�_�_�_�_&o!o 3oEonoio{o�o�o�o �o�o�o�oFA Se�������>�NOCODE �ZU���?�PRE_CHKg \U��pA �p��< ���pU�]�o�U� 	 <Q��������ۏ� Ǐ�#����Y�k�E� ����{�şן��ß� ���C�U�/�y����� s���ӯm���	��� ?��+�u���a����� ��ɿ�Ϳ߿)�;�� _�q�K�}ϧϝ����� �ω���%����[�m� Gߑߣ�}߯��߳��� �!���E�W�1�c�� g�y����������� ��A�S�-�w���c��� ����������+= asM_��� ���'�] o	����� �/#/�G/Y/3/e/ �/i/{/�/�/�/�/? �/?C?9Ky?�?%? �?�?�?�?�?	O�?-O ?OOKOuOOOaO�O�O �O�O�O�O�O)___ __q_K_�_�_a?�_�_ �_�_o%o�_Io[o5o Go�o�o}o�o�o�o�o �o�oEW1{� g���_���� /�A��M�w�Q�c��� �������Ϗ�+�� �a�s�M��������� ߟ���'���3�]� 7�I������ɯۯ�� �����G�Y�3�}� ��i���ſ������� �1�C���+�yϋ�e� ���ϛ���������-� ?��c�u�Oߙ߫߅� ���������)��M� _�U�G���A����� ���������I�[�5� ���k����������� ��3EQ{q� ���]���� /AewQ�� �����/+// 7/a/;/M/�/�/�/�/ �/��/?'??K?]? 7?�?�?m??�?�?�? �?O�?5OGO!O3O}O �OiO�O�O�O�O�O�/ �O1_C_�Og_y_S_�_ �_�_�_�_�_�_o-o o9oco=oOo�o�o�o �o�o�o�o__M _�ok�o��� �����I�#�5� ���k���Ǐ��ӏ�� ׏�3�E��i�{�5 c���ß�����ӟ� /�	��e�w�Q����� ��ѯ㯽�ϯ�+�� O�a�;��������Ϳ ߿y����!�K�%� 7ρϓ�mϷ��ϣ��� ������5�G�!�k�}� W߉߳ߩ������ߕ� �1���g�y�S�� ����������-� �Q�c�=�o���s��� ����������M _9��o��� ��7I#m Yk����� �!/3/)/i/{// �/�/�/�/�/�/�/? /?	?S?e???q?�?u? �?�?�?�?OO�?%O OOE/W/�O�O1O�O�O �O�O__�O9_K_%_ W_�_[_m_�_�_�_�_ �_�_o5oo!oko}o Wo�o�omO�o�o�o�o 1UgAS� �����	��� �Q�c�=�����s��� Ϗ�o������;�M� '�Y���]�o���˟�� ��۟�7��#�m� �Y����������� �!�3�ͯ?�i�C�U� ������տ����� ��	�S�e�?ωϛ�u�����ϫϽ�������$DCS_SG�N ]	�E���-���29�-NOV-25 ?20:38 ��N��27_�x�x� _[}�t��q�����xҚك�JѨ�E�ƼÞ� ���ǖ�  1�HOW� ^	�� x�/�VERSION =��V4.5.2���EFLOGIC� 1_���  	�����C��R��%�PROG_EN/B  ��:�{��s�ULSE  �X��%�_ACC�LIM������d��WRSTJ�NT��E��-�E�MO|�zя�$���I?NIT `2�����OPT_SL� ?		�	�
 ?	R575��]�74b�6c�7c�50��1���C���>@�TO  L���t �V�DEX���dE�x�PAT�H A=�A\�k}��HCP_�CLNTID ?<�:� D������IAG_GRoP 2e	�����z�	 @��  
ff?�aG���B�#  2��/�8[�I@c�ς!��7@�z�@^��@
�!���mp2m15 8�90123456�7����  �?��?�=�q?��
?޸�R?�Q�?��ׅ?�����(�?�z���x��@�  A_�ApX !7A�88v_�B4�� ���L�x�
�@��@��\@~�R�@xQ�@q��@j�H@c�
�@\��@U�@Mp��//'$��; �O)H��@�Ct >d 9��@}4�/\)@)� �#t {@���/�/�/�/�/P'?_���?����_ ?}p�?u¿�?n{?s ?\�Q�? ?2?�D?V?h8�
=?�����0w5�z��H?p�h��?^�R�?�?�?�?�?Th8��t0��Y�@�?��0� ;@&O8OJO\OnOP'� $_�_Y_k_�O?_�_ �_�_�_�_s_�_�_1o Co!ogoyoo�o��B�j"� �2{1�@"?����f�t0�d"5�!�
u4V���u"�B3t�A>u��?�@[q��@`,=�q�=b��=��E1>�J�>�n�>��H"�<�o �z�sT�q��� �x�C�@�<(�Uz� 4��� ����A@x�?*�o��m*�P� b���tn���2���Ώ����i>J���&�bN2�"��G�N��o@�@v���0����@ffrr!l ��33�(��"C��� ƒI�CH��)C.dBتA"8"����'�� �"~�A?�&"K����pf�B��@�p��������p��?}Wͽ��r�������@�~Ᵹ�-M��Cu=�TG��}�)D��C�Ҭ�D�xО�������3��N�T������1��@�G����Y�@Rs"����ǿ���ֿ�����<O3[>���P�_�Ǿ��J���#��!�o��CT_CONFIG f���|�eg�Y��STBF_TTS��
����О�t}���1�MAU�������MSW_CF���g�  # ��O�CVIEW��h!�-���s߅ߗ� �߻��ߟ�a����� ,�>�P���t���� ����]�����(�:� L�^������������ ��k� $6HZ ��~������ y 2DVh��������v�R%C�i���!�0. /S/B/w/f/�/�/�/���SBL_FAULT j*6��!GPMSK���'���TDIAG k���-�������UD1: 67�89012345 I2��=1���%P\υ? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�Od696�I�r
t?�O|ƟTRECP"?4:
 B44_[7M[s?p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�O�O��O�o7�UMP_O/PTIO=��.�a�TR����)uP�ME��Y_TE�MP  È�+3BC�gp�B�Qt�UNI����gq�Y�N_BRK l�L�7�EDITOR��a�a@�r_
PEN�T 1m) � ,&TPSN�AP^P ��l&M�TPG�p��T�ELEO+�f�&�/�����z����� ۏ����5��Y� k�R���v���ş��� П����C�*�g�N� v������������ޯ���?�Q���EMGDI_STAzu�V�gq�uNC_IN�FO 1n!��b���X���������vn�1o!� ��o(����
�d�oU� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߽߫��� u���� 
��*�B�*�P�b�t� ������������ �(�:�L�^�p����� ����2������� 9�CUgy��� ����	-? Qcu������ ��//1;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?m?? �?�?�?��?�?�?O )/OEOWOiO{O�O�O �O�O�O�O�O__/_ A_S_e_w_�_�_�_�? �?�_�_o�_3O=oOo aoso�o�o�o�o�o�o �o'9K]o ����_�_��� �+o5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� �ӟ���	�#�-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ���7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� �����������%�/� A�S�e�w����� ��������+�=�O� a�s������������� ���'9K]o �������� #5GYk}� 	������/ 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?��?�? �?�?/O)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�?�_�_�_�_O�_ !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew��_�_� ���o�+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ������ɟ۟�� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߝ��߹������� ���%�7�I�[�m�� ������������� !�3�E�W�i�{��߇� ���������/ ASew���� ���+=O as�������� ��//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?�� �?�?�?�?��?OO 1OCOUOgOyO�O�O�O �O�O�O�O	__-_?_ Q_c_u_�?�_�_�_�_ �?�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m�_ u����_��� !�3�E�W�i�{����� ��ÏՏ�����/� A�S�e�������� u������+�=�O� a�s���������ͯ߯ ���'�9�K�]�w� ��������ɿ���� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g߁��ߝ߯� ��ۿ����	��-�?� Q�c�u������� ������)�;�M�_� y߃������������� %7I[m ������� !3EWq�c�� �������//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? i{�?�?�?�?��? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_�?s?}_�_ �_�_�?�_�_�_oo 1oCoUogoyo�o�o�o �o�o�o�o	-? Qk_u����_� ����)�;�M�_� q���������ˏݏ� ��%�7�I�cQ�� �������ٟ���� !�3�E�W�i�{����� ��ïկ�����/��A�[� �$ENE�TMODE 1p���� + k�k�f������j�OATCFG� q�����Ѵ��C���D�ATA 1rw��Ӱ���*	�*@��'�9�K�]�l�dl���e��ϻ����� ����'ߡϳ�]�o� �ߓߥ߷�1���U��� �#�5�G�Y����ߏ� �����������u�� 1�C�U�g�y������ )�������	-�� ��cu������j�RPOST_L%O��t�[
׶�#5Gi�RROR�_PR� %w�%�L�XTABLE  w�ȟ�����RSEV_N�UM ��  ����  �_A�UTO_ENB � ���X_NON5! uw���"_  *�x �x %�x �x + +w �/x�/�/Q$FLTR=/O&HIS#]�J+_ALM 1vw�� �[x,e�+�/Q?c?u?�?�?�?r�/_"W   w��v!���:j�TCP_VER !w�y!x�?$EXT� o_REQ�&�H)�BCSIZKO=DST�KhIf%�?BT�OL  ]Dz��"�A =D_BWD�0�@�&�A���C;DI�A wķ�x��]�KSTEP�O��Oj�POP_DO��Oh�FDR_GR�P 1xw��!d �	�?�_��yPs��Y�Q'�M"����l��?T� ����VyS��_�]�TB CA���Az�m]�A^��_`���@՚��_�[Go 2oWo}oho�o�o�o�]�@\�G?�"��?k�)>��~�n
 F@c�`�bX.��o(2�o`�oZE~i|A@`��t@S33�uh}@ �q�g��yPq���|yPG�  @�Fg�fC�8RL���}?�  h��6��X����875�t��5���5�`+��~X����>� �y���_�|:� ��͓FEAT?URE y���@���Han�dlingToo�l �]En�glish Di�ctionary��4D St��a�rd��Anal?og I/O>�G��gle Shif�tZ�uto So�ftware U�pdate�ma�tic Back�up���ground Edit �~�CameraU��FY�CnrRnd�Im���ommo�n calib �UI��nˑ�M�onitor$�t�r�Reliab<n��DHCP �[��ata Acqu�is3�\�iagn�os��R�v�isp�layΑLice�nsZ�`�ocum�ent View�e?�^�ual C�heck Saf�ety��hanGced���s��Frܐ�xt. oDIO /�fi���@�end�Err�>�L��\�4�s[�r�P�K� �@
�FCT�N Menu��v|Z���TP In���facĵ�Gig�E־�Đp Ma�sk Exc�g�=�HT԰Prox�y Sv��ig�h-Spe�Sk�i�� Ť�O�mmuwnic��onsVȃur����q�V�ײc�onnect 2��ncrְstr�u!��ʴ�eۡ��J���X�KAREL �Cmd. L�u�a���Run-T�i<�Env�Ȟ�e�l +��s��S/�W�ƥ���r�Bo�ok(Syste�m)
�MACRO�s,M�/Offs	eu�p�HO���o�u��MR8�4���Mec_hStop+�t��D��p�im�q���x��R�����odo�wiGtch�ӟ�.��4�OptmF��,�'fil䬳�g��p�?ulti-T�Γ��PCM fun��Ǽ�o��������R�egie�rq���r�iݠF���S�Num Sel��/�:� Adjua�*�W�<q�h�tatu���ߪ�RDM Ro�bot�scov�e'���ea��<�F�req AnlyNq�Rem��O�n5�|����ServoO��!��SNPX b�-�v�SN԰Clixܡ?r�Libr&�D_�� ��q +oJ�=t��ssag��X��@ ����	�@/I|ս�MILIB�~�P Firm��:�P��AccŐ͛�TPTXk��el�n��������o�rquo�imul�a=��|u(�Pa�&��ĐX�B�&+�e3v.���ri��T�USB por[t �iPf�aݠ~&R EVNT�� nexcept������%5��VC"�rl�c���V���"��%q�+SR SC�N�/SGE�/�%U�I	�Web Pl ��>��A43��ۡ���ZDT App�lj�
�{1EOAT�����&0?�7Gr�id�񾡬=�?iR�".5� F���/ג�RX-10iA/�L�?Alarm �Cause/��e�d(�All Sm�ooth5���C�s�cii+�V�Loa9d䠌JUpl�@w��toS ��rityAvoidM(��s7�t�@�yc�n�����_�CS�+���. c��XJo���-T3_H�.RX���U���Xcollgabo����RA�0:�.9D��in����NRTHI
�On>��e Hel����`ֿ�����1trU�ROS Eth$р�A������;,�G 0�B�,|HUpV�%̸W�t ԰�_iR�S�ݐ�64MB �DRAM�o�cFR�O���L8F Fl�D�����2M �A:�o�pm�ԕex@V�
�sh�q��wce�u��Yp��|tyn�sA�
�%�r����J��^�1.v� P)Q/sbS��`���O�N��mai@��U���R�q�T1�^FC+Ԍ%̋�Fs9�ˌk̋��T[yp߽FC%�hױtV�N Sp�ForްK��Ԭ�lu!����c�p�PG j�֡�RtJ�[L`Sup"`}��֐f��crFPf��lu� ��al�����r��i�
q�4x@а�uest,?IMPLE ׀6�*|HZ���c0�BT�ea(�|���$rtqu���V�9HMI��ܤ��UIFc�po	no2D�BC�:�L� y�p���������ʿܿ 	� ��?�6�H�u�l� ~ϫϢϴ�������� �;�2�D�q�h�zߧ� �߰��������
�7� .�@�m�d�v���� ���������3�*�<� i�`�r����������� ����/&8e\ n������� �+"4aXj� �������'/ /0/]/T/f/�/�/�/ �/�/�/�/�/#??,? Y?P?b?�?�?�?�?�? �?�?�?OO(OUOLO ^O�O�O�O�O�O�O�O �O__$_Q_H_Z_�_ ~_�_�_�_�_�_�_o o oMoDoVo�ozo�o �o�o�o�o�o
 I@Rv��� ������E�<� N�{�r�������Տ̏ ޏ���A�8�J�w� n�������џȟڟ� ���=�4�F�s�j�|� ����ͯį֯���� 9�0�B�o�f�x����� ɿ��ҿ�����5�,� >�k�b�tφϘ��ϼ� �������1�(�:�g� ^�p߂ߔ��߸����� �� �-�$�6�c�Z�l� ~������������ )� �2�_�V�h�z��� ������������% .[Rdv��� ����!*W N`r����� ��//&/S/J/\/ n/�/�/�/�/�/�/�/ ??"?O?F?X?j?|? �?�?�?�?�?�?OO OKOBOTOfOxO�O�O �O�O�O�O___G_ >_P_b_t_�_�_�_�_ �_�_oooCo:oLo ^opo�o�o�o�o�o�o 	 ?6HZl �������� �;�2�D�V�h����� ��ˏԏ���
�7� .�@�R�d�������ǟ ��П�����3�*�<� N�`�������ï��̯ ����/�&�8�J�\� ����������ȿ��� ��+�"�4�F�Xυ�|� �ϻϲ���������'� �0�B�T߁�xߊ߷� ����������#��,� >�P�}�t����� ��������(�:�L� y�p������������� ��$6Hul�~����� � H552���21R78�50J614�ATUP'54�5'6VCAM�CRIbUIFv'28cNRE�52VR63S�CHLIC�DwOCV�CSU�869'02EI�OC�4R69�VESET?UJ�7UR68MA{SKPRXY{]7OCO#(3?h+ &3j&J6%�53�H�(LCH^R&OPLG?0�&�MHCRS&S�'MkCS>0.'552�MDSW+7u'OP�u'MPRv&��(0n&PCMzR0q7�+ 2� �'51J5u1�80JPRS"'�69j&FRDbFwREQMCN{93&SNBA�^�'SHLBFM1Gt�82&HTC>�TMIL�TP�A�TPTXcFELF� �8wJ95�TUTv'�95j&UEV"&U�ECR&UFRbV�CC
XO�&VIP�nFCSC�FCSGt��IWEB>7HTT>R6��Hl;RVCGiWIGQWoIPGS�VRCnF�DGu'H7�7R6�6J5'R�8R�51
(6�(2�(5�V�J8�86�L�=I% �84g66�2R64NVDv"&R6�'R84�gk79�(4�S5i'�J76j&D0�gFn xRTSFCR�gwCRXv&CLIZ8�ICMS�Sp>S�TYnG6)7CTOh>��7�NNj&�ORS�&C &FC�B�FCF�7CH�>FCR"&FCI��VFC�'J�PO7G�BfM�8OLaxEN�DS&LU�&CPR��7LWS�xC�SvTxTE�gS60�FVR�IN�7IHaF�я����� +�=�O�a�s������� ��͟ߟ���'�9� K�]�o���������ɯ ۯ����#�5�G�Y� k�}�������ſ׿� ����1�C�U�g�y� �ϝϯ���������	� �-�?�Q�c�u߇ߙ� �߽���������)� ;�M�_�q����� ��������%�7�I� [�m������������ ����!3EWi {������� /ASew� ������// +/=/O/a/s/�/�/�/ �/�/�/�/??'?9? K?]?o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�_�_�_�_�_	o o-o?oQocouo�o�o �o�o�o�o�o) ;M_q���� �����%�7�I� [�m��������Ǐُ��  Hg552��21��R78�50�J�614�ATUP�7�5457�6�VwCAM�CRI���UIF7�28��N�RE�52v�R6�3�SCH�LI�CƚDOCV�C�SU�8697�0^F�EIOCǛ4��R69v�ESET�W�u�J7u�R68��MASK�PR�XY��7�OCOB��3W����6�3�[J65�536�H$��LCHƪOPLGzW�0�MHCRǪ]S��MCSV�0��{55F�MDSW�v��OP��MPR��t�6�06�PCM���R0E˓�F���6�5�1f�51��0f�P�RS��69�FR�D��FREQ�M�CN�936�SN�BAכ%�SHLB��ME��ּ26�H{TCV�TMIL��6�TPAV�TPT�X��ELړ�6�8�%�#��J95��T�UT��95�UE�V��UECƪUF]R��VCCf�O��wVIP��CSC�ڧCSGƚ$�I�W�EBV�HTTV�Ra6՜��S���CG��{IG��IPGS'��RC��DG��H7.��R66f�5�u�]R��R51f�6�%2�5v�#�J׼�̅6��LU�5�s�v�4v��66F�R64��NVD��R6��R[84�79�4���S5�J76�Du0uFRTS&ڻCR�CRX��CsLI&�e�CMSV�\sV�STY��6�GCTOV�#�V�75�;NN�ORS�����6�FCBV�FCFv��CHV�FCR���FCIF�FC��J�#��G
M��OLn�ENDǪLU��WCPR��Lu�S��C$�StTE�S�60�FVRV�IN��IH���m?? �?�?�?�?�?�?�?O !O3OEOWOiO{O�O�O �O�O�O�O�O__/_ A_S_e_w_�_�_�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o �������� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������� #5GYk}� ������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ}�STD�?LANG�� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ߸�߰���RBT
�OPTN������'� 9�K�]�o�����8������DPN	�� �)�;�M�_�q����� ����������% 7I[m��� �����!3 EWi{���� ���////A/S/ e/w/�/�/�/�/�/�/ �/??+?=?O?a?s? �?�?�?�?�?�?�?O O'O9OKO]OoO�O�O �O�O�O�O�O�O_#_ 5_G_Y_k_}_�_�_�_ �_�_�_�_oo1oCo Uogoyo�o�o�o�o�o �o�o	-?Qc u������� ��)�;�M�_�q��� ������ˏݏ��� %�7�I�[�m������ ��ǟٟ����!�3� E�W�i�{�������ï կ�����/�A�S� e�w���������ѿ� ����+�=�O�a�s� �ϗϩϻ�������� �'�9�K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}���� ����������1�C� U�g�y����������� ����	-?Qc�f�������99��$FE�AT_ADD ?_	���?  	�# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ���������DEMO �y    �L�B�T߁�xߊ߷� ������������G� >�P�}�t����� ��������C�:�L� y�p������������� ��?6Hul ~������ ;2Dqhz� ����� /
/7/ ./@/m/d/v/�/�/�/ �/�/�/�/?3?*?<? i?`?r?�?�?�?�?�? �?�?O/O&O8OeO\O nO�O�O�O�O�O�O�O �O+_"_4_a_X_j_�_ �_�_�_�_�_�_�_'o o0o]oTofo�o�o�o �o�o�o�o�o#, YPb����� �����(�U�L� ^�����������ʏ� ���$�Q�H�Z��� ~�������Ɵ���� � �M�D�V���z��� ����¯ܯ��
�� I�@�R��v������� ��ؿ����E�<� N�{�rτϱϨϺ��� �����A�8�J�w� n߀߭ߤ߶������ ���=�4�F�s�j�|� ������������ 9�0�B�o�f�x����� ����������5, >kbt���� ���1(:g ^p������ � /-/$/6/c/Z/l/ �/�/�/�/�/�/�/�/ )? ?2?_?V?h?�?�? �?�?�?�?�?�?%OO .O[OROdO�O�O�O�O �O�O�O�O!__*_W_ N_`_�_�_�_�_�_�_ �_�_oo&oSoJo\o �o�o�o�o�o�o�o�o "OFX�| �������� �K�B�T���x����� ��ۏҏ����G� >�P�}�t�������ן Ο�����C�:�L� y�p�������ӯʯܯ 	� ��?�6�H�u�l� ~�����Ͽƿؿ��� �;�2�D�q�h�zϔ� �����������
�7� .�@�m�d�vߐߚ��� ���������3�*�<� i�`�r�������� �����/�&�8�e�\� n��������������� ��+"4aXj� �������' 0]Tf��� �����#//,/ Y/P/b/|/�/�/�/�/ �/�/�/??(?U?L? ^?x?�?�?�?�?�?�? �?OO$OQOHOZOtO ~O�O�O�O�O�O�O_ _ _M_D_V_p_z_�_ �_�_�_�_�_o
oo Io@oRolovo�o�o�o �o�o�oE< Nhr����� ����A�8�J�d� n�������яȏڏ� ���=�4�F�`�j��� ����͟ğ֟���� 9�0�B�\�f������� ɯ��ү�����5�,� >�X�b�������ſ�� ο����1�(�:�T� ^ϋςϔ��ϸ����� �� �-�$�6�P�Z߇� ~ߐ߽ߴ��������� )� �2�L�V��z�� �����������%�� .�H�R��v������� ��������!*D N{r����� ��&@Jw n������� //"/</F/s/j/|/ �/�/�/�/�/�/?? ?8?B?o?f?x?�?�? �?�?�?�?OOO4O >OkObOtO�O�O�O�O��O�O__0]  'XF_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?V?h?z?�?�? �?�?�?�?�?
OO.O @OROdOvO�O�O�O�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|� �������� 0�B�T�f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.�  /�)�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |������� ��0�B�T�f�x��� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� \�n������������� ����"4FXj |������� 0BTfx� ������// ,/>/P/b/t/�/�/�/ �/�/�/�/??(?:? L?^?p?�?�?�?�?�? �?�? OO$O6OHOZO lO~O�O�O�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_�_�_�_�_
o o.o@oRodovo�o�o �o�o�o�o�o* <N`r���� �����&�8�J� \�n���������ȏڏ ����"�4�F�X�j� |�������ğ֟��� ��0�B�T�f�x��� ������ү����� ,�>�P�b�t������� ��ο����(�:� L�^�pςϔϦϸ���@���� ��$�4�8�+�N�`�r߄ߖߨ� ����������&�8� J�\�n������� �������"�4�F�X� j�|������������� ��0BTfx ������� ,>Pbt�� �����//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?O O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h� zߌߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N�`�r������� ��������&8 J\n����� ���"4FX j|������ �//0/B/T/f/x/ �/�/�/�/�/�/�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�O�O��O�O�O __$_6Y��$FEAT_DEMOIN  ;T��fP�<PNTI�NDEX[[jQ��NPILECOMP z����Q�iRIU�PSETUP2 {�U��R�  N� �Q�S_AP2B�CK 1|�Y � �)7Xok%�_8o<P�P&oco9U �_�oo�oBo�o�oxo �o1C�og�o� �,�P���� �?��L�u����(� ��Ϗ^�󏂏�)��� M�܏q������6�˟ Z�؟���%���I�[� �������D�ٯh� �����3�¯W��d� �����@�տ�v�� ��/�A�пe����ϛ� *Ͽ�N���r���ߨ� =���a�s�ߗ�&߻� ��\��߀��'��K� ��o���|��4���X� �����#���G�Y��� }������B���f������1�Y�PP�_� 2�P*.VR8���*����0����l PC�>��FR6:�2�V�TzPz��w�]PG���G*.Fo/��	��:,�^/�ST�Mi/�/ /�-M/�/�H�/?�'?p�/�/g?�GIFq?��?�%�?D?V?�?�JPG�?O�%O�?�?�oO�
JSyO�O���5C�OMO%
JavaScript�O�?CS�O&_�&_�O� %Casca�ding Sty�le Sheet�sR_��
ARGN?AME.DT�_��� \�_S_�A�T�_��_�PDISP*�_���To�_�QLa�ZooCLLB.cZIwo2o$ :\�a�\�o�i�ACol�labo�o�o
T�PEINS.XML�_:\![o�Q�Custom T?oolbarbi�PASSWORD�Qo��FRS:\��dB`Passw�ord Config���/��(�e� �������N��r� ����=�̏a���� ��&���J���񟀟� ��9�K�ڟo������� 4�ɯX��|���#��� G�֯@�}����0�ſ ׿f������1���U� �y��ϯ�>���b� ��	ߘ�-߼�Q�c��� ��߽߫�L���p�� �ߦ�;���_���X�� $��H�����~���� 7�I���m���� �2� ��V���z���!��E ��i{
�.�� d����S� wp�<�`� /�+/�O/a/��/ /�/8/J/�/n/?�/ �/9?�/]?�/�?�?"? �?F?�?�?|?O�?5O �?�?kO�?�OO�O�O TO�OxO__�OC_�O g_y__�_,_�_P_b_ �_�_o�_oQo�_uo o�o�o:o�o^o�o �o)�oM�o�o� �6��l��%� 7��[����� ��� D�ُh�z����3� ,�i��������ßR���v������$F�ILE_DGBCK 1|������ �< �)
SUMMARY.DG!��͜MD:U����ِDiag S?ummary�����
CONSLOG���n���ٯ���C�onsole l�og���	TPA'CCN�t�%\������TP Acc?ountin;����FR6:IPKDMP.ZIPͿ�ј
�ϥ���Exception"��ӻ��MEMCHECCK��������-��Memory D�ata����&n{ )��RIPE�p~ϐ�%ߴ�%��� Packet yL:���L�$�c���STAT��߾�� %A�S�tatus��^�	FTP����	���/�mment �TBD2�^� >I�)ETHERN�Ew�
�d�u�﨡?EthernJ�1�?figuraAϩ�~�DCSVRF&����7����� v�erify alyl:��� 4��DIFF/��'���<;�Q�diff��r�|d���CHG01�������A����it�2���270���fx3���I� �p�V�TRNDIAG.�LSu&8����� Ope��L� ~��nostic���T�)VDEV�DAT�������Vis�D�evice�+IMG��,/>/�/:�=i$Imagu/+7UP ES/�/?FRS:\?Z=���Update?s ListZ?���� FLEXEV�EN��/�/�?����1 UIF Ev�M�M���-vZ)�CRSENSP)K�/˞�\!O����CR_TAOR_�PEAKbOͩPS�RBWLD.CM��O͜E2�O\?.�P�S_ROBOWEyLS���:GIG���@_�?d_��Gig�E�(O��N�@��)UQHADOW�__D_V_�_��Sh�adow Cha�nge����dt~�RRCMERR�_��_�_oo��4`CFG Erroro �tailo MA��k�CMSGLIBgoNo`o�o|R�e���z0ic�o�a�)�`ZD0_O�o�s��ZD�Pad��l �RNOT�I�Rd���N?otific����,�AG��P�ӟ t���������Ώ]�� ���(���L�^�폂� �����G�ܟk� ��� �6�şZ��~���� ��C�د�y����2� D�ӯh��������¿ Q��u�
�ϫ�@�Ͽ d�v�Ϛ�)Ͼ���_� �σ�ߧ�%�N���r� ߖߨ�7���[���� ��&��J�\��߀�� ��3����i����"� 4���X���|������ A�����w���0�� =f�����O �s�>�b t�'�K�� �/�:/L/�p/� �/�/5/�/Y/�/ ?�/ $?�/H?�/U?~??�? 1?�?�?g?�?�? O2O �?VO�?zO�OO�O?O �OcO�O
_�O._�OR_ d_�O�__�_�_M_�_ q_oo�_<o�_`o�_ mo�o%o�oIo�o�oo �o8J�on�o� �3�W�{�"� �F��j�|����/��ď֏e������0���$FILE_FR�SPRT  ��������?�MDONL�Y 1|S��� 
 �)MD�:_VDAEXTP.ZZZ1�⏹��ț6%NO� Back fi�le ���S�6P�����>��K�t� ����'���ί]�򯁯 �(���L�ۯp���� ��5�ʿY�׿ Ϗ�$� ��H�Z��~�Ϣϴ� C���g���ߝ�2��� V���cߌ�߰�?��� ��u�
��.�@���d���߈��C�VISB�CKq�[���*.�VD����S�FR�:\��ION\DOATA\��v�S��Vision VD���Y�k��� ��y��B�����x� ��1C��g��� ,�P���� ?�Pu�(� �^��/��M/ �q/�/>/�/6/�/Z/ �/?�/%?�/I?[?�/�??�?2?D?�?9�L�UI_CONFIoG }S���>�; $ �3v�{S�;OMO_OqO�O�O�I#@|x�?�O�O�O __%\�OH_Z_l_~_ �_'_�_�_�_�_�_o �_2oDoVohozo�o#o �o�o�o�o�o
�o. @Rdv��� �����*�<�N� `�r��������̏ޏ �����&�8�J�\�n� �������ȟڟ쟃� ��"�4�F�X�j���� ����į֯���� 0�B�T�f��������� ��ҿ�{���,�>� P�b����ϘϪϼ��� ��w���(�:�L�^� �ςߔߦ߸�����s�  ��$�6�H���Y�~� ������]������  �2�D���h�z����� ����Y�����
. @��dv���� U��*<� `r����Q� �//&/8/�\/n/ �/�/�/;/�/�/�/�/ ?"?�/F?X?j?|?�? �?7?�?�?�?�?OO �?BOTOfOxO�O�O3O �O�O�O�O__�O>_ P_b_t_�_�_/_�_�_ �_�_oo�_:oLo^o�po�o�o$h  �x�o�c�$FLU�I_DATA �~����a�(a�dRES�ULT 3�e�p �T��/wizard/�guided/s�teps/Expert�o=Oas ��������z��Contin�ue with =Gpance�:� L�^�p���������ʏX܏� � �b-�a|�e�0 �0`���c�a?��ps���������ҟ� ����,�>�P��0o w���������ѯ��� ��+�=�O�a�?�1��C�U�e�cllb s�ֿ�����0�B� T�f�xϊϜ�[����� ������,�>�P�b� t߆ߘߪ�i�{��ߟ�:]�e�rip(pſ -�?�Q�c�u���� ����������)�;� M�_�q����������� ����������`��e�#pTimeUS/DST	�� �����!3�E�Enabl (�y������@�	//-/?/Q/�b��)�/M_q24|�/�/??)?;? M?_?q?�?�?Tf�? �?�?OO%O7OIO[O mOO�O�Ob/t/�/�/�Z�"qRegion�O5_G_Y_k_}_�_��_�_�_�_�_�A?merica!�#o 5oGoYoko}o�o�o�o �o�o�o��Ay�O�O�3�O_qEditor�o����������+�=� � �Touch Pa�nel rs (recommenp�)K�������Ə؏�@��� �2�D�|��%��I[qaccesoܟ� ��$��6�H�Z�l�~������Connect �to Network��֯����� 0�B�T�f�x�����x���@��}����,!���s Introduct!_4�F�X�j� |ώϠϲ�������� ��0�B�T�f�xߊ���߮���������  ɿ��"�i�{� ������������� �/�A� �e�w����� ����������+D=�H�3��+� �O�����  2DVhz�K� �����
//./ @/R/d/v/�/�/Yk }�/�??*?<?N? `?r?�?�?�?�?�?�? ��?O&O8OJO\OnO �O�O�O�O�O�O�O�/ _�/1_�/X_j_|_�_ �_�_�_�_�_�_oo 0oBoS_foxo�o�o�o �o�o�o�o,> �O_!_�E_��� ����(�:�L�^� p�����So��ʏ܏�  ��$�6�H�Z�l�~� ��O��s՟����  �2�D�V�h�z����� ��¯ԯ毥�
��.� @�R�d�v��������� п⿡��ş'�9��� `�rτϖϨϺ����� ����&�8���\�n� �ߒߤ߶��������� �"�4��=��a�� Mϲ����������� 0�B�T�f�x���I߮� ��������,> Pbt�E��i� ���(:L^ p��������  //$/6/H/Z/l/~/ �/�/�/�/�/��� �/?�V?h?z?�?�? �?�?�?�?�?
OO.O �ROdOvO�O�O�O�O �O�O�O__*_<_�/ ??�_C?�_�_�_�_ �_oo&o8oJo\ono �o?O�o�o�o�o�o�o "4FXj|� M___q_��_��� 0�B�T�f�x������� ��ҏ�o���,�>� P�b�t���������Ο �����%��L�^� p���������ʯܯ�  ��$�6�G�Z�l�~� ������ƿؿ����  �2��S��w�9��� ����������
��.� @�R�d�v߈�G��߾� ��������*�<�N� `�r��Cϥ�g���� ����&�8�J�\�n� ���������������� "4FXj|� ��������� -��Tfx��� ����//,/�� P/b/t/�/�/�/�/�/ �/�/??(?�1 U??A�?�?�?�?�?  OO$O6OHOZOlO~O =/�O�O�O�O�O�O_  _2_D_V_h_z_9?�? ]?�_�_�?�_
oo.o @oRodovo�o�o�o�o �o�O�o*<N `r������_ �_�_�_#��_J�\�n� ��������ȏڏ��� �"��oF�X�j�|��� ����ğ֟����� 0����u�7����� ��ү�����,�>� P�b�t�3�������ο ����(�:�L�^� pς�A�S�e��ω���  ��$�6�H�Z�l�~� �ߢߴ��߅������  �2�D�V�h�z��� ������������� @�R�d�v��������� ������*;�N `r������ �&��G	�k -�������� /"/4/F/X/j/|/; �/�/�/�/�/�/?? 0?B?T?f?x?7�?[ �?�?�?OO,O>O PObOtO�O�O�O�O�O �/�O__(_:_L_^_ p_�_�_�_�_�_�?�_ �?o!o�OHoZolo~o �o�o�o�o�o�o�o  �ODVhz�� �����
���_ %o�_I�s�5o������ Џ����*�<�N� `�r�1������̟ޟ ���&�8�J�\�n� -�w�Q���ů����� �"�4�F�X�j�|��� ����Ŀ������� 0�B�T�f�xϊϜϮ� ����������ٯ>� P�b�t߆ߘߪ߼��� ������տ:�L�^� p�����������  ��$������i�+� ��������������  2DVh'�� �����
. @Rdv5�G�Y�� }���//*/</N/ `/r/�/�/�/�/y�/ �/??&?8?J?\?n? �?�?�?�?�?��?� O�4OFOXOjO|O�O �O�O�O�O�O�O__ /OB_T_f_x_�_�_�_ �_�_�_�_oo�?;o �?_o!O�o�o�o�o�o �o�o(:L^ p/_������  ��$�6�H�Z�l�+o ��Oo��sou�����  �2�D�V�h�z����� ������
��.� @�R�d�v��������� }�߯����ٟ<�N� `�r���������̿޿ ���ӟ8�J�\�n� �ϒϤ϶��������� �ϯ��=�g�)��� �߲����������� 0�B�T�f�%ϊ��� ����������,�>� P�b�!�k�Eߏ���{� ����(:L^ p����w���  $6HZl~ ���s�������/ ��2/D/V/h/z/�/�/ �/�/�/�/�/
?�.? @?R?d?v?�?�?�?�? �?�?�?OO��� ]O/�O�O�O�O�O�O �O__&_8_J_\_? �_�_�_�_�_�_�_�_ o"o4oFoXojo)O;O MO�oqO�o�o�o 0BTfx��� m_�����,�>� P�b�t���������{o ݏ�o��o(�:�L�^� p���������ʟܟ�  ��#�6�H�Z�l�~� ������Ưد���� ͏/��S��z����� ��¿Կ���
��.� @�R�d�#��ϚϬϾ� ��������*�<�N� `����C���g�i��� ����&�8�J�\�n� �����u������� �"�4�F�X�j�|��� ����q�������	�� 0BTfx��� ������,> Pbt����� ��/����1/[/ �/�/�/�/�/�/�/  ??$?6?H?Z?~? �?�?�?�?�?�?�?O  O2ODOVO/_/9/�O �Oo/�O�O�O
__._ @_R_d_v_�_�_�_k? �_�_�_oo*o<oNo `oro�o�o�ogOyO�O �O�o�O&8J\n �������� �_"�4�F�X�j�|��� ����ď֏�����o �o�oQ�x������� ��ҟ�����,�>� P��t���������ί ����(�:�L�^� �/�A���e�ʿܿ�  ��$�6�H�Z�l�~� �Ϣ�a����������  �2�D�V�h�zߌߞ� ��o��ߓ��߷��.� @�R�d�v����� ��������*�<�N� `�r������������� ����#��G	�n �������� "4FX�|� ������// 0/B/T/u/7�/[ ]/�/�/�/??,?>? P?b?t?�?�?�?i�? �?�?OO(O:OLO^O pO�O�O�Oe/�O�/�O �O�?$_6_H_Z_l_~_ �_�_�_�_�_�_�_�?  o2oDoVohozo�o�o �o�o�o�o�o�O_�O %O_v���� �����*�<�N� or���������̏ޏ ����&�8�J�	S -w���cȟڟ��� �"�4�F�X�j�|��� ��_�į֯����� 0�B�T�f�x�����[� m����󿵟�,�>� P�b�tφϘϪϼ��� ���ϱ��(�:�L�^� p߂ߔߦ߸�������  ￿ѿ�E��l�~� �������������  �2�D��h�z����� ����������
. @R�#�5�Y� ���*<N `r��U���� �//&/8/J/\/n/ �/�/�/c�/��/� ?"?4?F?X?j?|?�? �?�?�?�?�?�??O 0OBOTOfOxO�O�O�O �O�O�O�O�/_�/;_ �/b_t_�_�_�_�_�_ �_�_oo(o:oLoO po�o�o�o�o�o�o�o  $6H_i+_ �O_Q�����  �2�D�V�h�z����� ]oԏ���
��.� @�R�d�v�����Y�� }ߟ񟵏�*�<�N� `�r���������̯ޯ 𯯏�&�8�J�\�n� ��������ȿڿ쿫� ��ϟ�C��j�|ώ� �ϲ����������� 0�B��f�xߊߜ߮� ����������,�>� ��G�!�k��Wϼ��� ������(�:�L�^� p�����S߸�������  $6HZl~ �O�a�s�����  2DVhz�� ������
//./ @/R/d/v/�/�/�/�/ �/�/�/���9?� `?r?�?�?�?�?�?�? �?OO&O8O�\OnO �O�O�O�O�O�O�O�O _"_4_F_??)?�_ M?�_�_�_�_�_oo 0oBoTofoxo�oIO�o �o�o�o�o,> Pbt��W_�{_ ��_��(�:�L�^� p���������ʏ܏� ��$�6�H�Z�l�~� ������Ɵ؟꟩� �/��V�h�z����� ��¯ԯ���
��.� @���d�v��������� п�����*�<��� ]����C�EϺ����� ����&�8�J�\�n� �ߒ�Q����������� �"�4�F�X�j�|�� Mϯ�q�������� 0�B�T�f�x������� ��������,> Pbt����� �������7��^ p�������  //$/6/��Z/l/~/ �/�/�/�/�/�/�/?  ?2?�;_?�?K �?�?�?�?�?
OO.O @OROdOvO�OG/�O�O �O�O�O__*_<_N_ `_r_�_C?U?g?y?�_ �?oo&o8oJo\ono �o�o�o�o�o�o�O�o "4FXj|� ������_�_�_ -��_T�f�x������� ��ҏ�����,��o P�b�t���������Ο �����(�:��� ��A�����ʯܯ�  ��$�6�H�Z�l�~� =�����ƿؿ����  �2�D�V�h�zό�K� ��o��ϓ���
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ������#���J�\�n� ���������������� "4��Xj|� ������ 0��Q�u7�9� ����//,/>/ P/b/t/�/E�/�/�/ �/�/??(?:?L?^? p?�?A�?e�?�?�/  OO$O6OHOZOlO~O �O�O�O�O�O�/�O_  _2_D_V_h_z_�_�_ �_�_�_�?�?�?o+o �?Rodovo�o�o�o�o �o�o�o*�ON `r������ ���&��_/o	oS� }�?o����ȏڏ��� �"�4�F�X�j�|�; ����ğ֟����� 0�B�T�f�x�7�I�[� m�ϯ������,�>� P�b�t���������ο �����(�:�L�^� pςϔϦϸ����ϛ� ����!��H�Z�l�~� �ߢߴ����������  �߿D�V�h�z��� ����������
��.� �����s�5ߚ����� ������*<N `r1����� �&8J\n �?��c������ /"/4/F/X/j/|/�/ �/�/�/�/��/?? 0?B?T?f?x?�?�?�? �?�?��?�O�>O PObOtO�O�O�O�O�O �O�O__(_�/L_^_ p_�_�_�_�_�_�_�_  oo$o�?EoOio+O -o�o�o�o�o�o�o  2DVhz9_� �����
��.� @�R�d�v�5o��Yo�� ͏����*�<�N� `�r���������̟� ���&�8�J�\�n� ��������ȯ��я�� ����F�X�j�|��� ����Ŀֿ����� ݟB�T�f�xϊϜϮ� ����������ٯ#� ��G�q�3��ߪ߼��� ������(�:�L�^� p�/ϔ���������  ��$�6�H�Z�l�+� =�O�a���������  2DVhz�� ������
. @Rdv���� �������/��</N/ `/r/�/�/�/�/�/�/ �/??�8?J?\?n? �?�?�?�?�?�?�?�? O"O��/gO)/�O �O�O�O�O�O�O__ 0_B_T_f_%?w_�_�_ �_�_�_�_oo,o>o Poboto3O�oWO�o{O �o�o(:L^ p������o�  ��$�6�H�Z�l�~� ������Ə�o珩o� �o2�D�V�h�z����� ��ԟ���
��� @�R�d�v��������� Я�����׏9��� ]��!�������̿޿ ���&�8�J�\�n� -��Ϥ϶��������� �"�4�F�X�j�)��� M����߅������� 0�B�T�f�x���� ���������,�>� P�b�t���������{� �ߟ�����:L^ p�������  ��6HZl~ �������/ ����;/e/'�/�/ �/�/�/�/�/
??.? @?R?d?#�?�?�?�? �?�?�?OO*O<ONO `O/1/C/U/�Oy/�O �O__&_8_J_\_n_ �_�_�_�_u?�_�_�_ o"o4oFoXojo|o�o �o�o�o�O�O�O	�O 0BTfx��� ������_,�>� P�b�t���������Ώ ������o�o�o[� ��������ʟܟ�  ��$�6�H�Z��k� ������Ưد����  �2�D�V�h�'���K� ��o�Կ���
��.� @�R�d�vψϚϬϾ� Ͽ������*�<�N� `�r߄ߖߨߺ�y��� ������&�8�J�\�n� ������������� ���4�F�X�j�|��� �������������� -��Q���� ����,> Pb!������ ��//(/:/L/^/ /A�/�/y�/�/  ??$?6?H?Z?l?~? �?�?�?s�?�?�?O  O2ODOVOhOzO�O�O �Oo/�/�/�O_�/._ @_R_d_v_�_�_�_�_ �_�_�_o�?*o<oNo `oro�o�o�o�o�o�o �o�O_�O/Y_ �������� �"�4�F�X�o|��� ����ď֏����� 0�B�T�%7I�� mҟ�����,�>� P�b�t�������i�ί ����(�:�L�^� p���������w����� ����$�6�H�Z�l�~� �Ϣϴ��������ϻ�  �2�D�V�h�zߌߞ� ����������
�ɿۿ �O��v����� ��������*�<�N� �_������������� ��&8J\� }?�c����� "4FXj|� ������// 0/B/T/f/x/�/�/�/ m�/��/�?,?>? P?b?t?�?�?�?�?�? �?�?O�(O:OLO^O pO�O�O�O�O�O�O�O  _�/!_�/E_?	_~_ �_�_�_�_�_�_�_o  o2oDoVoOzo�o�o �o�o�o�o�o
. @R_s5_��mo �����*�<�N� `�r�������gȍޏ ����&�8�J�\�n� ������c��џ�� �"�4�F�X�j�|��� ����į֯������ 0�B�T�f�x������� ��ҿ�������ٟ#� M��tφϘϪϼ��� ������(�:�L�� p߂ߔߦ߸�������  ��$�6�H���+� =ϟ�a����������  �2�D�V�h�z����� ]���������
. @Rdv���k��}�����$FM�R2_GRP 1���� ��C4  B]��	 ��9�K6F@ a@��6G�  �Fg�fC�8R�y?�  ��6�6�X���87�5t��5����5`+�yA�  /+BH�w-%O@S339%�5[/l-6@6!�/xl/ �/�/�/�/?�/&?? J?5?G?�?k?�?��_CFG ��TK�?�? OO�9N�O 
F�0FA K@�<RM_�CHKTYP  ���$&� R{OMa@_MINg@������@�R X�SSB�3��? 7�O���C�O�O�5TP_�DEF_OW  ���$WIRC�OMf@_�$GE�NOVRD_DO2�F��E]TH��D� dbUdKT_EN�B7_ KPRAV�C��G�@ ��Y�O�_�?oy�o&oI* �QOUU�NAIRI<�@��o`Go�o�o�o��C�p�3��O:��B��+sL�i�O�PSMT��Y(�@
t�$HOSTC�2s1��@��5 MC��R{����  27�.00�1�  e�]�o�������K��ď֏��������	�anonymou�s!�O�a�s����� �4�������� D�!�3�E�W�i����� ����ï柀�.��� /�A�S���课�П�� ��Ŀ����+�r� O�a�sυϗϺ��� ������'�n����� ���ϓ�ڿ�������� ��F�#�5�G�Y�k�� �υ����������B� T�f�C�z�g��ߋ��� ���������	- P�����u���� ��(�:�<)p�M _q������� �/$ZlI/[/m/ /�/����//�/ D!?3?E?W?/?�? �?�?�?�/�?./OO /OAOSO�/�/�/�/�? �O?�O�O__+_r? O_a_s_�_�_�O�?O��_�_oo'o�t�qE�NT 1�hk sP!�_no  �p\o�o�o�o�o�o�o �o�o:_"� F�j����� %��I��m�0���T� f�Ǐ��돮��ҏ3� ��,�i�X���P���t� ՟��៼�
�/��S� �w�:���^�������������ܯ=� �Q�UICC0J�&�!�192.168�.1.10c�X�1 ��v�8��\�2�ƿ�ؿ9�!ROUT3ER:��!��a�~�PCJOG�Ͼe�!* ��0���U�CAMPRT��϶�!�����R�TS���x� !�Software� Operator PanelU������7kNAME �!Kj!ROB�O����S_CFG� 1�Ki ��Auto-started�D/FTP�Oa�O �_���O���������� E_�.�@�R�u�c�	� ����������cN:�L� ^�;r���R��� �����%H �[m���jO |O�O�O4!/hE/W/ i/{/�/T�/�/�/�/ �//�//?A?S?e?w? �?����??�?</ O+O=OOO?sO�O�O �O�O�?`O�O__'_ 9_K_�?�?�?�?�O�_ �?�_�_�_o#o�OGo Yoko}o�o�_4o�o�o �o�of_x_�_g �o��_�����o ��-�?�Q�tu�� ������Ϗ�(:L ^`�2��q������� ����ݟ���%�H� ʟ[�m���������� � �ί4�!�h�E�W� i�{���T���ÿտ� 
�Ϟ�/�A�S�e�w�����_ERR ��ڇϗ�PDUS_IZ  �^6�����>��WRD� ?(���� � guest���+�=�O�a����SCD_GRO�UP 3�(� �,�"�IFT��$�PA��OMP��� ��_SH��E�D�� $C��CO�M��TTP_AU�TH 1��� �<!iPend�anm�x�#�+!KAREL:*x����KC��������VISION SET��(����?�-�W�R���v��� ��������������G�CTRL ����a�
�F�FF9E3���FRS:DEFA�ULT�FA�NUC Web ?Server�
t dG����/� �2DV��WR_C�ONFIG �.��������IDL_CPU_kPC� �B����� BH�MIN�����GNR_I�O������ȰHM�I_EDIT =���
 ($/C/ ��2/k/V/�/z/�/�/ �/�/�/?�/1??U? @?y?d?�?�?./�?�? �?�?OO?OQO<OuO `O�O�O�O�O�O�O�O�__;_�NPT_�SIM_DO��*NSTAL_S7CRN� �\UQ�TPMODNTOqL�Wl[�RTYbXp�qV�K�ENB�W��ӭOLNK 1�����o%o7o�Io[omoo�RMAS�TE��Y%OSLAVE �����eRAMCACH�E�o�ROM�O_CcFG�o�S�cUO'���bCMT_OPp�  "��5sYCL�o�u� _ASG 19����
 �o� ������"�4��F�X�j�|����kwrN�UM����
�bI�P�o�gRTRY_�CN@uQ_UP)D��a��� �bp�b��n��M��а�P}T?��k ��._������ɟ۟� �S���)�;�M�_�q�  �������˯ݯ�~� �%�7�I�[�m���� ����ǿٿ�����!� 3�E�W�i�{�
ϟϱ� �������ψϚ�/�A� S�e�w߉�߭߿��� ������+�=�O�a� s���&�������� ����9�K�]�o��� ��"����������� ����GYk}�� 0����� CUgy��,> ���	//-/�Q/ c/u/�/�/�/:/�/�/ �/??)?�/�/_?q? �?�?�?�?H?�?�?O O%O7O�?[OmOO�O �O�ODOVO�O�O_!_ 3_E_�Oi_{_�_�_�_ �_R_�_�_oo/oAo �_�_wo�o�o�o�o�o `o�o+=O�o s�����\n ��'�9�K�]�����������ɏۏi�c�_�MEMBERS �2�:� �  $:� ����v���1���R�CA_ACC 2��� �  [}�� �:�2 Y �p )5�l��(l�l���� ����� {���a�B�UF001 2��n�= ��?�?  ��=��=�  �>�>�V��=8{=8��=�=����?H?H.�V�>(>����
����=�=�  ��@�@�N�VK�0K0  � *�*��@
����@�@m��j��u�0u]��8=�=}���x?�?؆��J�����8H�����xX�XM������K�L��8���Mu08�<x��[��u0�iڤu�ڤ�ڤ�ڤ�ڤ��ڤ�ڤ�ڤ�ڤ��ڤ�ڤ�ڣ�Zn�Z�	���J�U�J��J��J��J���ڣ�z�z��z�*z�Vu0?�5@��=�=U���I����V���������X�X�����ߙ2���� "�4�F�X�j�|����� ��ĭ��ء������ ������������	� ��������!���)� ��1���9���@�B�H� ��P�U�Y�U�a�U�i� U�q�U�y������҉� �ґ��ҙ��ҡ��ҩ���Ϳ߿�3���l� �l���"��*�� 2�l�9�>�B�>�J�>� R�l�Y�^�b�l�i�n� r�n�z�n��n��l� �����������l� �����������T�ƣ ��Ѡ��٢������� �������	����� '���)�7���9�G�l� H�W�V�Y�g�V�i�w� V�y��ӎ򉲗ӎ� �ӎ�Ў�[������� ��������������~a�CFG 2�n�� 4l��
l�
l�<l�47%�a��HIS钜n� ��� 2025�-11-29l� 珚�������l�;g� � % �� � -i�B�� �r������ �//K]J/\/n/ �/�/�/�/�/�/�/#/ 5/"?4?F?X?j?|?�? �?�?�?�/?�?OO 0OBOTOfOxO�O�O�? �?�?�O�O__,_>_ P_b_t_�_�O�O�_�_ �_�_oo(o:oLo^o L	��[m�o�o�o@�o�o!3!: Ic��Ƒd��@d�_ �_<������ ��+��_t�s��� ������͏ߏ��� L�^�K�]�o������� ��ɟ۟�$�6�#�5� G�Y�k�}�������ů �������1�C�U� g�y�����ԯ���� ��	��-�?�Q�c�u� coue�Ѐo�o�o���� ���"�4�F�X�!o� F�}Ӳ�Ŀa��� ��������,�>�P� �ߙ߫ߘ������� ����(�:�q��p� ��������������  I�[�HZl~� �����!3  2DVhz��� ��
//./@/�R/d/v/�/�/��u`I_CFG 2���� H
Cycle Time��Busy�I�dl�"�minz�+1Up�&��Read�'�Dow8? �2�#Count>�	Num �"�����<��~�qaP�ROG�"�������)/sof�tpart/ge�nlink?cu�rrent=me�nupage,1133,1�/OO�/OAO3b5leSDT�_ISOLC  ���� �@�.J�23_DSP_ENB  vK0�@?INC ��M����@A   ?� � =���<#��
�A�I:�o ��A__���O<_�GOB�0C�C5�FVQ�G_GROUP �1�vK<Zq<���C��_D_?"��?�_��Q�_o .o@o�_dovo�o�o��,_NYG_IN_�AUTOcT�MPO�SRE^_pVKANJI_MASK v��HqRELMONG ��˔?��y_o x�����.6r�3%��7�C���u�o��DKCL_L�`N�UM�@�$KEYLOGGING�����Q�E�0LAN�GUAGE ���~��DE?FAULT �����LG�!��:2e���x�@{�80oH  ���'0��� 
������|GOUF ;��
��(UT1:\��  �-�?�Q�h� u���������ϟ������(g4�8i�N_DISP ��O�8�_�_��LOCT3OL����Dz|�A��A��GBOOK ���d�1
�
�۠X����#�5��G�Y�i���3{�W�	��쉞QQJ¿Կ1���_BUFF ;2�vK ����25
�ڢVB&�7� Collaborativ�=�O� �ώϠϲ��������� '��0�]�T�fߓߊ�����DCS � �9�B�Ax�����%��-�?�Q���IO 2��� ���Q��������� ����*�<�N�b�r� ���������������&:e�ER_ITMsNd�o��� ����#5G Yk}�����p����hSEV���MdTYPsN��c/u/�/
-�aRS�T5���SCRN__FL 2�s��0����/??1?C?U?�g?�/TPK�sOR">��NGNAM�D���~�N�UPS_AC�R� �4DIGI��8+)U_LOA�D[PG %�:%�T_NOVIC�Et?��MAXUA�LRM2��1���2�E
ZB�1_P�5�0� ��y�Z@CY���˭�O+���ۡ�D|PPw 2�˫ ��	R/_
_C_._g_y_ \_�_�_�_�_�_�_�_ oo?oQo4ouo`o�o |o�o�o�o�o�o) M8qTf�� �����%��I� ,�>��j�����Ǐُ �����!���W�B� {�f�������՟���� ܟ�/��S�>�w��� l�����ѯ��Ư�� +��O�a�D���p����RHDBGDEF ���E�ѱO��_L?DXDISA�0�;�c�MEMO_AP޻0E ?�;
 ױ��3�E�W�i��{ύϟϱ�Z@FRQ_CFG ��Gm۳A ��@�����<��d%�� ���t���B��K���*i�/k� **:tҔ�g�y�� ���߱��������� �J�Es�J d������,(H���[� ����@�'�Q�v�]� ���������������*NPJISC 31��9Z� ���� ��ܿ�����	Z�l_MSTR ��#-,SCD 1�"͠{��� �����//A/ ,/e/P/�/t/�/�/�/ �/�/?�/+??O?:? L?�?p?�?�?�?�?�? �?O'OOKO6OoOZO �O~O�O�O�O�O�O_ �O5_ _Y_D_i_�_z_ �_�_�_�_�_�_o
o oUo@oyodo�o�o�o �o�o�o�o?*�cN�MK���;љ$MLT�ARM���N��r ��հ��>İMETPU��zr���CNDSP?_ADCOL%�ٰ�0�CMNTF� �9�FNb�f�7�FS�TLI��x�4 �;ڎ�s����9�_POSCF��q��PRPMe��STvD�1�; 4�#�
v��qv����� r��������̟ޟ � ��V�8�J���n����¯�������9�SI�NG_CHK  }��$MODA����t�{�~2�DE�V 	�	M�C:f�HSIZE���zp�2�TASK� %�%$12�3456789 �ӿ�0�TRIG ;1�; lĵ��2ϻ�!�bϻ�YP蠱��H�1�EM_�INF 1�N��`)AT&F�V0E0g���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ��2�ԁH6�^���Rφ��A��߶�q��������  ��5������ߏ�B� ������������1� C�*�g��,��P�b� t������R�?�� �u0������ ���������M q ���Z���/ �%/��[/ 2 �/�/h�//�/�/� 3?�/W?>?{?�?@/�? d/v/�/�/O�//OAO x?eO?�ODO�O�O�O|�O_�NITORÀ�G ?z�   	EXEC1~s�&R2,X3,X4,X5�,X��.V7,X8,X9~s'R�2�T+R�T7R �TCR�TOR�T[R�TgR��TsR�TR�T�R�S2��X2�X2�X2�X2��X2�X2�X2�X2��X2h3�X3�X3�7R2�R_GRP_�SV 1��� �(�=�ĝ<����=�9P�w�п����3jca���_D�B��~�cION_DB<���@�zq  �J2p<2p=Y�1u�2p��>w�ZpyZpz�Y��@N   �Xrp]p@yq$�rY�-ud1������8�PG_JOG� �ʏk�
�2��:�o�=���?����@0�B��~\�n���������H�?��C�@�pŏ׏���  ������qL_NAM�E !ĵ8���!Defaul�t Person�ality (from FD)qp�0�RMK_ENOgNLY�_�R2�a� 1�L�XL��8�gpl d����şן���� �1�C�U�g�y����� ����ӯ���	��n� 
�<�N�`�r�������p��̿޿� :� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w���������������+��<�Se w�������x��A�a��AB�Bw��Pf ������/!/ 3/E/W/i/{/�/�/�/ ���/�/??/?A? S?e?w?�?�?�?�?�? �?�?�/�/+O=OOOaO sO�O�O�O�O�O�O�O __'_9_&O�S��#�x_�]�rdtS�� �_�]�_�_�W�����S�"oe_oXoa  ��qogoyo�o�o�o�o@�ouP�p"|����	`[oUgy8qK��A\����s� AA ��y@h�Q�Q��e"���Tk\$���  ��P��PE�xC�  �I�@oa�<o��p��� ����ߏ
f�Q,�������0��PCr� �� 3r �.� �@D�  A�?��G�-�?.I�.@I��A����  ;��	lY�	 ��X  ������� �,? � ������uPK�o������]K��K]�_K	�.��w��r_	����@
��)�b�1�����I��Y�����T;�fY�{S���3����I�>J���;�Î?v�>��=�@�����E��R ѯעZ���wp��u��� D!�3���7pg  �  ��9�͏W���	'�� � u�I�� �  ���u��:�È��ß�=��ͱ���@��ǰ�3��{"3�E�&���N�pC�  'Y�&�Z�i�bb�@f�i�n�C��D��I�C����b��r���`����B�p�Ŕq���}ر�.DzƏ<ߛ�`�pK�pߖ����������А G4P����.z���d  �Pؠ?�ff�_��	��C 2p>�P���8.f�t�>L���U���	(.��P���٨������É��� x��;�e�m��KZ;��=g;�4�<�<����%�G���3����p?fff�?ذ?&S���@{=0e�?��q� �y�rN�Z���I���G� ��7���(�����! E0iT�����x��F�p��� #��D��w� ������// =/(/a/L/�/p/��/ �p�6�/Z#?�/ ? Y?k?}?��?�?>?�?��?�?�?�?1O�����KD�y{CO�OO�O���ذO�O�O�O�y���J��}�D#D1���.�D��@�A�mQa��9N,ȴA�;�^@��T@�|j@$�?��V�>�z������=#�
>�\)?��
=��G�-]�{�=���,��C+��Bp���P���6��C98R����?N@���(��5-]G��p�Gsb�F��}�G�>.E�VD�Kn����I�� F��W�E��'E���D��;n����I��`E��G��cE�vmD���-_ �oQ_�o�o�o �o$ H3X~i�� �������D� /�h�S���w������� �я
���.��R�=� v�a�s�����П���� ߟ��(�N�9�r�]� ��������ޯɯۯ� ��8�#�\�G���k��� ����ڿſ���"�� F�1�C�|�gϠϋ���@����������P(�Q�34�] ������Q�	�9�Oߵ53~�qmm��aҀ5Q����aғ����ߵ1�������1��U�C�y�g��%P�P���!�/��'���
�x��.������4� ;�t�_����������� ����:%��/0�/d����� ���7%[@Im���027�  B�S@J@�KCH#PzS@�0@ZO /1/C/U/g/y/�-�#��/�/�/�/�/�3�?�3�� @�3J��0�0�13��5
 ?f?x? �?�?�?�?�?�?�?O�O,O>OPO�Z@1 ����ۯ�c/�$�MR_CABLE� 2ƕ� ��TT�����ڰO ���O�Y�@���C_�� ��_O_u_7_I__�_ �_�_�_�_o�_�_o Koqo3oEo{o�o�o�o �o�o�o�o�oGm /�K!�"���O� ���ذ�$�6���w*Y�** �C�OM ȖI�����":&�%�% 234567O8901���� ��HÏ��� � !� ��!
���M�not sent� b��W���TESTFECS�ALGR  egD)
!d[�41�
k�������$pB����������� 9U�D1:\main�tenances�.xmlğ�  �C:�DEF�AULT�,�BGR�P 2�z�  ����%  �%!�1st clea�ning of cont. v��ilation +56��ڧ�!0�����+B��*������+��"%��me�ch��cal c�heck1�  ��k�0u�|�� ԯ����Ϳ߿�@���?rollerS�e�w�ū��m�ϑϣ����@�Basic� quarterCly�*�<�ƪ,\��)�;�M�_�q�8�MXJ��ߓ "8��� ���ߕ �����+�=��C�g�ߋ���߹���������@�Overha�u�ߔ��?� x� I�P����}���������� $n���� ��aIl�ASew� ����� � +=O�s��� ����/R�9/ �(/��/�/�/�/�/ /�/�/N/#?r/G?Y? k?}?�?�/�???�? 8?OO1OCOUO�?yO �?�?�O�?�O�O�O	_ _jO?_�O�Ou_�O�_ �_�_�_�_0_oT_f_ ;o�__oqo�o�o�o�_ �oo,oPo%7I [m�o��o�o� ���!�3��W�� ������ÏՏ�6� ���l����e�w��� ������џ�2��V� +�=�O�a�s���� ��ͯ����'�9� ��]�������⯷�ɿ ۿ���N�#�r���Y� ��}Ϗϡϳ������ 8�J��n�C�U�g�y� ���ϯ������4�	� �-�?�Q��u����� �ߞ���������f� ;������������ �����P���t�I [m����� �:!3EW� {��� ��� //lA/��w/���/�/�/�/�/X*�"	� X�/?.?@?�)B a/o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�_�_�_�_�_	o�o" Џ!?� ; @�! M?Ho Zolo�&4o�o�o�o�(�*�o** F�@ i!k&�`o�'9�o]o�����/^&�o��� ��/�A�S�e��� #�����я����� +�q�����7������� k�͟ߟ��I�[��� K�]�o���C�����ɯ���o$�!�$M�R_HIST 2��g%#�� 
 �\7"$ 2345?6789013�;���b2�90/���� [���./����ǿٿ F�X�j�!�3ρϲ��� {��ϟ�����B��� f�x�/ߜ�S����߉� �߭��,���P��t����=��$�SKCFMAP  g%�&��b
�� ����ONREL  �$#�������EXCFENB��
����&�FNC�-��JOGOVL�IM�d#�v���K�EY�y���_�PAN������R�UNi�y���SFSPDTYPM�<���SIGN���T1MOTk�����_CE_GRP7 1�g%��+� 0�ow�#d�� ����&�6 \�7y�m� ��/�4/F/-/j/ !/t/�/�/�/{/�/�/�/?�+��QZ_E�DIT
����TC�OM_CFG 1����0�}?�?�? }
^1SI �NB����?�?���?�$O����?XO78T__ARC_*��X�T_MN_MO�DE
�U:_S�PL{O;�UAP_�CPL�O<�NOCHECK ?��/ �� _#_ 5_G_Y_k_}_�_�_�_��_�_�_�_oo��N�O_WAIT_L�	S7> NTf1�����%��qa_ERMRH2������� ?o�o�o�o��O�Gj�@O�cӦm| �:�6GA@g���A����PF������W/�-`���<���?���)��n�b_PARAM�b����vHO��w
�.�@� = n�]�o� w�Q�����������`Ϗ�)���w�[��m� �����ODRD�SP�C8�OFFSET_CARI0��OǖDISԟœS;_A�@ARK
T9�OPEN_FIL�E��1T6�0OPTION_IO�����K�M_PRG ;%��%$*�����'�WO��N�s�ǥ�� ���u����	� ����Ӧ������RG_DSBL'  ����jN����RIENTTO����C�����A� ��U�@IM_D�S���r��V��LCT �{mP2ڢȪ3̹��dҩ��_P�EX�@���RAT��G d8��̐UOP װ�:�����S�e�Kωϗ��$��r2G�L�X�LȚ�l 㰂�������'�9� K�]�o߁ߓߥ߷��� �������#�5�G���2��v������� ������e�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?�q1�~?�?�?�? �?�?�?�?O O2ODO^�yA�a�m? ~N��~O�O�P�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�O �Oo$o6oHoZolo~o �o�o�o�o�o�o�o  �_oVhz�� �����
��.��@�R�d�QOES��(����B�d�ӏ� ʏ��������Y�D�}�0��r������� ��ԟڟ���p���=�4M��q�	`����x����c�:�o��¯ԯ����A�C  �k�C�C�ڰe"ڰ���O���  ����-���)�C�  �t�k���g�����Կ ��ѿ
�5���^:�ĳ��OU��� �� �H��n��� � ^��\� @D�  &p�?�v�\�?:px��:qC4r�p�(�� � ;�	l��	 ��X � ������ ��, � �x������Hʪ�������H���Hw�zH����ϝ�8�B���B��  Xѐ�`�o�*��'3����t�>u����fC{ߍ��:pB\��
�Ѵ9:qK�t�� �����$���*��� D�P�^��b�g  �  �h������)�	'� �� ��I� ��  ��'�=��������t�@����!�b��^;bt�U�(�N��r� ' '��E�C�И�t�C�И��ߗ���jA��@�����%�B �� ��,���H:qDz�k�ߏz����������А 4P���:uz:���	�f��?�faf'�&8� ]��m�8:p��>!L�����$�(:p�P��	������:�� x�;e�m�"�KZ;�=g�;�4�<<�0��E/Tv��b����?fff?�?y&� )�@=0�%?��%`9��}! ��$�x��/v��/f'�� W,??P?;?t?_?�? �?�?�?�?�?O�?(O OLO�/�/�/EO�OAO �O�O�O�O_�O_H_ 3_l_W_�_{_�_�_1� �_A���eO+o�ORoo Oo�o�o�oK/�o�omo �o*'`+�,�zt���CL�H<��}?����X�
������u�����D1�/n�t�x�p�q��@I�h~�,ȴA;�^@���T@|j@�$�?�V�n��z�ý��=�#�
>\)?��
=�G�����{=��,���C+��B�p����6���C98R����?}p��(��5���G�p�G�sb�F�}�G��>.E�VD��KL����I��� F�W�E���'E���D���;L����I���`E�G���cE�vmD���\�՟��ҟ� ��/��S�>�w�b��� ����ѯ������� =�(�:�s�^������� ��߿ʿ�� �9�$� ]�Hρ�lϥϐϢ��� ������#��G�2�W� }�hߡߌ��߰����� ���
�C�.�g�R�� v��������	��� -��Q�<�u�`�r��� ����������'�M�(�34�]O!���8h~�%3~�m���ǀ5Q��������!���   `N�r��J	eP@"P��Q�_�/V/9/$/]/H)����c/j/�/�/�/ �/�/�/�/!??E?0? i?T?"&�_�_�?�?�8��?�?O�?OBO 0OfOTO�OxO�O�O�O��O2f?_  B���pY�$QCHR�z�p@�N_`_r_�_�_�_�]c�O�_�_0oo+o?�Bc�� @d4��QJc�D
 2o�o�o�o�o�o�o %7I[m���oa ������c/�$PARA�M_MENU ?� � � DEF�PULSE��	�WAITTMOU�T�{RCV� �SHELL_�WRK.$CUR�_STYL�p�"�OPT8Q8�PT�BM�G�C�R_DECSN�p�V<�� ���������-�(� :�L�u�p��������q�SSREL_ID�  ��̕U�SE_PROG �%�z%���͓C�CR�pޒ��s1�_HOST !�z#!6�s�+�T�=����V�h���˯*�_�TIME�rޖF�~�pGDEBUGܐ��{͓GINP_F�LMSK��#�TR\2�#�PGAP� ���_b�CH1�"�TWYPE�|�P�� ������0�Y�T� f�xϡϜϮ������� ���1�,�>�P�y�t� �ߘ��߼�����	�� �(�Q�L�^�p��%�WORD ?	�{
 	PR��p#MAI��q"3SUd���TE��p#��	1���COL�n%��!���L�� �!��F�d�T�RACECTL �1� �q }�� �#�����_�DT Q�� ��z�D �� �La ��k`����������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_�T� �_�_�_ �W��Uoo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�.�oP�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/Dϒ/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D��V�h�z�����������$PGTRACE�LEN  �� � ������Ά_UP _�����������΁_CFoG ����*��
���*�*�D��O���O�  ��O��DEFSPD� ��������΀H_CONF�IG ����� ����dĔ�&݂ ��ǑP^�a�l㑹��΀IN�?TRL ��=��8^���PE��������*�ÑO��΀LID���	~T�LLB 1ⳙ_ ��BӐsB4��O� �𼧶��Q� <<7 ��?��� ����M�3�U���i� ��������ӿ��	�7�T�Ϣk�b�tϡπ诚��������S�G�RP 1爬����@A!���4�I���A �C�u�C�OCWjVF�/��Ȕ`a�zي�ÑÐ�t�0�ޯs���´�ӿ���B������������A�S�&�B3�4�_������j���������	� B�-���Q���M�������  Dz����.� ����&L7p[ ��������6!Zh)w�
V7.10be�ta1*�Ɛ@��*�@�) @ߺ+A Ē?���
?fff>�����B33�A�Q�0�B(���A���AK��h����//('/9/P�p*�W�ӑ��n/�/�%���R��fh���� *���P2�LR��/�/@�/�/�/H?�Ĕ�I�u�&:���?��x?��?A���P!\3 Bfu�B��?�5BH�3�[4��o��4�I�[45��/B\3x3Dx�?YO�?aOkO}O�<<�R@��O�C�O�O��O�O�DA�X�KNO?W_M  Z�%��X�SV 賚ڒ���_�_�_?��_�_�_o����W�M�+�鳛 ��	~<�3#���_��o�\=��
]bV4�@u��u��e��o�l,�X�MR+��JmT3?��W�1C{��OADBANFW�DL_V�ST+�1 k1����P4C� ��[��i/��� ��?�1�C���g�y� �������ӏ�*�	�@�`�?�Q�c��w2�|8Va�up�<ʟ����p3��Ɵ؟Ꟃw4 ��+�=��w5Z�l�~����w6����ѯ㯂�w7 ��$�6��w8`S�e�w����wMAmp�������OVL/D  ��yo���rPARNUM � �{+þ�?υqS[CH�� �
��pX���{s��UPDX��)ź��Ϧ�_CMPa_@`���p|P'yu~�ER_CHK���yqbb3��.��RSpp?Q_MO�m��_}ߥ�_REWS_G�p쩻
� e�����0�#�T�G�x� k�}��������������׳�������� �:�Y�^���Y�y��� ���Ӭ����������� ����R�6UZ��ӥ�u����V �1�FvpVa@k��p��THR_ICNRp��(byudoMASS Z)�MNGMON_�QUEUE �P�uyvup\!��N��UZ�NW��ENqD��߶EXE�����BE���O�PTIO��ۚP�ROGRAM %z%��~Ϙ?TASK_I��.OCFG �zx+�n/� DATACcM�+�1#s2ae ?"?4?F?X??|?�? �?�?�?o?�?�?OO^�/INFOCc��-���?wO�O�O�O�O �O�O�O__+_=_O_ a_s_�_�_�_�_�_�_4:GFD��, 	��!6��K_�!�)fN!fENB��0m��Pfi2YokhG�!2�0k X,		d�o=��·o���e�a$�pd��i�i�g�_EDIT ��/%7����*S�YSTEM*upV�9.40107 �cr7/23/2021 A���Pw��PRGAD�J_p  h �$X[�p $Y�xZ�xW�xқt�ZқtSPEED_��p�p$NEXT�_CYCLE�p����q�FG�p� ��pALGO�_V �pNYQ�_FREQ�WI_N_TYP�q)��SIZ1�O�LA!P�r!�[��M+�����qCREATED��r�IFY�r@!N�AM�p%h�_G>J�STATU��J��DEBUG�rMA�ILTI����E�VEU��LASTx�����tELEM�� � $EN�AB�rN�EASI�򁼁AXIS�p�$P߄�����qR�OT_RA" �rM�AX ��qE��L�C�AB
���C D�_LVՁ`�BAS ��`�1�{���_� ��g$x���RM� 9RB�;�DIS�����X_SPo�΁�� ��u�P� | �	� 2 6\�AN�� �;������Ӓ�� |�0�PAYLO��<3�V�_DOU�qS�x��p�tPREF�� ( $GR�ID�E
���R����Y�  �pO�TOƀ�q  ��p��!�p��k�O�XY� � ;$L��_PO|��נVa�SRV��)����DIRECTS_1� �2(�3(�U4(�5(�6(�7(��8��qF��A�>� $VALu�GROUP�����}F�� !��@!�������GRAN泲���R��</���TOTA��,F��PW�I=!%�REGEN#�8��������/���ڶnT0zЉ���#�_S����8�(�V[�'���4���GGRE��w���H���D�����V_H��D�AY3�V��S_Y��Œ;�SUMMA�R��2 $C�ONFIG_SEpȃ���ʅ_RUN��m�C�С�$CMPuR��P�DEV��4�_�I�ZP�*������ENHANCUE�	�
����1���INT��qM�)b�q�2K����O�VRo�PGu�IX8��;���OVCT���|��v�
 4 �����a˟��PSLG|"�� \ � ;��?�1���SƁϕc�U�����Ä��4�U�q]�Tp�� (`�-��rJ�<�O� CK�IL_�MJ���VN�+��TIQn{�N5���C�SULȀD�V(�C6��P_�຀@�MW�V�1V�V1d�2s�2�d�3s�3d�4s�4 d��'�	�������p�	�IN	VIB1qp1� 2!pq/,U3 3,4 4, �p?��;��A���N��������PL��TORr3�	��[��SAV��d��MC_FOLD~ 	$SL�(����M,�I���L� �pL�b��K�EEP_HNAD�D	!Ke�UCCOMc�k��
�lOP���p�l��lREM�@k��΢���U���ekHPW� �KSBM��ŠCOLLAB|�Ӱn��Zn�+�IT�O���$NOL�FCA9LX� �DON�r����� ,��F�L���$SYNTy,M�C=�����UP_DLY�qs"DELA� �����Y(�AD��$T�ABTP_R�#���QSKIPj%3 ����OR� �E�� P_��� �)� ��p7��%9��%9A� $:N�$:[�$:h�$:u��$:��$:9�q�RA�� X������MB�NFLIC�]��0"�U!�o���N�O_H� �\�< _�SWITCHk�R�A_PARAMG�� ��p��U���WJ��:Cӣ�N/GRLT� OO�U������X�<A��T_J�a1F�rAPS�WE�IGH]�J4CH��aDOR��aD��O!O��)�2�_FJװ����sA�AV��C�HOB�.�.�l�J2�0�q�$�EX��T$�'QIT��'Q�pG'Q-�GΨ�RDC�m" G� ��<��
R]���
H���RGEAp��4��U�FLG`�g��H��ER	�SsPC6R�rUM_'P>��2TH2No��@~Q 1 @�ED����  �D �وIi�2_P�25cS�ᰁ+�_L10_CI��pe� �pk�� ��UՖD��zaxT�p�Q(�;a��c���޲+�i���e��`� P`DESIG\Rb$�VL1:i1Gf��c�g10�_DS���D��w�POS11�q l�pr��x1C/#AT�Br��U
WusIND�Ѐ}�mqCp�mq`B	�H7OME�r 	aBq2GrM_q��(��!@s3Gr��@� ��$�`!@s4GrG�Y�k�}�����6�5Grď֏�������6GrA�S�e�Pw�����6�7Gr��@П�������8Gr;�M�_�q��������S �q     �@sM��P�!�K@��! T`M��M��IO��m�I��2�OK _OPy��� »Q�6�POWE"� 7�x EQ�1E� � #s%Ȳ$D;SBo�GNA�b� C�P2�BS23�2S�$ �iP���xc�ICE<@%�P1E`2� @IT��P��OPB7 1�FLO�W�TRa@2��U�$�CUN��`�AUX�T��2Ѷ�ERFAiC3İUU��;CH��% t<�_9�EЎA$FR?EEFROMЦ��A�PX q�UPD�"YbA�PT.�pEE�X0����!�FA8%b�/��RV�aG� &  ��E�" 1�AL�  ��+�jc'��D�  ?2& �S\PcP?(
  �$7P�%��R�2� ��T�`A9XU���DSP���@@�W���:`$��RNPн%�@����K��_McIR�����MT��AP���P"�qD��QSYz������QP=G7�BRKH����� AXI�   ^��i���1 ����OBSOC���N��DUMMY16�1o$SV�DE���I�FSPD_OV%R79� D���ӓOR��֠N"`��F�_����@OV��SFN�RUN��"F0�̊���UF"@G�TO�d�LCH�"�%REGCOV��9@�@W�`@&�ӂH��:`_0��  @�RTINsVE��8AOFS��9CK�KbFWD���`���1B��TR�a�B �FD� ��14= B1pBL� �6� A1L�V��Kb�����#��@+<�AM�:��0��j��_M`@ ~�@h���T$X`�x ��T$HBK ���F��A�����PPA�
��	�������DVC_DB�3@pA�A"D��X1`�X3`@��S�@�`�0��U���h�CABPP
R�S  #��c�B�@���G�UBCPU�"��S �P�`R��11)A�RŲ�!$HW_�CGpl�11� F&A1�Ԡ@8p�$UNI�Tr�l e ATT�RIr@y"��CYC�5B�CA��FLTR_2_FI�������2bP��CH�K_��SCT��F�_e'F_o,�"�*FqS�Jj"CHA�Q��'91Is�82RSD�����1���_T`g�`� i�EM��NPMf�T&2 8px&2- �6DIAGpE?RAILACNTB�Mw�LO@�Q��7&��PS��� � ���PRBSZ`�`�BC4&�	��FUuN5s��RIN�P`Zaߠ�07Dh�RAH@���`� `C�@�`C��Q�CBLCUR�uH�DA�K�!�H�HD�Ap�aA�H�C�ELD@������C��jA�1��CTIBUu�8p$CE_RIA�QVJ�AF P��>S,�`DUT2�0C��}�;OI0DF_aLC�H���k�LML}F�aHRDYO���RG�@HZ0��ߠ|�@�UMULSE�Pt�'3iB$J���J����FAN_�ALM�dbWRNeHARD��ƽ�	P��k@2aN�r�J�Y_}�AUJ R+4~�TO_SBR���~b�Іje 6?A�cM/PINF��{!�d��A�cREG�NV���ɣZ�D��NF9LW%6r$M�@� ���f� �0 h'uC�M4NF�!�ON 	 e!e#�(b*r3F�3G �	 ���q)5�;$�$Y�r���Zu�_��p*$ �/�EGE�����F�qAR��i���2�3��u�@<�AXE��R�OB��RED��W�R��c�_���SY�`��q� ?�SI�WR1I���vE STհ��(� d���Eg!��t8��^a��B���񐆹9�3� OTO�a���ARY��ǂ�1�����FIE����$LINK�QGT5H��T_�������30���XY�Z���!*�OFF������ˀB��,Bl������m�FI� ��C@Iû�,B��_J$�F������S`����3-!$ 1�w0���R��C��,�DU���3�P�3TUR`XS.�Ձ�b1XX�� ݗFL�d�`��pL�0���34��^�� 1)�K��	M�5�5%B'��ORQ�6��fC����0B�O;�D�,��p����a�OVE��rM�����s2��s2� �r1���0���0�g /�AN=!�2�DQ�q� ��q�}R�*��6���0�s��V���ER��jA�	�2E��.�C��A���0��XE�2Ӈ�A��AAX��F��A� N!�SŴ1_��Q_Ɇ� ^ʬ�^ʴ�^��0^ʙ�^ʷ�^�1&�^ƒP[� �PkɒP{ɒP�ɒP�� �P�ɒP�ɒP�ɒP������ɪ �R>�DEBU=#$8ADc�2����
�AB�7����9V� <" 
��i �q��-!��%��׆��� ���״����1�י������JT��DR�m�LA�B��ݥ9 FGR�O� ݒ=l� B_ �1�u���}��`����pޥ��qa��AND������qa�  �Eq��1��A@�� ��NT$`��c�VEL �1��m��1u���QP��Fm�NA[w�(�CN1�� ��3줙�  ��SERVEc�p+� $@@d@��!���PO
�� _�0T� !�򗱬p�,  $T�RQ�b
(� -�DR2,+"P�0_ . l"@!�&'ERR��"I� q𜍴~TOQ����L��p]�e���0G��%l�����RE�@ / ,��/I �-��RA� 2�. d�&��_n! 0�p$&�0�2tPM��OC�A8 �1  pCO�UNT�� ��FZ�N_CFG2 4B �f�"T�:#��Ӝ� � `�s/3 ���M:0�R��qC@��/�:0�FA1P��?V�X������r���� �P�:b��HELpe�4 5��B_wBAS�cRSR�f� @�S�!QY 1T�Y 2|*3|*4|*U5|*6|*7|*8��L!RO�����NL�q �AB���0Z �ACK��INT�_uUS`�Pta9_cPU�>b%ROU��PH@�h9#�u`w�9��TPFWD_KA1R��ar RE���PqP��A]@QUE�i@&��	�f�>`QaI`���9#�j3r��f�SCEME��6��PA�7STY4SO�0�DI'1�`���18�rQ�_TM�cMANR�QXF�END��$KEYSWIT�CHj31:A�4HE�	�BEATM�3PE�pLE��1��H�U~3F�42S?DD_O_HOMBPO:a60EF��PRr��(*�v�uC�@O�Qo ��OV_Mϒ��E�q�OCM���7��p8%HK�q5 DH��g�Uj�2M�px�4R��FORC�cgWAR��NYOM�p 6 @�Ԣ�v`U|�P�p1�V'p�TE3�V4��OR#O�0�L�R7��hUNLiOE0hdEDVa�  �S�@d8� <pAQ9�l1M�SUPG�UaCALC_PLANccM1��AYS1�1:b>�9 � X`��P �q;a�թ�w��2��j�M$P�㣒�fXyt$��rSC�M�p m�q ���aq��0�t5YzZzEU�Q�b�� T!�Hr�pPv	�NPX_ASf:; 0g ADD���$SIZ%a$�VA��MULTKIP�"ns�PA�Q; � $T9�op�B���rS��j!C<~ �vFRIF�2aS�0�YT�pNF[DODBUX�B��u&��!���CMtA�Е� ��������+Z ��< � �p�T�Eg�����$SGL��T��X�&{����<����STMTe�Ѓ�PSEG�2��BW<���SHOW؅�17BAN�`TPO����gᣥ��������V��_G�= ��$�PC���O�FBZ�QP\�SP�0A&0�^�� VDG��>�� �cA00 �����P���P���P��T�P��5��6��7��8��9��A��b`��@�P��w᧖��F����h���1��v�h�יU1�1�1��1�U1�1%�12�1?�U1L�1Y�1f�2��U2��2��2ʙ2יU2�2�2��2�U2�2%�22�2?�U2L�2Y�2f�3��U3��3��3ʙ3י�3�3�����3��3%�32�3߹3�L�3Y�3f�4��4���4��4ʙ4י4��4�4��4�4��4%�42�4߹4�L�4Y�4f�5��5���5��5ʙ5י5��5�5��5�5��5%�52�5߹5�L�5Y�5f�6��6���6��6ʙ6י6���6�6��6�6�(�6%�62�6߹6�L�6Y�6f�7��7���7��7ʙ7י7���7�7��7�7�(�7%�72�7߹7JL�7Y�7f�[V�`�_UPD��? <�c 
ZB�����@ x $T�OR�1T�  �cO�P �, ZQ_7RAE^��� J��SsiC�A��_U�p���YSLOA"A � �u$�v���w�@���@��bVA�LUv10�6�F��ID_L[C:H�I5I�R$FILcE_X3eu4$�C�7 �SAV��B �hM �E_BLC�K�3�ȁ�D_CPU��p��p5h�z��@S2R C? � PW��� �	�!LAށSRp�#.!'$RUN�`G@%$D!'$�@G%e!$e!'%HR03$� '$v7aT2Pa_LI�R�D  � G_�O�2�0P_ED�I�R�"SPD�#�E�"i0ȁ�p�Q��DCS9@G)F� � 
$JPC�71��� S:C;C�9$MDL7�$5P>9TC�`@7U�F�@?8S� ?8CO�Bu �@�"|�L�G��P;;� 9�:;�qTABUI�_�!L�HGb�% sFB3G$�3�A�sR�LLB_AVAI�B���3�!��wI $� SEL� sNẼ�@RG_D �N��Ta���4S=C�PJ �1/A�B�PT�R?�w@_M]`L�K \M f/Q�L_��FMj��PG�i�U9R�6��PS�_�P\� �p�EE�7B�TBC2�eL� ���``�`b$�!FT�P'T�`TDCg�� BPLp�sLNU;WTH��qhT�gtWR�2$�pERVE.S�T;S�Tw��R_ACkP MX -$�Q�`.S �T;S�PU@�`IC�`7LOW�GF1�QR�2g�`��p�S�ERTIA�d^0iP��PEkDEUe�LA7CEMzCC#c��V�BrpTf�edg�aT�CV�l�adgTRQ �l�e�j|�Scu��edcBu�J7_ 4J!���Se@qde�Q2��0���1�PRcuPJKlvVK<�~qcQ~qw�bspJ0��q�sJJ�s;JJ�sAAL�s�p �s�p�v���r5sS�`N1�l�p�k�`5dXAa_́� PCF�B�N `M GROUP ��bh�NPC0s~D�REQUIR�R�� EBU�C�Q�6g0 2Mz��Pd�VQSGUO�@�)/APPR0C7@� �
$� N��CLO�� ǉS^U܉Se>@BuC�@A�"P �$P�M]P�`�`sR�_M	Ga!�C���+��0��@,�BRK*�NO�LD*�SHORTCMO�!m�Z��JWA�SP�tp`�sp`�sp`@�sp`�sp`�A��7���8sQIR_�RTQ�� m��R.Qx�cQ�PATH��*� �*��X&���P�NT|@A�"p���6 �IN�RUC4`aZ��C�`UM��Y
`�)p��>�Q��cP����p��PAYLO�Ah�J2L& R_	Am@�L ������+�R_F2LS3HR�T/�LO���p0���>���ACRL0 z�p�y�ޤsRH5b�$H+���FLE�X��#�JVR P��_._�_�_Q}J�US :�_ �Vd`0�G��_tQd`�_�_lF1G��ũ�o@0oBoTofoxo��E�o �o�o�o�o�o�o  ����wz3lt����3�EWF�^zT!��X ���ju��uu~�W� ����p�u�u�u�u0����UM��(�T �P5�G�Y��' AT��l�pELP0�_B��s�J�Sz�;JEW�CTR7B`�NA��d�HAND_VB����TEUO@`+�`T�SW8F�A�V� $$M��e G��AV�Qs�De�oA@A��@�	$�A5�G�AU�Ad�� 6�T�G�DU�Dd�PD�G/ -STI�5V�5Ng�DYF ��+� x����P&�G�&�A�@�lw�o�Q�k�P�������ʕӕܕ��D9X�TW 7 Ć� ��3%�?!A'SYMT�(�m�T��V*�o�A�t�_SH �~������$����Ưد�J񬢐�#3�9"���_VI���`8�q0V_UNIrS�4��.�Jmu�2� �2A��4X��4�6a�p@t�������&E_������RE��CH( X ̱���[TOc�PP�VsS(vD�US�RU�P���� �z@�D�A}@_5�U���P�EyAa��RPROoG_NA��$��$LAST���C�ANs�ISz@XYZ_SPu�DW]R@�Ͱ,VSV@�E1QENc��DCUR�H#���oHR_T��YDtQ9S�d��O�T� 
Z�tQ?�Z) ��I�!A�D�� �Q���#�S���� �3��vP [ � ME�O��R#B�!T�PPT0F@1�a-�1�̰� h1a�%iT0� $�DUMMY1��o$PS_��RF���!�$lfװFL�A*�YP�bc?$GLB_TI �Up�e`ձ��LIF(!�\����g`OW��P��eVOL#qLb �a_2��[d2[`����b�P�cZ`T�C��$BAUD,v��cST��B�2g`�ARITY0sD_[WAItAIyCJ�2�OU6�ZqyyT�LANS�`�{S�SyZc��BUF_�r��fиx�PyyCHK]_�@CES��� +JO`E�aA�x�bUBYT���� �r�.�.� ��aA���M�������Q] �Xʰ����ST����SBR@M21�_@��T$SV_cER�b����CL�`ʐ�A1�O�BpPGL�h0EW(!^ 4 �$a$Uq$�q$W�9�A��@R����ӃU�م_ "��D$�GI��}$ف �^��(!` qL�.��"}$F�"=E6�NEAR��B'$F}��TQL����J�@R� a�mP$JOINT�a�)�&ՁMSET.(!b  +�Ec�2ъ^�ST��H�_�(!c��  ��U�?����LOCK_F�O@� �PBGLV���GL'�TE�@X9M���EMP����qK��b�$U��؂a�2_���q�`�<� �q�^��CE�/�?��� $KAR�b�M�STPDRA8܀����VECX���֪�IUq�av�HE��TOOL���Vv��REǠIS3�2�6��ACH̐m Mb^QONe[d3����IdB�`@$RAIL_BOXEa���ROB�@D�?����HOWWAR�0Aa�i`-�ROLM tb��$�*���T��`��n��O_FU�!��HTML58QS��@ e�"Հ�(!d��#��@�(!e��Ļ���І}p(!f 	t��m�^a��t��VB�PO��AIPE�N���O����q�|�AORDED��m �z�XT`��A)� ��P�O�P �g D �`OB �����ǯ�Uc�`���� ��SYS��AD�R��pP`U@^  �h ,"��f$A���E��EтVW�VA�Qi � 1�@ق�UPR�B��$EDI�Ad�V/SHWRU�z���cIS�Uq�pND�Px7���G�HEAD�!h @���!i�KEUq�O`CP)P��JMP���L�U�TRA[CE�Tj����IL�S��C��NEx���TICK�!M4�_N��H=Nr�k @���HWC��P�FF��`S3TYeB+�LO�a9�P' ��[�C�l3�
�@��F%$A��D=��S�!$�1�p a�e��q�ePv �FSQU̩�#LO�b_1TE�RC`!oPS?�m 5���R�m@3����ܡ�O`	c IZ�d�A�eha�qtb�}�hA}pP~r��_D)O�B�X�pSSQ�S'AXI�q��v�bS��U�@TL���RE3Q_ܠ��ET���`@�CY%�P��Z&��Af�\!\d9x�P �MBSR$$nl-�w �����c
��uV
Qh(�A ���dC`�A�� 	�Y��D��pH�E"�	CC�C���/�/�/	4ISC��` o h��D1Smడ[`SP�@�AT� 
R��L���XbADDR�s$�Hp� IF�Ch�_2CH���pO����- ��TUk�Ir �p�CUCp�V
��I�Rq�4���c
��
K�
��^ ���P'r \z�D����|,K� P�"CN��*�CƮ��!�TXSCREE��s�Pp@��INA˃<�4�Dp������`t T� ���b����O Y6������U4h�RR��������R1�T  �UE��u �j �qz`9Ś��RSML���U����V�1tPS_ ��6\��1�9G\���qC��2@4 2���0Ov�R��&F�A�MTN_FL*��`Q��W� ��BBL�_/�WB`�Pw �ԫ��BO ��BLE�"�Cg�R"�DRIG�HtRD��!CKGRB`�ET���G�AWIDTHs���RxB��a�r�UI��sEYհRx d��ʰ�����`y�BACCK��tb>U���PsFO��QWLAB��?(�PI��$�URm�~P�P�PH�y1 y 8 $�PT_��,"�R�PRUp�s5�da���Q)O%!t�zV�ȇ�p�U�@�SR ���LUqM�S�� ERVJ��SP��T{ � " GE�Rh� ��&��LPAeE��)^g�lh�lh�ki5ik6ik7ikpP`@�Z�x����$u1���p�Q zQU{SRل| <z�b�PU2�a#2�FOO .2�PRI*m9�[��@pTRIPK�m��UNDO��}�)���Yp��y���q�h����p ~�R\p�qG ��T����-!�rOS2��vR ��2�s�CA��H���ro���Pi�UIaCA����3Ibn�s�OFFA�D@���Ob�r���L�t��GU��Ps���������+QSUBo� }��E_EXE���VeуsWO� e�#��w��WAl��p΁fP
 V_CDB���pT�p�O�V░���3OR�/�5�RAU@6�T�K���__����s |j �OWNj�>34$SRC�0`����DA���_MPFqI����ESP�� T�$0��c��g�Y�8q�z�E!� `%�ۂr34J���COP��$���p_���/�+�6���CT�Cہ��ہ�D �DCS���P4�C3OMp�@�;�@�Oo�=���K��^�/�VT�q'�
��Y٤Z��2����@p�w#SB����2�\0˰_��M��%!]�gDIC#��AY�3.G�PEE�@T�QS�#VR1���eQL�� a��P�D ��f�z���f�> ���6�FP��A�t�b# �L2SHADOW��#ʱ?_UNSCAd�׳�OWD�˰DGDE>#LEGAC)�q'��VC\ C��� v����だ�m�RF07���7d`C�2`7�DRIVo���ϠC�A]�(�` ��~�MY_UBY�d ?Ĳ��s��1��$0飈����_ఆ���L���BM�A$�DEY	�EXp@C�/��MU��X��,��0U1S��.�;p_R"1��0p#�2�GPAgCIN*���RG�� c�y�:�y��sy�C/�CRE�R"!�q��Üy�D@� L !�GB�P�"�г��R�p�D@�&P�Px1Q��	l.���RE��SWqГ_Ar��+�{�ODq�AA/�3�hEZ�9U���� P�+HK���PJ��p_/�Q0{�EAN���ۀ2�2��P�MRC�VCA� �:`ORG��Q�dR	��L�����REFoG����� !�+`	�p����� ���<���q�_����r��� S�`C��Ú�8G�@D� ��0�!`��#q�š�OU��<��?� ��Վ�2�J@0� 1�*p�����0 UL6�@��CO�0)�3�� NT�[���Z�Qf�af% L�飏��Q��a��VIAچ� ��@HD7 6P$J�O�`oB�$Z�_UPo��2Z_LOW��$�QiBn��1$EP�s�y@�� 1!f m� |1¦4� 5��PA�A �CACH&�LO�w��ВQB���Cn�I#F^��Tm����'$HO2�32{��Uÿ2O�@���Ro0��=a��ƐVP��X@�A"_SIZ&�K$Z�$�F(�G'���CMP�k*FAIo�G��AD�)/�MRE���"P'GP�0е��9�ASYNBUFǧRTD�%�$P!�COLE_2D_4�"5W�sw�~�UӍyQO��%ECCU�؇VEM��v]2�VIRC�!5�#�2�!�_>�*&�pWp��AG:	9R�XYZ@�3�W���8��4+Qz0T"��IM�16�2|P�GRABB�q\��;�LERD�C �;�F_D��F�f5!0MH�PE�R�[��� ��KQLAS��@��[_GEb�� �H൑~23�ET@����"���b��I�D��ҙ6m�BG_LEVnQ{�PK|Л6\q���GI�@N\P4� n��A��!g�dr��S� �NRT�V	Lʁc�Ų��#a�4�c"!D�qDE��� �Xа�X�����1��d��pzZ���dT�c���D4qȲ��2pT��U&�� $�ITPr9p[Q�ŜՓV�VSF$�d��  fp/�f�URl&ҿ�SMZu�dr���ADJ`C�� Z�DVf� D�XA�L� � 4 PER�IKB$MSG_Q3$Q!o%[���p'��dr:g�qQ�^ �XVR\t��B�pT_\��R��ZABC"����Sr����
W��aACTV�S' � � �$|u�0�cCTIV�Q!IOu¥s&fD�IT�x�DVϐ#
x�P���!��M�pPS���� �#༒!���q!LST`D�!�  �_ST�c��aq�CHx�� L-�@��u�Ɛp*���P GNA#��C�!q�_FUN��� uqIPu���HR�$L����XZMPCF"���`bƀ�rX�ف��LN�K��
Ł�0#�� $ !��ބ�CMCMk�C8�C�"����P{q '$J8�2�D6!>� O�H���T���2������M���UX�1݅UXE1Ѡ��1C���Y���ੑ����˗7�FTFpG>�������Z���� �k�� ���YD'@ W� 8n�R� Uӱ$HEIGHd�F:h?(! 'v���|���� � Gd��qp$B% � E���SHIF��hRVBn�F�`�HpC�  3�(�8H`O�ѡ�Cd��+%D	�"�CE�p�V���SPHER>s� � ,! M��c�u��$POW�ERFL �R|�2���|�p�RG�`����������A�  ��?h`��`d��NSb� ���?�  Bz|�} l�  <@�|��%���˃�p���ŵ�� 2ӷ^�� 	H��l&����>����A |��t$���*��/�� **�:��`�ϥ��͘����������ɘ� �|�����5������ �%ߟ�I�[߉�ߑ� ����������w�!� 3�a�W�i������� ����O����9�/�A� ��e�w�������'�� ���=O} s������� k'UK]�� ����C/��-/ #/5/�/Y/k/�/�/�/ ?�/�/?�/?�?1? C?q?g?y?�?�?�?�? �?�?_O	OOIO?OQO�� 	 �O�O�O _�E��3_���O`_�O��_�_÷PREF SӺ``
��IORITY `�|���`����pSP0L`z����WUT�Vq�Έ�ODU~������_?�OG��Gpx��R��,fHIBq�Oy�|kTOENT� 1��yP(!�AF_b�`�o�g�!tcp�o}�!ud�o)~!�icm�0bXuY̳�k �|��)� ����������u���� ��N�5�r�Y����� ��̏�����*/c̳�ӹ���E�W�|�>W�^�F��/��H4���|��,�7�A���,  ��P@����%�|�'����Z��h�z�����|���ENHANCE� 	#�7�A9�dx�����  �,f��T
�_�S����P�ORTe�rb����U��_CART�REP�Pr|brSK�STAg�kSLGmS�`�k������Unothing������Ϳ�>�P�b�To��TEM�P ?isϨE�/�_a_seibanm_��i_����� 0��T�?�x�cߜ߇� ���߽�������>� )�N�t�_����� ��������:�%�^� I���m�����������  ��$H3lW i������ �D/hS�w���uϪ�VER�SI�P=g  �disable���SAVE �?j	2670/H705��k/�!�m//*�/ 	��(%b�O�+�/�Se@?6?H?Z?l?z:%<Т/�?4�*'_j` 1�kX �0ubuE��?OqG�PURGEb��Bp`�ncqWF<@�a�TӒ*fW�`]Da�a�WRUP_DE?LAY z�f��B_HOT %�?e'b��OnER_NORMAL�HGb�O<%_�GSEMI_*_|i_�QQSKIP�3	.��3x��_��_ �_�_�]?eo+goKo ]ooo5o�o�o�o�o�o �o�o�o5GY i�}����� ��1�C�U��y�g� ��������я�����-�?�7%�$RACFG �[ќ�3��]�_PARA�M�Q3y��S @�И@`�G�42C�۠��2��C�bFB�B]�BTIF����J]�CVTMO�U�����]�D�CR�3�Y ���Q>�g�@���B�@�jx��S��{�����5�?C����0�_��~\� ;e�m����KZ;�=g;�4�<<���pf@����� � 5�G�Y�k�}��������ſ׿���xURDI�O_TYPE  ��V�5��EDPR�OT_a�&Y>��4BHbCEސ�SǆQ2c� ��B�ꐪϸ���� �����&�ݹ�W�V_ ~�o����߱����� ����A�O�m�r��� 9����������� ���=�_�d����� ������������' I�Nm���� �����#EJ i+k���� ��//4/F//g/ /�/y/�/�/�/�/�/ 	?+/0?O/?c?Q?�? u?�?�?�?�?�??;?�,O��S�INT 2��I���l�G;�� jO|K��鯤O�f�0 �O�K�?�O�? ___N_<_r_X_�_ �_�_�_�_�_�_�_&o oJo8ono�ofo�o�o �o�o�o�o�o"F 4j|b����������B�O�E�FPOS1 1~"�  xO ��o×O����ݏ鈃� ��Ϗ0��T��x�� ��7���ҟm������ ��>�P����7����� ��W��{�����:� կ^����������S� e��� ��$Ͽ�H�� l��iϢ�=���a��� ��� ߻����h�S� ��'߰�K���o���
� ��.���R���v��#� 5�o���������� <���9�r����1��� U�����������8# \����?�� u��"�FX� ?���_�� /�	/B/�f//�/ %/�/�/[/m/�/?�/ ,?�/P?�/t??q?�? E?�?i?�?�?O(O�? �?OpO[O�O/O�OSO �OwO�O_�O6_�OZ_ �O~_�_+_=_w_�_�_ �_�_ o�_Do�_Aozo<cf�2 1r�o .oho�o�o
o.�o R�oO�#�G� k�����N�9� r����1���U����� �����8�ӏ\���	� �U�����ڟu����� "����X��|���� ;�į_�q������	� B�ݯf����%����� [���ϣ�,�ǿٿ �%φ�qϪ�E���i� �ύ���(���L���p� ߔ�/�A�Sߍ����� ��6���Z���W�� +��O���s����� ����V�A�z����9� ��]���������@ ��d��#]�� �}�*�'` ���C�gy ��&//J/�n/	/ �/-/�/�/c/�/�/? �/4?�/�/�/-?�?y? �?M?�?q?�?�?�?0O �?TO�?xOO�O�o�d3 1�oIO[O�O _�O7_=O[_�O__ |_�_P_�_t_�_�_!o �_�_�_o{ofo�o:o �o^o�o�o�o�oA �oe �$6H� ����+��O�� L��� ���D�͏h�� �������K�6�o�
� ��.���R���퟈�� ��5�ПY�����R� ����ׯr�������� �U��y����8��� \�n�������?�ڿ c�����"τϽ�X��� |�ߠ�)�������"� ��nߧ�B���f��ߊ� ��%���I���m��� ,�>�P��������� 3���W���T���(��� L���p����������� S>w�6�Z ����=�a � Z���z /�'/�$/]/��/�/�/@/�/�O�D4 1�Ov/�/�/@?+? d?j/�?#?�?G?�?�? }?O�?*O�?NO�?�? OGO�O�O�OgO�O�O _�O_J_�On_	_�_ -_�_Q_c_u_�_o�_ 4o�_Xo�_|ooyo�o Mo�oqo�o�o�o�o �oxc�7�[ ����>��b� ���!�3�E����ˏ ���(�ÏL��I��� ���A�ʟe���� ���H�3�l����+� ��O���ꯅ����2� ͯV����O����� Կo�����Ϸ��R� �v�Ϛ�5Ͼ�Y�k� }Ϸ���<���`��� ��߁ߺ�U���y�� ��&���������k� ��?���c������"� ��F���j����)�;� M���������0�� T��Q�%�I��m��/�$5 1 �/���mX�� �P�t�/�3/ �W/�{//(/:/t/ �/�/�/�/?�/A?�/ >?w??�?6?�?Z?�? ~?�?�?�?=O(OaO�? �O O�ODO�O�OzO_ �O'_�OK_�O�O
_D_ �_�_�_d_�_�_o�_ oGo�_koo�o*o�o No`oro�o�o1�o U�oyv�J� n������� u�`���4���X��|� ޏ���;�֏_����� �0�B�|�ݟȟ��� %���I��F����� >�ǯb�믆������ E�0�i����(���L� ��翂�Ϧ�/�ʿS� � ��LϭϘ���l� �ϐ�ߴ��O���s� ߗ�2߻�V�h�zߴ� � �9���]��߁�� ~��R���v����#�<	6 1&�� �������������}� ��<��`��� �CUg�� &�J�n	k� ?�c��/�� �	/j/U/�/)/�/M/ �/q/�/?�/0?�/T? �/x??%?7?q?�?�? �?�?O�?>O�?;OtO O�O3O�OWO�O{O�O �O�O:_%_^_�O�__ �_A_�_�_w_ o�_$o �_Ho�_�_oAo�o�o �oao�o�o�oD �oh�'�K] o�
��.��R�� v��s���G�Џk�� �����ŏ׏�r�]� ��1���U�ޟy�۟� ��8�ӟ\������-� ?�y�گů����"��� F��C�|����;�Ŀ _�迃������B�-� f�ϊ�%Ϯ�Iϫ��� �ߣ�,���P�6�H�7 1S����I� �߲�������3��� 0�i���(��L��� p�����/��S��� w����6�����l��� ����=������6 ���V�z�  9�]��� @Rd���#/� G/�k//h/�/</�/ `/�/�/?�/�/�/? g?R?�?&?�?J?�?n? �?	O�?-O�?QO�?uO O"O4OnO�O�O�O�O _�O;_�O8_q__�_ 0_�_T_�_x_�_�_�_ 7o"o[o�_oo�o>o �o�oto�o�o!�oE �o�o>���^ �����A��e�  ���$���H�Z�l��� ��+�ƏO��s�� p���D�͟h�񟌟� ��ԟ�o�Z���.� ��R�ۯv�د���5��ЯY���}�c�u�8 1��*�<�v���߿ ��<�׿`���]ϖ� 1Ϻ�U���y�ߝϯ� ����\�G߀�ߤ�?� ��c����ߙ�"��F� ��j���)�c���� ������0���-�f� ���%���I���m�� ����,P��t �3��i�� �:���3� �S�w /��6/ �Z/�~//�/=/O/ a/�/�/�/ ?�/D?�/ h??e?�?9?�?]?�? �?
O�?�?�?OdOOO �O#O�OGO�OkO�O_ �O*_�ON_�Or___ 1_k_�_�_�_�_o�_ 8o�_5ono	o�o-o�o Qo�ouo�o�o�o4 X�o|�;�� q����B��� �;�������[��� ����>�ُb������!�������MASKW 1 ��������ΗXNO  �ݟ���MOTE � ���S�_CFG !Z���N������PL_RANG�V�N������OWE/R "��Ϡ���SM_DRYPRoG %���%W���եTART �#Ǯ�UME_P�RO���q���_E�XEC_ENB � ����GSPD�J�������TD�B����RMп��I�A_OPTION��������N�GVERS���`�řI_AIoRPUR�� R��+���ÛMT_֐T� X���ΐOBOT_ISOLC�A�������u�����/NAME8��H�Ě�OB_CATEG�ϣ,��S�[�.��ORD_NUM �?Ǩ��H705  N��ߨߺ�ΐPC_T�IMEOUT�� �xΐS232s�1�$��� L�TEACH PENDAN��o�������V�T�M�aintenance ConsN��&�M�"B�P�No Use6�r�8�������̒��N�PO$��Ҋ�"�^��CH_LM�Q�朕	a�,�!U�D1:��.�RՐVgAILw��粥�*�SR  t�� ���5�R_INoTVAL����� ���V_DAT�A_GRP 2'|���� D��P�������	�� ����B0 RTf����� �/�/>/,/b/P/ �/t/�/�/�/�/�/? �/(??L?:?p?^?�? �?�?�?�?�?�?O O "O$O6OlOZO�O~O�O �O�O�O�O_�O2_ _ V_D_z_h_�_�_�_�_ �_�_�_o
o@o.oPo�vodo�o��$SA�F_DO_PUL�SW�[�S���i�SC�AN�������S�Cà( ��!���S�S�
���Ķ�(q�q�qN� �L ^p���5��`� ��$��+�E�r2M�qX�dM��h�J�	t/� @���������ʋ|��� �r ք��_ @N�T ��'�9�K�~X�T D��X� ��������ɟ۟��� �#�5�G�Y�k�}������䅎�p����Ǧ  "�;�oR� ���p�"�
�u���Di���q$q�  � ���uq�� \�������ҿ���� �,�>�P�b�tφϘ� �ϼ���������(� :�L�^�p߂ߔߦ߸� ������ ��$�6�H�Z����珈���� ��������g�;�D� V�h�z���������������(�Ӣ0�r�i� y���$�7I[m ������� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/?r�+?=?O? a?s?�?�?�?�?�?8� �?OO'O9OKO]OoO �O��$�r�O�O�O �O	__-_?_Q_c_u_ �_�Y�_�_�_�_�_o o&o8oJo\ono�o�o �o�o�o�o�o�o"�4FXj|�c�� ��g������� 0�B�T�f�x������� ��ҏ������\:�Ҧ��y�3��	�	12345�678��h!B�!�� 
\��p0����Ο �����(�:�@�� c�u���������ϯ� ���)�;�M�_�q� ����R���ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����ϖ����� 1�C�U�g�yߋߝ߯� ��������	��-��� Q�c�u������� ������)�;�M�_� q���B���������� %7I[m �������� !3EWi{�� �����//// �S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?D/�?�?�?�? �?OO'O9OKO]OoO��O�O�O�O�O�O*� ���O	_�E�?5_G_Y_��yCz  A���z   ��x2��r }��)�
�W�  	�*�2�O�_�_H oo"l�#\��_ hozo�o�o�o�o�o�o �o
.@Rdv ����Mo��� �*�<�N�`�r����� ����̏ޏ����&�8�J��X #P$P�Q�R�<u� k��Q  ������S��P���Q�Qt  ��PÙ۟�P(� `,b����]�PFl��$SCR_GR�P 1*!+�!4� � }�,a �U�	 v��~������d����%���ɯ���h]���P�D1� D�7n��3��Fl
�CRX-10iA�/L 23456�7890�Pd� 4r��Pd�L ��,a�
1o��������[ ¶~�+fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@�R�d�~t���H�~�Ă�m��ϴ������ϼ��,a��1��ϨU�[�G�imXhuP,�[}��P0���B�  BƠߞҷ�r��A�P��  @1`��՚�@����� ?	���H����ښ�F@ F�`A� I�@�m�X��|���� ��������������`:�%�7�I�[�B�i� ��������������� -Q<u`��@En�ٯ���W�P�"+f@_�5��1`4b���x����ͣ�O�,dA����$���Fa�,a �#!"/4/E-!�Z(f/x/G/ (�P�!(� �/�/�/��/�/?#9b�����S7س�M�ECLV�L  ,a���ݲ�Q@f1L_D?EFAULTn4b1_�1`�3?HOTSTR�=���2MIPOWER�Fm0pU�5�4W7FDO�6 �5L��ERVENT 1�+u1u1�3 L!�DUM_EIP�#?5H�j!AF�_INE�0SO,d!'FT)O�NIO�O9!���O ��O�O�!RPC_MAIN�O�H��O>_S'VIS_�I�-_�_?!OPCUf�_�Wy_�_!TMP�PPU�_<Id�_�"o!
PMON_�PROXY#o?Fe ono�R<o8Mf]o�o�!RDM_SR�V�o<Ig�o!�R��"=Hh�oR!%
PM�o9LiA��!RLSYNC̟�y8��!gROS(O��4��6�!
CE�PMT'COM7�?Fk%���{!	K�CONS���>Glq�Ώ!K�WOASRC�o?Fm��v�!K�USB��=Hn	�f�!STM�0��;JoU����O�֟�c����CICE�_KL ?%K� (%SVCPRG1��G�1���c�FN�G3o�t�6�4��D��6�5��į6�6��6�7��6���W�R�9_�d�3��� 6�9���6�a�ܿ6��� �6���,�6�ٯT�6� �|�6�)���6�Q��� 6�y���^����^�ʿ D�^��l�^�ϔ�^� Bϼ�^�j���^���� ^���4�^���\�^�
� �2���6��/� ���V��<�'�`�K� ��o����������� ��&J5nY� ������� 4F1jU�y� ����/�0// T/?/x/c/�/�/�/�/ �/�/�/??>?)?P?�t?_?�?
�_DEV� I�M{C:�84���4?GRP 2/E�0�+�bx 	�/ 
 ,@�?O ��ODO+OhOOOaO�O �O�O�O�O�O�O__ @_R_9_v_]_�_�_O �_�_�_o�_*ooNo `oGo�oko�o�o�o�o �o�o&8\�_ Q�I����� ��4�F�-�j�Q��� ����ď���Ϗ�� uB�T�;�x�_����� ��ҟ����ݟ�,�� P�7�t���m�����ί �7����(�:�!�^� E�����{�����ܿÿ տ���6��Z�l�S� ��篅���}������  ��D�+�h�z�aߞ� �����߻������� �R��v��o��� ��������*��N� `�G���k��������� ��k�8��\n U�y����� �	F-jQ� ������/ /B/T/;/x/_/�/�/ �/�/�/�/?�/,??�P?7?I?�?�3d ��6	t?�?�?�?�?O�?)O8K%�8O]O����vA"AvE�O �G~O�O�O�O�O�O
Y JO/_rI�O\_J_�_n_ �_�_�_�__o@_�_ 4o"oXoFo|ojo�o�_ o�oo�o�o0 TBx�o��oh� d���,��P�� w��@�����Ώ��ޏ ��(�j�O������ p�����ʟ��ڟ �B� '�f��Z�H�~�l��� ��Ư������د��  �V�D�z�h����ſ �������
��R� @�vϸ���ܿf��Ͼ� �������Nߐ�u� ��>ߨߖ��ߺ�����  �V�|�M��&��n� ��������.��R� ��F���V�|�j����� �����*���B 0Rxf���� ���>,N t���d��� �//:/|a/s/*/ L/&/�/�/�/�/�/? T/9?x/?l?Z?|?~? �?�?�?�?,?OP?�? DO2OhOVOxOzO�O�O O�O(O�O_
_@_._ d_R_t_�O�O�_ _�_ �_�_oo<o*o`o�_ �o�_Po�oLo�o�o�o 8zo_�o(� �������R 7�v �j�X���|��� ���*��N�؏B� 0�f�T���x�����՟ 矞������>�,�b� P���ȟ���v��ί ���:�(�^����� įN�����ܿʿ��  �6�x�]Ϝ�&ϐ�~� �Ϣ�������>�d�5� t��h�Vߌ�z߰ߞ� �����:���.���>� d�R��v������� �����*��:�`�N� �������t����� ��&6\����� L������" dI[4|� ����<!/`� T/B/d/f/x/�/�/�/ /�/8/�/,??P?>? `?b?t?�?�/�??�? O�?(OOLO:O\O�? �?�O�?�O�O�O _�O $__H_�Oo_�O8_�_ 4_�_�_�_�_�_ ob_ Go�_ozoho�o�o�o �o�o�o:o^o�oR @vd���� �6�*��N�<�r� `������Ϗ������ ��&��J�8�n����� ԏ^�ȟ��؟ڟ�"� �F���m���6����� į��ԯ֯��`�E� ���x�f��������� п&�L��\���P�>� t�bϘφϼ�����"� ��ߨ�&�L�:�p�^� ���ϻ��τ������  �"�H�6�l�ߓ��� \������������ D���k���4������� ������
L�1C�� ��d����� $	H�<*LN `����� � //8/&/H/J/\/�/ ��/��/�/�/?�/ 4?"?D?�/�/�?�/j? �?�?�?�?O�?0Or? WO�? O�OO�O�O�O �O�O_JO/_nO�Ob_ P_�_t_�_�_�_�_"_ oF_�_:o(o^oLo�o po�o�o�_�oo�o  6$ZH~�o� �n�j���2�  �V��}��F����� ��ԏ
���.�p�U� �����v��������� П�H�-�l���`�N� ��r��������4�� D�ޯ8�&�\�J���n� ���˿
�������� 4�"�X�F�|Ͼ���� l���������
�0�� Tߖ�{ߺ�D߮ߜ��� �������,�n�S�� ��t�������� 4��+������L��� p����������0��� $46H~l� ������  02Dz���j ����/
/,/� �y/�R/�/�/�/�/ �/�/?Z/??~/?r? ?�?�?�?�?�?�?2? OV?�?JO8OnO\O~O �O�O�O
O�O.O�O"_ _F_4_j_X_z_�_�O �__�_�_�_ooBo 0ofo�_�o�oVoxoRo �o�o�o>�oe �o.������ ��X=�|�p�^� �����������0�� T�ޏH�6�l�Z���~� ������,�Ɵ �� D�2�h�V���Ο��� |��x����
�@�.� d�����ʯT������ п���<�~�cϢ� ,ϖτϺϨ������� �V�;�z��n�\ߒ� �߶ߤ�������� ����4�j�X��|�� ����������� 0�f�T��������z� ������,b �����R���� �j�a�: ������ /B '/f�Z/�j/�/~/ �/�/�//�/>/�/2?  ?V?D?f?�?z?�?�/ �??�?
O�?.OORO @ObO�O�?�O�?xO�O �O_�O*__N_�Ou_ �_>_`_:_�_�_�_o��_&oh_Mo�_�Q�$�SERV_MAI�L  �U�`�~rhOUTPUT�h_�P@vd�RV 20f  �` (a\o�ovd�SAVE�l�iTO�P10 21�i d �_HZl ~������� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d�v������� ��П�����*�<��euYPscFZ�N_CFG 2e�c�T�a�e~|�GRP 23���q ,B   �AƠ�QD;� B}Ǡ�  B4�S�RB21�fH7ELL�4ev��`�o��/�>�%RSR>�?�Q���u� ����ҿ������,π�P�;�t�_Ϙϩ�~���  � �����Ϸͻ��P��&�'�ސW��2Pd��g��HKw 15�� ,� �߫ߥ��������� @�;�M�_���������������OMM� 6��?��FT?OV_ENB�d�a�u�OW_REG�_UI_�tbIMI_OFWDL*�7.��ɥ��WAIT\� `ٞ����`���d��wTIM�������VA�`����_UNcIT[�*yLCy�WTRY��uv`ME�8���aw�rdt ��9� ������<���X�Pڠ6p`?� � ��o+=1`VL�l�f�MON_ALIA�S ?e.��`heGo������ /)/;/M/�q/�/�/ �/�/d/�/�/??%? �/I?[?m??�?<?�? �?�?�?�?�?!O3OEO WOO{O�O�O�O�OnO �O�O__/_�OS_e_ w_�_�_F_�_�_�_�_ �_o+o=oOoaoo�o �o�o�o�oxo�o '9�o]o��> ������#�5� G�Y�k��������ŏ ׏������1�C�� g�y�����H���ӟ� ��	���-�?�Q�c�u�  �������ϯᯌ�� �)�;��L�q����� ��R�˿ݿ��Ͼ� 7�I�[�m��*ϣϵ� �����ϖ��!�3�E� ��i�{ߍߟ߱�\��� ��������A�S�e� w��4�������� ���+�=�O���s��� ������f����� '��K]o��> �����#5 GY}�����l�$SMON_�DEFPROG �&����� &*S?YSTEM*����RECALL �?}� ( ��}-copy f�rs:*.dt �virt:\te�mp\=>192�.168.56.�1:36372 �q%�/�/�/�/}
x�yzrate 11 V/h/z/??/?�%�'�/�!�/�/�?�?�?�"8K&ord�erfil.da~�&mpback�/p}?O#O5O }/K"mdbS *�?�?�?��O�O�O�$3xK$:\TO�@fOv0O_"_4_� 4�Ea�O�Oq5  _�_�_�_�?�?cO~O o!o3oFO�_jO�_�o �o�o�OW_i_�O /B_�o�ox_�����'tpdisc 0kv0hz���/��%tpconn 0 ����� ����@��sS�e�w�� �,��_�_Zo�_���� ��=oOoj�so��(� �o�o`�o7�����9 K\���$�6��* ֯���������B?T?400 j�|��� 1��ؿ����ϝϯ� B�T�f�x�	��-�@� �!�����ϋߝ߯�¿ Կ�x�	��-�@��! �����ߋ������� f�x�	��-�@�R�۟ ���������̟g��� {�0C���h��� �����ǯXj�� �#5H���� �����nj|/ /1/D�����/�/ �/B(���d/v/?? +?>�P���t��?�?�? ����i?��OO'O: L_pO�O�O8O� [OmO�O_#_5_H?Z? �?�?�_�_�_�?a_�?�|_oo1oDR�$S�NPX_ASG �2:���Va?� � DP�%�7o~o  ?��GfPARAM �;Ve`a �U	lkP>TDP>X~�d� ��I`�OFT_KB_CFG  CS\eFc�OPIN_SIMW  Vk�b+�=OYsI`RVNO�RDY_DO  ��eukrQST_P_DSB~�b|�>kSR <Vi� � & TELEO�e�{v>T�W`I`TOP_ON�_ERRxGb�P_TN VeP���D:�RIN�G_PRM'��rV�CNT_GP 2�=Ve�ac`x 	 ���DP��я����Bg�VD�RP 1>�i�`�Vq؏0�B� T�f�x���������ҟ �����,�>�e�b� t���������ί�� �+�(�:�L�^�p��� ������ʿ�� �� $�6�H�Z�l�~ϐϷ� ����������� �2� D�V�}�zߌߞ߰��� ������
��C�@�R� d�v��������� 	���*�<�N�`�r� �������������� &8J\n�� ������" 4[Xj|��� ����!//0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�?�O�PRG_CO7UNT�f�P�)I'ENBe�+EMUC�d�bO_UPD 1?>�{T  
ODR �O�O�O�O�O__A_ <_N_`_�_�_�_�_�_ �_�_�_oo&o8oao \ono�o�o�o�o�o�o �o�o94FX� |������� ��0�Y�T�f�x��� �����������1� ,�>�P�y�t������� ��Ο��	���(�Q� L�^�p���������� ܯ� �)�$�6�H�q� l�~�������ƿؿπ��� �I�D�V�"L_INFO 1@�E��@��	 �yϽϨ����ɿ��z�>�3=��n��w~�� �@k�?���@i*,�]/�H��r��
=�q��  ?�` �>@��i� �D�C�Ҭ��D	�1���@�G���Y��p߂�-@YSDEBSUG:@�@�o�d�I���SP_PASS�:EB?��LOG� A���A  �o�i�v�  ��Ao�UD1:�\��}���_MPC �ݚEk�}�A&��� �AK�SAV �B��IA���*�i��1�SVB�TEM�_TIME 1C����@ 0o���i�#�+��"���ME?MBK  �EA��������X�|�@� V�i�����������h�,9
�� ��@�a s���ϻ���nà@Rd�v�����
Le �//(/:/L/^/p/ �/�/�/�/�/�/�/ ?�?$?6?H?Z?��SK V�[�EAj��?�?�?��+:o�X]2���?
i� �po��
:O .@R�O�O�O}N�o�� ��OBi���?_&_8_,M2�Y_�_�_�_�_�_o�$�_�_�o'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk�_?T1SVGUNwSPD�� '�����p2MODE_?LIM D���2�t2�p�qE�݉u�ABUI_DCS' H}5���0�G ��D�D��|-�X�>�ލ�*���� 
��e��i���r�i������uEDI�T I��xSC_RN J���rS�G K�.�(���0߅SK_OPT�ION��^����_�DI��ENB  ��E���BC2_�GRP 2L��0���&AMPC�ʓ�|/BCCF/�N����c ����`� >�W�B�g���x����� կ��������S� >�w�b���������Ͽ �����=�(�a�L� �ϗ�Ň�϶������� v��
�/�U�@�yߧ� ��`�iМ��߰����� 
���.��>�@�R�� v����������� *��N�<�r�`����� ����������̀ 4FX��|j�� �����B 0fTvx��� ��/�,//</b/ P/�/t/�/�/�/�/�/ �/�/(??L?d?v? �?�?�?6?�?�?�?O  O6OHOZO(O~OlO�O �O�O�O�O�O�O __ D_2_h_V_�_z_�_�_ �_�_�_
o�_.oo>o @oRo�ovo�ob?�o�o �o�o<*Lr `������� �&��6�8�J���n� ����ȏ���ڏ��"� �F�4�j�X���|��� �����֟��o$�6� T�f�x���������ү �������>�,�b� P���t��������ο ��(��L�:�\ς� pϦϔ��ϸ�������  ��H�6�l�"��ߖ� ������V������2�  �V�h�z�H����� ����������
�@�.� d�R���v��������� ����*N<^ `r������� &8�\Jl� �������"/ /F/4/V/X/j/�/�/ �/�/�/�/?�/?B? 0?f?T?�?x?�?�?�? �?�?O�?,O�DOVO tO�O�OO�O�O�O�O��O_ V4P�$TB�CSG_GRP �2O U��  �4Q 
 ?�  __q_[_ �__�_�_�_�_�_o�%k8R?SQF\dאHTa?4Q	 �HA���#e>�w��>$a�\#e?AT��A WR�o��hdjma�G�?L�fg�bp�o�n�ff�hf��ͼb4P|j���o*}@��Rhf�?ff>�33pa#eB<qB�o+=xrRp�qUy�rt~��H`�y rIpTv�pBȺ t~	xf	x(�;��� f���N�`���ˏڋ�����	V3.0�0WR	crxlڃ	*��3R~td��HH��� \��.�]�  cC�.�����8QJ2?SR�F]����CFG [T UPQ SPVܚ��r�ܟ1��1�W�e�	P e���v�����ӯ���� ����Q�<�u�`� ��������Ϳ�޿� �;�&�_�Jσ�nπ� �Ϥ�������WRq@ �0�B���u�`߅߫� ���ߺ������)�;� M��q�\������ 4Q _���O ���J� 8�n�\����������� ������4"XF hj|����� �.TBxf ��nO����/ />/,/b/P/�/t/�/ �/�/�/�/�/�/?:? (?^?p?�?�?N?�?�? �?�?�?�? O6O$OZO HO~OlO�O�O�O�O�O �O�O __D_2_T_V_ h_�_�_�_�_�_�_
o �_o@o�Xojo|o&o �o�o�o�o�o�o* N`r�B�� �����&��6� \�J���n�����ȏ�� ؏ڏ�"��F�4�j� X���|���ğ���֟ ���0��@�B�T��� x�����ү䯎o��� ̯ʯP�>�t�b����� ���������Կ&� L�:�p�^ϔϦϸ��� ������� �"�H�6� l�Zߐ�~ߴߢ����� �����2� �V�D�z� h������������ �
�,�.�@�v��� ����\������� <*`N���� x���8J \(����� ���/4/"/X/F/ |/j/�/�/�/�/�/�/ �/??B?0?f?T?v? �?�?�?�?�?�?OO ��2ODO�� O�OtO�O �O�O�O�O_�O(_:_ L_
__�_p_�_�_�_ �_�_ o�_$oo4o6o Ho~olo�o�o�o�o�o �o�o D2hV �z�����
� �.��R�@�b���v� ��&OXO֏菒���� �N�<�r�`������� ̟ޟ🮟��$�&� 8�n�������^�ȯ�� �گ��� �"�4�j� X���|�����ֿĿ� ���0��T�B�x�f� �ϊϜ���������� �>�P���h�zߌ�6� �ߪ����������:� (�^�p���R���p���� ���  &��*� *�>�*���$TBJOP_G�RP 2U����  ?_���C*�	V��]�Wd������X  �*��� �,? � ���*� @&�?��	� �A�����C�  DD������>v�>\?� ��aG�:��o��;ߴAT3������A�<���MX����>��\�)?���8Q������L��>̼0 &�;iG.���Ap< � F�A�ff�v��� �):VM�.��� S>o*�@��R�Cр	����p�����ff��:�6/�?�3=3�B   �� /������>)/:�S���� <�/�/@��H�%&/и/��=� <#��
*��v�;/��ڪ!?���4B� 3?'?2	��2?hZ? D?R?�?�?�?F?�?�? �?�?OAOO�?`OzO`dOrO�O�O*�C�*����A��	V3.�00{�crxl��*P��%�%c�5Z F� �JZH F6� �F^ F�� �F�f F� �G� G5 �G<
 G^] �G� G����G�*�G�S G�; G��ER�Du�\E[� �E� F( �F-� FU` �F}  F�N �F� F�� �Fͺ F� �F�V G� �Gz Ga O9ѷ�Q�LHe�fJ4�o,b*��0c1���OH�ED_?TCH Xd�+X�2S�&�&�dA$'X�o�o*�1F��TESTPARS�  ��cV�HR�pABLE 1Yd� N`*����R�g$j�g�h�h�)�1��g	�h
�h��hHu*��h�h:�h%vRDI0n�GYk}��u	�O�#�-�?�Q�c�u�)rS�l� �z6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z���I���m�Fwͩ ��ȏڏ쏘������x)r��NUM [ ��n����2� Ep�)r_CFG Z��I����@V�IMEBF_�TTqD��e޶V�ER�����޳R� 1[8{ 8$�o*�%�Q� ��د  9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}��ߡ߳� ����������1��� E�W�i�{������ ��������/�A�S� e�w����������������+=O�_Ԗ��@��`LIoF \��D`B����DR�(FP�
�!p�!p� �d� ��MI_CH�AN� � D_BGLVL��f�ETHERAD� ?u��0`�1�_}�ROUmT�!�j!���SNMASK�Y�j255.�%S///A/S�`O�OLOFS_DI�p�CORQC?TRL ]8{��1o�-T�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OL�/6O�%OZOcPE_DE�TAI7�*PGL�_CONFIG �c������/�cell/$CID$/grp1^O@�O�O�O
__|��� G_Y_k_}_�_�_0_�_ �_�_�_oo�_CoUo goyo�o�o,o>o�o�o �o	-�oQcu ���:���� �)���_�q���������׮}N�����%�7�I�a�KOq�P�� M�����ʟܟ� �G� $�6�H�Z�l�~���� ��Ưد������2� D�V�h�z������¿ Կ���
ϙ�.�@�R� d�vψϚ�)Ͼ����� ���ߧ�<�N�`�r� �ߖ�%ߺ�������� �&��J�\�n��� ��3����������"� ��F�X�j�|���������@�User� View �I}�}1234567890����+`=Ex �e����2��B������`r��3�Oa�s����x4 >//'/9/K/]/�~/x5��/�/�/�/ �/?p/2?x6�/k? }?�?�?�?�?$?�?x7Z?O1OCOUOgOyO�?�Ox8O�O�O�O�	__-_�ON_TR �lCamera���O�_�_�_�_�_�_˂E�_o)o;n ��Uogoyo�o�o�o�)  mV�	�_�o# 5GY o}���o�������F_� mV=�k�}������� ŏl����X�1�C� U�g�y���2�D��"� ן�����1�؏U� g�y�ğ������ӯ� ����D��k��E�W�i� {�����F�ÿտ�2� ��/�A�S�e��nU Y9������������	� ��-�?�Qߜ�u߇ߙ� �߽���v�D�If�� -�?�Q�c�u�ߙ�� ���������)�;� ��D��I��������� ������)t�M�_q���N�`�9 3��0B�� Sx�1����P�//�J	oU0� U/g/y/�/�/�/V�/ �/�/�?-???Q?c? u?/./tPv[?�?�? �?OO(O�/LO^OpO �?�O�O�O�O�O�O�? oU�k�O:_L_^_p_�_ �_;O�_�_�_'_ oo $o6oHoZo_;%N��_ �o�o�o�o�o �_$ 6H�ol~��� �moe��]�$�6� H�Z�l�������� ؏���� �2��e &�ɏ~�������Ɵ؟ ���� �k�D�V�h� z�����E�e��5�� ��� �2�D��h�z� ��ׯ��¿Կ���
���  ��9�K� ]�oρϓϥϷ�����<����   �� 5�G�Y�k�}ߏߡ߳� ����������1�C� U�g�y�������� ����	��-�?�Q�c� u��������������� );M_q��  
��(  }�-�( 	 � ������# 35G}k���:�
� �Y�
/ /./��R/d/v/�/�/ �/����/�/�/A/? 0?B?T?f?x?�/�?�? �??�?�?OO,O>O �?bOtO�O�?�O�O�O �O�O_KO]O:_L_^_ �O�_�_�_�_�_�_#_  oo$ok_HoZolo~o �o�o�_�o�o�o1o  2DVh�o�o� ��	��
��.� @��d�v�������� Џ���M�*�<�N� ��r���������̟� %���&�m�J�\�n� �������ȯگ�3� �"�4�F�X�j����� ������ֿ����� 0�w���f�xϊ�ѿ�� ���������O�,�>� Pߗ�t߆ߘߪ߼��� �����]�:�L�^��p����߻@  ����������� ���"frh:\�tpgl\robots\crx!��10ia_l.xml��D�V�h�z������������������ ��0BTfx� �������� ,>Pbt��� �����/(/:/ L/^/p/�/�/�/�/�/ �/��/?$?6?H?Z? l?~?�?�?�?�?�?�/ �?O O2ODOVOhOzO �O�O�O�O�O�?�O
_ _._@_R_d_v_�_�_ �_�_�_�O�_oo*o <oNo`oro�o�o�o�o��o�n �6� |���<< 	� ?��k!�o; iOq����� ����%�S�9�k�@��o�����я�����(�$TPGL_�OUTPUT �f������ �&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��������į�p�ր2�345678901�����1�C�K� ���r���������̿ d�п��&�8�J��}T�|ώϠϲ���\� n�����0�B�T��� bߊߜ߮�����j��� ��,�>�P����߆� ��������x���� (�:�L�^���l����� ������t���$6 HZlz��� ���� 2DV h ����� ��/./@/R/d/v/ /�/�/�/�/�/�/�/~ۂ $$�� ί<7*?\?N?�?r?�? �?�?�?�?�?OO4O &OXOJO|OnO�O�O�O �O�O�O_�O0_"_T_}�an_�_�_�_�_�_��]@�_o	z ( 	 V_Do2o hoVo�ozo�o�o�o�o �o
�o.R@v d������� ��(�*�<�r�`����ܦ�  <<I_ˏݏ����� ��:�L�֪��}���)� ��ş�������k�� C�ݟ/�y���e����� ��������-�?�� c�u�ӯ]�����W�� �Ϳ��)χ���_�q� �yϧρϓ�����M� �%߿��[�5�Gߑ� ��߫���s����!� ��E�W��?���9� ��������i���A� S���w���c�u���� /�����=) s�����U�� �'9�!o	 [�����K� #/5/�Y/k/E/w/�/ �/�/�/�/�/?�/ ?U?g?�/�?�?7?�?��?�?�?	OO��)�WGL1.XML��_PM�$TPOF?F_LIM ���P����^FNw_SVf@  �T�xJP_MON �g��zD�P��P2ZISTRTC�HK h��xF�k_aBVTCOMP�AT�HQ|FVWV_AR i�M:X.�D �O R_�P��BbA_DEFPROG %�I�%TELEO�P Pi_VM_DISPLAYm@�N�R�INST_MSK�  �\ �ZI�NUSER_�TL�CKl�[QUIC�KMEN:o�TSC�REY`��Rtpsc�Tat`hyixB�`_�iSTZ�xIRACE_CF�G j�I:T��@	[T
?��hHNL 2k�Z���aA[ gR-?Qcu�����z�eITE�M 2l{ ��%$123456�7890 ��  �=<
�0�B�J�  #!P�X�dP��� [S���"���X�
� |���W���r�֏���� .��0�B�\�f����� 6�\�n�ҟ������ ��>���"���.��� ��ίR����Ŀֿ:� �^�p�9ϔ�Tϸ�x� ����d���H�� l��>�Pߴ�\����� ��v� ������h�(� �ߞ߰�4�L��ߦ�� ���@�R��v�6��� Z�l���������*� ��N��� �������� ����X���J 
n���b� ���"4F�/ |</N/�Z/���/ /�/0/�/?f/?�/ �/e?�/�?�/�?�?�? ,?�?P?b?t?�?�?DO jO|O�?�OOO(O�O �O^O_0_�O<_�O�O �_�O�__�_�_H_�_Pl_~_Go�dS�bm�o>Lj�  �rLj� �a�o�Y
 �o�o�o�o{jUD�1:\|��^aR_GRP 1n�{�� 	 @ �PRd{N�r����~��p���q�+��O�:�?�   j�|�f���������� ҏ����>�,�b�P����t���������	�e���\cSCB ;2ohk U�R� d�v���������Я��RlUTORIAL� phk�o-�WgV�_CONFIG qhm�a�o�o��<��OUTPUT yrhi}����� ܿ� ��$�6�H�Z� l�~ϐϢϴ�z�ɿ�� �� ��$�6�H�Z�l� ~ߐߢߴ��������� � �2�D�V�h�z�� �����������
�� .�@�R�d�v������� ��������*< N`r������ ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/��/�/? ?0?B?T?f?x?�?�? �?�?�/�?�?OO,O >OPObOtO�O�O�O�O �?�O�O__(_:_L_ ^_p_�_�_�_�_�_f� x�ǿoo,o>oPobo to�o�o�o�o�o�o�O (:L^p� ������o �� $�6�H�Z�l�~����� ��Ə؏��� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ���*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b� t���������������>�X���# ��N�_r��� ����&8 J��n����� ���/"/4/F/X/ i|/�/�/�/�/�/�/ �/??0?B?T?e/x? �?�?�?�?�?�?�?O O,O>OPOa?tO�O�O �O�O�O�O�O__(_ :_L_^_oO�_�_�_�_ �_�_�_ oo$o6oHo Zok_~o�o�o�o�o�o �o�o 2DVgo z������� 
��.�@�R�d�u�� ������Џ���� *�<�N�`�q������� ��̟ޟ���&�8��J�\�k��$TX_�SCREEN 1}s% �}�k�����ӯ���	���Z��I�[� m�������,�ٿ� ���!�3Ϫ�W�ο{� �ϟϱ�����L���p� �/�A�S�e�w��� � �߿��������~�+� ��O�a�s���� � ��D�����'�9�K� ��������������� R���v�#5GYk�}����$UAL�RM_MSG ?5����� �n� ��	:-^Q c������ /~�SEV  ��2&�ECFG� u���� � n�@�  A�b!   B�n�
 /u����/�/�/ �/�/�/??%?7?I?�W7>!GRP 2v�H+ 0n�	 �/�?� I_BBL�_NOTE w�H*T���lu���w�T �2D_EFPRO� %� (%�Ow�	O BO-OfOQO�OuO�O�O��O�O�O_�O,_�<F�KEYDATA �1x���0p W'n��?�_�_z_�_��_�Z,(�_on�(�POINT  �]onc NCEL�@oko�PNDIRE�CTlono EXT� STEP�om?TOUCHU�o�o��PORE INFO�o�o0B)fM �����������>�P� ���/frh/gu�i/whitehome.pngQ�`������ŏ׏�h�pointz����/�A�S��  FR�H/FCGTP/�wzcancel ��������ʟܟk�i�indirec����'�9�K�]�h�z�nex�������ϯ���h�touchup���/�A�S�e���h�arwrg ������ÿտ�n�� �(�:�L�^�p����� �ϸ�������}��$� 6�H�Z�l��ϐߢߴ� �������ߋ� �2�D� V�h�z�	������� ������.�@�R�d� v���_����������� ���2DVhz ������
 �@Rdv�� )����//� </N/`/r/�/�/%/�/ �/�/�/??&?�/J? \?n?�?�?�?3?�?�? �?�?O"O�?4OXOjO |O�O�O�OAO�O�O�O __0_�OT_f_x_�_ �_�_=_�_�_�_oo ,o>o�_boto�o�o�o��oW��k�b�����o}�o8J$v,6�{.�� �������/� �S�:�w���p����� я�ʏ��+��O� a�H���l�������ߟ ���'�9�Ho]�o� ��������ɯX���� �#�5�G�֯k�}��� ����ſT������ 1�C�U��yϋϝϯ� ����b���	��-�?� Q���u߇ߙ߽߫��� ��p���)�;�M�_� �߃��������l� ��%�7�I�[�m��� ������������z� !3EWi���� �����П/ ASew~��� ���/�+/=/O/ a/s/�//�/�/�/�/ �/?�/'?9?K?]?o? �?�?"?�?�?�?�?�? O�?5OGOYOkO}O�O O�O�O�O�O�O__ �OC_U_g_y_�_�_,_ �_�_�_�_	oo�_?o Qocouo�o�o�o:o�o �o�o)�oM_ q���6������%�7�9�}����b�@t���^�������,�� 돞����3�E�,�i� P�������ß����� ����A�S�:�w�^� ������ѯ����ܯ� +�
O�a�s������� �Ϳ߿���'�9� ȿ]�oρϓϥϷ�F� �������#�5���Y� k�}ߏߡ߳���T��� ����1�C���g�y� ������P�����	� �-�?�Q���u����� ������^���) ;M��q���� ��l%7I [������ h�/!/3/E/W/i/ @��/�/�/�/�/�/� ??/?A?S?e?w?? �?�?�?�?�?�?�?O +O=OOOaOsOO�O�O �O�O�O�O_�O'_9_ K_]_o_�__�_�_�_ �_�_�_�_#o5oGoYo ko}o�oo�o�o�o�o �o�o1CUgy ������	� ��?�Q�c�u����� (���Ϗ������ ;�M�_�q�������~ ����~ ���ҟ���Ο�*��,�[���f��� ����ٯ�������3� �W�i�P���t���ÿ ���ο��/�A�(� e�Lωϛ�z/������ ����(�=�O�a�s� �ߗߩ�8�������� �'��K�]�o��� ��4����������#� 5���Y�k�}������� B�������1�� Ugy����P ��	-?�c u����L�� //)/;/M/�q/�/ �/�/�/�/Z/�/?? %?7?I?�/m??�?�? �?�?�?���?O!O3O EOWO^?{O�O�O�O�O �O�OvO__/_A_S_ e_�O�_�_�_�_�_�_ r_oo+o=oOoaoso o�o�o�o�o�o�o�o '9K]o�o� �������#� 5�G�Y�k�}������ ŏ׏������1�C� U�g�y��������ӟ ���	���-�?�Q�c� u��������ϯ��h���0���0���B�T�f�>�����t�,��˿~� �ֿ�%��I�0�m� �fϣϊ��������� ��!�3��W�>�{�b� �߱ߘ��߼�����? /�A�S�e�w��� ������������=� O�a�s�����&����� ������9K] o���4��� �#�GYk} ��0����/ /1/�U/g/y/�/�/ �/>/�/�/�/	??-? �/Q?c?u?�?�?�?�? L?�?�?OO)O;O�? _OqO�O�O�O�OHO�O �O__%_7_I_ �m_ _�_�_�_�_�O�_�_ o!o3oEoWo�_{o�o �o�o�o�odo�o /AS�ow��� ���r��+�=� O�a����������͏ ߏn���'�9�K�]� o���������ɟ۟� |��#�5�G�Y�k��� ������ůׯ����� �1�C�U�g�y���� ����ӿ������-�@?�Q�c�uχ�^P����^P���������ͮ���
���, ��;���_�F߃ߕ�|� �ߠ����������7� I�0�m�T������ �������!��E�,� i�{�Z_���������� ���/ASew ������ �+=Oas� �����//� 9/K/]/o/�/�/"/�/ �/�/�/�/?�/5?G? Y?k?}?�?�?0?�?�? �?�?OO�?COUOgO yO�O�O,O�O�O�O�O 	__-_�OQ_c_u_�_ �_�_:_�_�_�_oo )o�_Mo_oqo�o�o�o �o���o�o%7 >o[m���� V���!�3�E�� i�{�������ÏR�� ����/�A�S��w� ��������џ`���� �+�=�O�ޟs����� ����ͯ߯n���'� 9�K�]�쯁������� ɿۿj����#�5�G� Y�k����ϡϳ����� ��x���1�C�U�g� �ϋߝ߯�����������`����`���"�4�F��h�z�T�,f���^���� �����)��M�_�F� ��j����������� ��7[B� x�����o! 3EWixߍ�� �����///A/ S/e/w//�/�/�/�/ �/�/�/?+?=?O?a? s?�??�?�?�?�?�? O�?'O9OKO]OoO�O O�O�O�O�O�O�O_ �O5_G_Y_k_}_�__ �_�_�_�_�_o�_1o CoUogoyo�o�o,o�o �o�o�o	�o?Q cu��(��� ���)� M�_�q� �������ˏݏ�� �%�7�Ə[�m���� ����D�ٟ����!� 3�W�i�{������� ïR������/�A� Яe�w���������N� �����+�=�O�޿ sυϗϩϻ���\��� ��'�9�K���o߁� �ߥ߷�����j���� #�5�G�Y���}��� ������f�����1��C�U�g�>�i��>>�������� ����������,� �?&cu\�� �����) M4q�j��� ��/�%//I/[/ :�/�/�/�/�/�/�� �/?!?3?E?W?i?�/ �?�?�?�?�?�?v?O O/OAOSOeO�?�O�O �O�O�O�O�O�O_+_ =_O_a_s__�_�_�_ �_�_�_�_o'o9oKo ]ooo�oo�o�o�o�o �o�o�o#5GYk }������ ��1�C�U�g�y��� �����ӏ���	��� -�?�Q�c�u�����p/ ��ϟ�����;� M�_�q�������6�˯ ݯ���%���I�[� m������2�ǿٿ� ���!�3�¿W�i�{� �ϟϱ�@�������� �/߾�S�e�w߉ߛ� �߿�N�������+� =���a�s����� J�������'�9�K� ��o�����������X� ����#5G��k�}���������������&�HZ4,F/�>/���� �	/�-/?/&/c/J/ �/�/�/�/�/�/�/�/ ?�/;?"?_?q?X?�? |?�?�?���?OO%O 7OIOXmOO�O�O�O �O�OhO�O_!_3_E_ W_�O{_�_�_�_�_�_ d_�_oo/oAoSoeo �_�o�o�o�o�o�oro +=Oa�o� �������� '�9�K�]�o������ ��ɏۏ�|��#�5� G�Y�k�}������ş ן������1�C�U� g�y��������ӯ� ��	��?-�?�Q�c�u� ��������Ͽ��� Ϧ�;�M�_�qσϕ� $Ϲ��������ߢ� 7�I�[�m�ߑߣ�2� ���������!��E� W�i�{���.����� ������/���S�e� w�������<������� +��Oas� ���J�� '9�]o��� �F���/#/5/�G/�$UI_IN�USER  ����h!��  H/L/_�MENHIST �1yh% � (u  �)�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,1133,A1�/�/??�'�/�.71�/{?�?�?�?��+E?�%edit~�"TELEOPj?@OO'O�?D?V?2�/ �O�O�O�O�(MO�/48,2�O
__._x@_�/�O,163i?��_�_�_�_Q_c_uR2 {_o"o4oFo�O�_�!�5qO�o�o�o�o�����!�a�o�o!3EW �o|�� ���e���0� B�T��x��������� ҏ�s���,�>�P� b�񏆟������Ο�� o���(�:�L�^�p� ��������ʯܯ��o �$�6�H�Z�l�~��� ����ƿؿ����� � 2�D�V�h�z�	Ϟϰ� ��������
ߙ�.�@� R�d�v߈�߬߾��� ������*�<�N�`� r���%�������� �����J�\�n��� �������������� "��FXj|�� /����0 �Tfx���= ���//,/�=/ b/t/�/�/�/�/K/�/ �/??(?:?%��/p? �?�?�?�?�?�/�? O O$O6OHO�?lO~O�O �O�O�O�OgO�O_ _ 2_D_V_�Oz_�_�_�_ �_�_c_�_
oo.o@o Rodo�_�o�o�o�o�o �oqo*<N`�K;�$UI_PA�NEDATA 1�{����q�  	�}�  frh/cg�tp/flexd�ev.stm?_�width=0&�_height=�10�p�pice=�TP&_line�s=15&_columns=4�p�font=24&�_page=wh�ole�pmI6) � rim�9�   �pP�b�t�������� ����Ǐ��(�:�!� ^�E�����{�����ܟ��՟�I6� ��    	 :�J�O�a�s� ��������ͯ@��� �'�9�K���o���h� ����ɿۿ¿���#� 5��Y�@�}Ϗ�vϳ�&��Ɠs����� )�;�Mߠ�q�䯕ߧ� ��������V��%�� I�0�m��f����� ��������!��E�W� ���ύ����������� :�~�/ASew ������  =$asZ� ~����d�v�'/ 9/K/]/o/�/��/�/ *�/�/�/?#?5?�/ Y?@?}?�?v?�?�?�? �?�?O�?1OCO*OgO NO�O�/�/�O�O�O 	__-_�OQ_�/u_�_ �_�_�_�_6_�_o�_ )ooMo_oFo�ojo�o �o�o�o�o�o%7 �O�Om���� �^_�!�3�E�W� i�{������Ï��� ������A�S�:�w� ^�������џDV� �+�=�O�a������� 
���ͯ߯���|� 9� �]�o�V���z��� ɿ���Կ�#�
�G�0.�k�ޟ�}�|ϵ� ���������)��4� ��#�`�r߄ߖߨߺ� !����������8�� \�C���y������������������$�UI_POSTY�PE  ��� 	 ��s�B�QUICKM_EN  Q�`��v�D�RESTOR�E 1|���  ��*default���  INGL�E��PRIM���meditp�age,TELEOP,1Sew �,������ �/ASe��� z������/ !/�E/W/i/{/�/0/ �/�/�/�/�/�?? *?�/e?w?�?�?�?P? �?�?�?OO+O�?OO aOsO�O�OB?�O�O�O :O__'_9_K_�Oo_ �_�_�_�_Z_�_�_�_ o#o�O�_BoTo�_xo �o�o�o�o�o�o 1CU�oy�����{�SCRE��?���u1s]c��u2�3�U4�5�6�7��8��sTATM��� ����:�USE�R�p��rT�p�k�s���4��5��6ʝ�7��8��B�ND�O_CFG }�Q�����B�PDE����Non�e��v�_INFOW 2~��)���0%�D���2�s�V� ������͟ߟ�� '�9��]�o�R���z���OFFSET �Q�-���hs�� p�����G�>�P� }�t���Я��׿ο� ���C�:�L�^Ϩ����͘���
����av���WORK �!�����.�@ߢ��u�UFRAM ����RTOL_�ABRT�����E�NB�ߣ�GRP �1�����Cz  A������ *�<�N�`�r��֐��U�����MSK � �)���N���%!��%z����_'EVN�����+�vׂ3�«
 h��UEV��!�td:\event_user\�Fu�C7z���jpF���n�SPs�x�sp�otweld��!C6��������!���G|'��5 kY����� >���1�U g���/��	/ ^/M/�/-/?/�/c/�/ �/�/�/$?�/H?�/:�J�W�3�����8C?�?�? �?�?�? �?O+OOOOaO<O�O �OrO�O�O�O�O_�O '_9__]_o_J_�_�_��_�$VALD_�CPC 2�« ��_�_� w��qd�R�*o_oqo��hsNbd�j�`�� �i�da{�oav�_�oo o3BoWi{�o�o �o�o��o�P A�0�e�w����� �����(�=�L� a�s�
�������ʏ�� ���$�ޟH�:�o� ��������ڟ؟��� �� �2�G�V�k�}��� ����¯ԯ����� .��R�S�yϋϚ��� �������	��*�<� Q�`�u߇ߖϨϺ��� ������&�8�M�\� q���߶���n��� ���"�4�F�[�j�� �������������� !0�B�Wf�{�� ���������, >teT���� ���/+/:L a/p�/�/./��� ��//'?6/H/?l/ ^?�?�?�/�/�/�/�/ ?#O�?D?V?kOz?�O �O�?�?�?�?�?_O 1_@ORO9_vOw_�_�_ �O�O�O_�__-o<_ N_`_uo�_�o�o�_�_ �_�_o&o;Jo\o q�o����o�o�o � �"7�FXj� ���������� !�0�E�T�f�{����� ��ßҏ����
�,� A�P�b�����x����� Ο�����(�*�O� ^�p���������R�ܯ � ��Ϳ6�K�Z�l� &ϐ��Ϸ���ؿ��� "� �2�G���h�zϏ� �ϳ���������
�� 1�@�U�d�v�]�ߛ� ���������,��<� Q�`�r�������� ������&�;J�_ n����������� ���$F[j| ������� 0E/Ti/x��/ ��/�/�/�//,/ .?P/e?t/�/�/�?�? �?�?�/??(?:?L? NOsO�?�?�O�?�O�O vO OO$O6O�OZOo_ ~O�OJ_�O�_�_�_�O�_ _F_D_V[�$V�ARS_CONF?IG ��Pxa�  F�P]S�\lCMR_GRP 2�xk' ha	`�`�  %1: S�C130EF2 �*�o�`]T�VU�P��h`�5_Pa?_�  A@%pp*`��Vn No9x CVXdv��a��N<uA�%p�q�_R���_R B���#�_Q'��H� �l�;���{�����؏ ÏՏ�e��D�/�A��z�-�����ddIA_WORK �xe�ܐ�Pf,	�	�Qxe���G�P� ���YǑRTS�YNCSET  �xi�xa-�WIN?URL ?=�`�����������ȯ�گSIONTM�OU9�]Sd� ���_CFG ��S۳�S۵�P�` FR�:\��\DATA�\� �� �MC3�LOG@� �  UD13�E�Xd�_Q' B@ ����x�e_�ſx�ɿ�VW �� n6  ���VV��l�q?  =���?�]T�<�y�Y�TRAI�N���N� 
g!p?�CȞ��TK��:�b�xk (g��� ��_���������U� C�y�g߁ߋߝ߯���\���_GE��xk7�`_P�
�P�R,ꋰRE��xe*�.`hLEX�xl`�1-e�VMPH?ASE  xec��ecRTD_F�ILTER 2�.xk �u�0�� ��0�B�T�f�x��� ��VW�������� �$6HZl_iSH�IFTMENU {1�xk
 <�\1%�������� ��=&sJ \��������'/�	LIVE�/SNA�c%v�sfliv��9/�+�� 7�U�`\"menur/w//�/��/�����]��M�O��y��5`h`Z%D4�V�_Q<��0���$WAITDINEND��a2p6OK  �i�<��r�?S�?�9TIM�����<Gw?M�?�*K�?
J�?
J�?�8RELE��:G6p3��<�r1_ACTO 9Htܑ�8_<� �ԙ��%�/:_af�BRD�IS�`�N�$X�VR��y��$oZABC�b1�S;� ,��j�I�2�B_ZmI1�@VSPT� �y��eG�
�*�/o�*!o7o��WDCSCHG ��ԛ(��P\g@m�PIPL2�S?�i��o�o�o�ZMPCF_G 1��ii�0'¯S;Ms�Si��i��p'��g��e2��  ?�}Wν�s������I��~ꞽ-M���C�=TH��}�)D�C�Ҭ�D	I��1�҃ĝ<Ŧ��=�9H�w�п����jYc��ur��p�pUG�t�p��p�x���p���}P����Z�~���Ï��y��1��@�G��G�Y�ڈE�ꄙ��҉�����*�@��N�x��vv�L�R���2���d���x�}���܏��@=���7�{"�Þ��B��DL�W�I�&���B.�g�L�?����=k�5�q? �glp����o�_CYLI�ND�� { ���� ,(  * =�N�G�:�w�^����� ��ѯ���7�� ��<�#�5�r������� ����޿y�_����8�@ύ�nπ�㜻ã wQ �5�����S �����(�ٻ�X���r�A��SPH�ERE 2��� ҿ��"ϧ������P� c�>�P�̿t���ߪ� �����'���]�o� L���p�W�i�������������PZZ�F � 6