��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1RTU4QQ�Rx1R�� � $TIT91� ��� �Td��T0�ThP�T5�V6��V7�V8�V9�W0 �W�WOQ�U�WgQ�U�WU1�W1�W1�W1�W�2�R  �ASBoN_CF�!@$<!J� ; ;2�1�_CMNT�$�FLAGS]�C�HEK"$�b_O�PTJB6 � ELL�SETUP � `@HO8@9 P�R�1%�c#�aREPR�hu0D+�@���b{uHM9 MN�B;1 UTOB�J U�0 }49DEVIC�STI/@�� �@b3�4pB�d�"VAL��#ISP_UNI�tp_DOcv7�yFR_F�@|%u13���A0s�C_WAx�t,q�zOFF_T@]N�DEL�Lw0pdq�1�Vr?^q��#S?�o`Q"U��t#*�QTB����MO� �E �� [M�����R;EV�BIL����XI� v�R � !D�`��/$NOc`M�|���ɂ/#ǆ� �ԅ���1X�@Ded� p E RD_�E��h�$FSS�B6�`KBD_S�E�uAG� G�2BQ"_��2b�� V!��k5p`(��C 0q_E�D� � � �t2�$!S�p-D%$$� �#�B�ʀ�_OK1��0] P_�C� ʑ0t��U �`LACI�!�a�Y�<� �qCOMM� # $D
� ��@����J_\R��IGALL;OW� (Ku2:-B�@VAR���!�AB �BL�@� �� ,K�q���`S�p�@M_O]˥���CCFS_U	T��0 "�A�Cp'���+pXG��b�0 =4� IMCM ��#�S�p�9���i �_@�"t��6 ��M�1� h$�IMPEE_F�s��s��0� t����D_���J��D��F����q_����0 T@L��L�DI�s@G�^� �P��$I�'�� ��CFed X@G�RU@��Mb�NF�LI�\Ì@UIR�E�i42� SWIYTn$`0_N�`S 2�CF�0M� 	�#u�D��!��v`(����`J�tV��[ �E��.p�`�ʗELBOF� �շ �p`0���3����� F�2T��A`�rq1�J1��z _To!@��p��g���G�� �r0WARNM�p#tC�v`�ç` �� COR-UrF�LTR��TRAT�9 T%p� $AC�CVq��� ��r$�ORI�_&�RTr��S<��0CHG�0I���TW��A�I'�T��!D��� �202�a1���HDR�2��2�2JP; S���3��4��U5��6��7��8���9KD׀
 �2 ]@� TRQ�$vfh��'�1�<�_U<��G�]`COec  <� P�b�t�53>B_�LLEC��!~�MULTI�4�"u�Q|;2�CHILD���;1���@T� "'�STY92	r��=��)2�������ec# |r056$J� ђ��`���uT�O���E^	EXT�t����2��22Q"M����$`@D	��`&�ᣡ����� %�"��`%�ak�� ���s�����&'�E��Au��Mw�9 �%� ��TR�� ' L@U#9 ��z�At�$JOB�����P��}IG��( dp������^'�#j�~�L�pOR��) t$�FL��
RNG%Q@�TBAΰ �v&r�*`1t(@��0 �x!�0�+P�p��%ذ�`��*��@͐U��q�!�;2J�S_R��>�C<J�T8&<J D`5CF9����x"�@J��P_�p�7p+ \@RaO"pF�0��IT�s�0NOM��>Ҹ4s(�2�� @U<PPgў�P8,|Pn��0�1P�9�͗ RA���pl�?C�� �
$TͰ.tMD3�0T��pQU�`�΀+AHlr>�T1�JE�1\�J����PQ��\Q��hQCY�NT�P��PDBG�D̰�0-���PU�6$$Po�|�u�AX�����TAI�sB�UF,�]��A�1. �����F�`PI|�U-@PvWMuXM�Y��@�VFvWSIMQ�STO�q$KEE�SPA��  ?B�BP>C�BWQ��/�`�ˏMARG�u2�F�ACq�>�SLEW�*1!0����
��A_MCW$0'���p�JB�Ї�qDEC�j�e�s�V%1� Ħ�CHNR�MPs�$G_@�gD��_�@s��1_FP�5�@TC�fFӓC�� ����qC��+�VK�*���"*�JRx���SE7GFR$`IOh!�0;STN�LIN>�cs�PVZ�N�Ц@�D2 ����r 2��hr�rذ�P��3` + ^?���եq�`��q|`������t��|aSI!Z#�!� �T�_@%�I��qRS�*s���2y{�Ip{�pTpLpF�@�`��CRC����CCTѲ�Ipڈ�a8���b��MIN��aP1순���D<iC �C/���!uc�OP4�n �j�EVj���F��_
!uF��N����|a�֔=h?KNLA�C=2�AVSCA�@�A��R�@�4�  cSF�$�;�IrC �3�a�05��	D-Oo%g��,,m�����ޟ�:co��ǀD�6� @n���sυ�U��R�0�HANC��$LG���ɑDQ$t�ND,ɖ��AR۰N��aq0g��ѫ�X�ME��^ИY�[PS�RAg�X�A�Z�П���rEOB�F�CT��A��`�2t!S\h`0ADI��O�� y�s"y�n!��������~#C�G3t!��BM�Pmt@�Y�3�afAcES$�����W_;��BAS#XYZW�PR��*�m!��	�VQU�87  "ƀI@d���8\�pc_C:T���# ��s_L
 � 9 ����C�/�(zJ�LB�$�3�D��5��FORC�b�_A�V;�MOM*�q�SaԫBP`Ր�y�HBP��ɀE�F����AYLwOAD&$ER�t&3�2�Xrp�!��R_FD�� :� T`I�Y3��Ed�&��Ct��MS�PU
$(kpD���9 �b�;�B�	E�VId�
�!_7IDX��$����B@X�X<&�SY�5� �R_H�OPe�<��ALAR1M��2W�r����0= h�@Pnq�`yM\qJ@$PL`A&�M#�$�`��� �8�	���V�]�0æ`��CU�PM{�U��>n�TITu�
1%�![q��Z_;���? �B pQk��6�NO_HEADE ^az��}ѯ��`􂳃 ���dF�ق�t�����@�@��uCIR#TR�`��ڈL��D��CB@4�RJ��:�[Q���A�2>���OR�r��O����T`�UN_OO�Ҁ$@����T�����I��VaCnpVPDBPX�WOY���B#�$�SKADR��DBT��TRL��C���րfpbDs��~�DJ$j4 _�DQ}�։PL�qwbWA����WcD�A��A�=�2�UMMY9���10���DBd����D;[QPR��� 
,�Z���E� O�Y1$�a�$8��L)FL!/��9����0GG/.�2�PC�1Hf/_c�PENEA@Tf�I��/3#�RECOR>`"JH @ �oE$L�#F$#�PR���+jp��nq�_yD$�qPROSS]��
���R�r�` u�$T�RIG96PAU�S73ltETURN�72�MR:�U 0�Ł0EW$��`SI�GNALA�QR$L�A�З5�1G$P�D�H$Pİ�AI��0�A�C�4�C��D�O�D�2�!�6G�O_AWAY2M�OZq�Z�� CSޏ�CSCBg�K qԻa#���ERI�0�Nn�T�`$������FCBPL�@QBGAGE���P��ED|BD�wA[CD�OF�q[F0�F�oC��MPMAB0X�oC�$FRCIN��2Dk��@��$N)E�@�FDL8�� L� ����=���Rw�_��P� OV�R10���lҠ��$ESC_�`uDSBIO����pTe�.E�VIB�� `s���Z��V��pSSW���$�VL��:�L k��X���ѣ�bQ���&�USC�P��A=�	Q��MP1%e&S*`��(bt`'c5۳ESU d��-cWg&SWg?cWd�����Wd��Wd.���AUTO$�Ya҃�ac�SB����-d��&SwB�[��GB�f$VO�LT�g �� � �GAOD!�q��\�@:�ORQҀKr�a�$DH_TH�E&0�Rgp� qtnwALPHnt��o��w0! Vp]�$�.�Ra�[Ӏ�s�5�`r�CQ#BUD��S� F1M��sV
��;��Lb�tk�:��BRTHR��L���T`�Z��V0ɖ��DE  �1��2�⋅������ ��kѯ�aәTt0V� ꆸ������̈Я�-�"�N~��sS2�����INHB��ILTG0ɡ�T?��3$�w� �E��PqQxQ�TqPe�Z�0Y�AF}�O�� ����ڗ��qPڳ�ē����bPܙ���P�L?���3���TMOU��ēS���� ��s� /�S18���O�Aܙ��1I����CDIƑ˩�o�STI��գ�O`:ҋ�,0���AN���Qg�S��+r�#x!$�����w�_���&�PRA�P`vC�����MCNeQe���=��VERS��r�oPIw�FPåǲ�Ш۷G.�DN��G>�����F�2�Ƿ��M�7�F��_�MN�D̠,����d�{��a����OB���U˱z���DI���#Ā��3�����A���w�F0x���3�ON�5���Q��VAL�CR[�_SIZ��b�;Qn�REQ�Rb��]2b���CHq�΂Āڃ�Ռ�����:�n�S�_U��X��wWFLG����wU$CV��iMGP�QδFLX�P�923R�u���EA�L�P-�C	��+rT��W��� �R�c���NDMS7� �љK>S�P_M'0h�S�TWv������AL�P���Q���U���U�IAG,�o��d(�U�-�T"A-`� ���A�����H`��dQ`��6��Pq_D& ��1s��.�P�F��"2�T�� ? 7 1A>��#�#L��?_=i @@>LD�c���0n�FRI�0 ``Ѐ��1}ѲIV\10�*�^1�UP`��0a��C�LW��
`L=S&-c&&S�C.w�� L���! ����d�Q$w�҇��$w����
�P�5RSM���V0�h � r��d^2AMW�a_TRp}�8@?NS_PEA����8< ��$�SAVG�8��6G]%���CAR� �`�!�$���"CR a���$ d�#E�@��N�"STD���!Fpo��'QOF��%�f�"RC���&RC۠ �(F�2A�R#7���%, gMA�Q_�a��
Q�Q��al2��u4Ib�r7I�R�9wQ�7�R�8M/��!CpR� � �p�2F<�ScDN�a0   W�2QM P $Mi��s$cA�$C�c@m�9���4�AT��0CY_ N LS!IG1x'yB��hy@@H2Y�NO�x���SDEVI�@� O@$�RBT:VSP�3�CuT�DBY|�A	W`3C�HNDGDAP ]H@GRP�HE iXL�U��VS�Fx2�: DL1p Q6ROp���FB�\]�FEN�@��S��ChA7R d�@DOd�PMCSb�P薇P|�R��HOTSWz4:2�DMpELE�1/e8x\8`�RS T�@��`�r� hf��`OL�GCHA�Fk�Fs����C�A@T � �$MDLUb 2S@�E���q�6�q	0P�i�c�e�cJ��	u�ݢ�#~5t+w�PTO©�� �byU DSL�AVS� U  ��INP �	V�Њy�A_;�ENUAV; $R�PC_�q�2� 1bL�w���tSHO+� WA ���A�a�q�2�r��v�u�v�rCF�� X` ,f��r�OG gE��%XD�h��pC�Iߣ�i�MA��D�x AYr?�W� p�NTV	��D�VE�0@�SKIB��T�`g?Ň2��" JZs�! Cꆻ���f�_SV/ �`X�CLU��H���O�NL��'�Y�T��O=T:eHI_V,11 �APPLY��HI�4`;�U�_ML�� $VRFY8��	�U�M{IOC_�I���J 1/��߃O��@X�LSw"`@$?DUMMY4����ڑ�Cd L_TP����kC��^1CNF f���E��@T�y� 	D_#UQ_��ݥ�YPCP��=�� �������d���� Ys +�
0RT_;PިRVI�rNO�CCb Z�r�TAE���=�פ�DG��@[ D�P_B�Ae`kc�!I��_��H���u�� \�p�Ab=cARGI�!�$���`[ ~T_wSGNA] ��`U��IGN�Տ��� ��V������ANNUN��&�˳�EU�J'�ATCH���J�ƣu�u^� <@g�����:c	$Va�������QEF] I�� �_ @@FͲIT>b�	$TOTi �C��O�c�t�M�@N�I�a`tB��c�r��A>���DAY@CLOAD�D\�n�����q��EF7�XIJ�Ra��K���O%���a��ADJ_R�!@b��>�H2�"A[�
 c�%��`a͠�MPI�J��D �A8��?�Ac 0��ѐ��� ��Z�ϡ�U|i ��CTRL� �Yp d��TRA�8 ?3IDLE_PAW  �Ѡ��Q�V�G�V_���`c ��o�;Q@e� 1q$��6`<cTAC-3@��P�LQ�Z�Rz�\ A-u:ɰSW;�A\���/J��`�b�K�OH�(OP9P; �#IRO� �"gBRK��#AB � �O������� _ ���F���`d͠, j@S�oRQDW��MS��P6X�'z��IFEgCAL�� 10^tN��V��豊�V�(0L}f�CP
��N� 9Yb�0FLA_#�3OVL ��HE���"SUPPO��ޑ\B�L�p��&2X�*$Y-
Z-
W-
��`/��0GR�XZ�q6�$Y2�CO�PJ�SA�X2R��*r�!���:��"��I�0)�f{ `�@CACHE���c��0�s0LA�Z SUFFI, �C��q\���6���QMSW�g �8�KEYIMA-G#TM�@S��n�
2j�r���ROCVsIE��~�h �a�BGL����`�?�� 	Q���i��6!`STπ!�����������E�MAI�`N�����NY�FAU� �j�$"�qa��U�3���� }�k< �$I#�US�� �IT'�BUF`��D9NB���SUBu$�D�C_���J"��"SAV�%�"k������'�;��P�$�UORD���UP_u �%��8O�TT��_B`��8@LaMl�F4��C7AX@C�v���Xu 	��#_G:��
�pYN_����l6���D�E��M�����T��F���caC�DI`BEDT�)@C��~�m�rI�GD�!c�&��l`��-���P��FZP n (�pSV� )d\�ρ���A��o�� ����>"$3C_R�IK��kB��hD�{pRfgE.(ADS�P~KBP�`�IIM@�#�C�Aa�A��U�Gh���iCM! IP��0KC��� �DTH� �Sd�B*�T��CHS�3��CBSC��� ��V`�dYVSP�#[T_Drc/CONV�Grc[TH� �Fu F�ቐd�C�0j1��SC5�e]C�MER;dAFBC�MP;c@ETBc �p\FU DU�i ��+�~�CD�I%P702# �EO����qWӏ�SQ��QǀSU��MSS�1ju�D4`�T�RB`��A�1r� "�Й��4$ZO@s���l��U6�&��eP���eC�Nc�l��l�l�iGR#OU�W)��S c�MN�kNu�eNu�eNpR|b|�i�cH�pi��z
 �0CYC���s�w��c��zDEL�_D��RO�a���qVf���v{�O�2��� 1��t��:R�ua�.#�L ��AL� �1sˢ I1¡�J0�PB����"�R^�T�Gbt �,!@��5��aGI1L�cR1s 
�0ԠN	O��1u��������R�P����Cڠ	�<����DMA��J0��0vH *	�L U�1#J�Q��V
�[�7A z���z��z��z�Ѩz�Fz�7w�8w�9Pw���y���1��1��U1��1��1Ě1њU1ޚ1�2��2�����2��2��2��2�Ě2њ2ޚ2�3J��3��3����3��U3��3Ě3њ3ޚe3�4���2XTF��1w6�.(�0�f�0�U�0ŷ�e� FDR�5�xTU VE���?1���SR��REr�F���OVM~Cz)�A2�TROV2ɳDT� R�MXa�I�N2���Q�2�IND�p�r�
���0�0�0G@u1��[�G`��{�D_֎[�RIV�P��G�EAR~AIOr�K"N�0�y�p�5`�@�a�Z_MCM܀ ���F��UR��Ryǀ��!?� ��p?nЋ�?n�ER�v�!�!��P��zI:�PXq�B�RI0%�Ђ#ET�UP2_ { ����#TDPR�%T�Bp������3���BAC�2| T��"�4E)�:%	`^B��p�WIFI��� Mc����.�PT���LU=I�} � ��K UR�c!���B�18SPx E�EMP�p�2u$��S^�?x��qJق0
3VRT����0x$SHO��Lq�6 ASScP=1��PӴBG_���-�����FO�RC3"Ag�d~�)"FUY�1�2\�2�
A�h� p� |n��NAV�a��������S!"��$�VISI��#�SC�M4SE����:0E�V�O��$���M����$��I��@��FMR2��� �5`�r� @�� �2�I�9 �F�"�_���LI�MIT_1�dC_�LM������DGC�LF����DY�L	D����5������J�� ����u	 �T�FS0Ed� �P��QC�0$E#X_QhQ1i0�PԪaQ3�5��G�oQ��� ����RS�W�%ON�PX�EBcUG��'�GRBpگ@U�SBK)qO1nL� ��POY �
)��P��M��O,Xta`SM��E�"R�����`_E � y
@��TERMZ%9�c%��ORI�1_ -�c)SMepO��_ ��c&>`�`�(�c%���?�UP>� ��� -���bQ���q#� ���G�*� ELTOQ�p�0�PFIrc�1Y��P|�$�$�$UFR�$��1L0e� OTY7�PT4q�k3wNST�pPAT�q=4PTHJ�a`�EG`*C�p1ART�� !5� y2$2REyL�:)ASHFTR(1�1�8_��R�PcJ�& � $�'@��  ��s�1 @I�0��U�R G�PAYLyO�@�qDYN_k����.b�1|��'PERV��RA��H��g7�p��2�J�E-�J�RC����ASYMFL3TR�1WJ*7�����E�ӱ1�I��aU�T�pbA�5�F�5P��PlC�Q1FOR�pMF��I!���W���/&�0F0�a_C�9H��Ed� �m2N�,��5`OC1!?�$OP����c������bRE��PR.3�1a�F��3e��R�5e�X�1(�e$PWR��_����@R_�S�4��et$3�UD��N�Q72 ]���$H'�!�`�ADDR�fHL!G �2�a�a�a��R��U�w� H��SSC����e-��e���e��S�EE����HSCD���� $���P_"�_ B!rP�����DTR�HTT�P_��HU�� (��OBJ��b(�-$�fLEx3Us�� � ���ะ%_��T?#�rS�P���z�KRN�LgHIT ܇5��P���P�r���0���PL��PSS<�Ҵ�JQUERY_F�LA 1�qB_WE�BSOC���HW��1U���`6PIONCPU���Oh� �q����d���d����� �IHMI_E�D� T �RHv�?$��FAV� �d�Ł��IOLN.
� 8��R�@�$SLiR$I�NPUT_($t
`��P�� ـwSLA� ����5�1��C��B {IO6pF_AS7��$L%�}w%�A��\b.1�����T@HYķ�������h�UOP4� ` y�ґ�f�¤�������`PCC
`����#�|��QIP_ME��n��� Xy�IP�`<�U�_NET�9����Rĳs�豟D�SP(�Op=��BG�`�T���M�A���3 lp:CTAjB�pAF TI�-U��Y lޥ�0PSݦBUY IDI�rF ��P�0�a�� �y0�,����Ҥ�NQ�Y R���IRCA�i� �� ěy0�CY�`EA��������CC����R�0�A��7QDAY_���NTVA����$��5� ���SCAd@��C9L���� ��������8�Y��2e�o�N_�PCP�q��ⱶ��,�N����
�xr����:p�N� 2��Ы�(ᵁ����xr۠LABy1��Y �ǗUNIR��Ë ITY듭��eK0s�#��5���R_UR�L���$AL0 EAN��ҭ� ;�T���T_U��ABKY9_z��2DISԐ�NA��Jg����P�C$���E��g�R�D�З A�/���J����FLs��7 Ȁ�Ѿ�
�UJR� ���F{0G��E7X��J7 O R/$J8I�7��$R�d�7��E�8{�H�oAPHIQS�z��DeJ7J8Bޱ�L_KE*� o �K��LM[�� � <X�XR�l�u���WATCH�_VA��o@D�tvF'IELc��cyN��&4� o1Vx@���-�CT[�9�m�t�p�LGH���� $��LG_SIZ�t�z�2y�p�y�FD��Ix���+! ��w�\ ����v��S� ��2��p�������\ ����A�0_gCM ]3NzU
RFQ\�vv�d(u�"B��2�p�����I��+ �\ �̥v�RS���0  >�ZIPDUƣ�aSLN=��ސ�p �z6���f�>sD�P�LMCDAUiE�AFp���TuGH��RE�|�BOO�a��� C��I�IaT+���`��RE����SCR� �s��D�I��SF0�`RGIO"$D�����T("$�t|�S�s{�W$|��X��JGM^'MN3CH;�|�FN��a&1K�'uЅ)UF�(1@n�(FWD�(HL�)STP�*V�(%Г(,��(RS9HIP�+��C[T�# R��&p:'^9U=q�$9'�H%C�d���"Gw)�0PO�7��*��#W}$���)E]X��TUI�%I�� �Ï���rCO#C� N*�$S��	)���B@�NOFAN1A|��Q
�AI|�t:��EDCS��c�CT�c�BO�HO�GS����B�HS�H(IGN������!O���DD�EV<7LL��H�-��Ц(�;�T�$��2�p���=��#A���(�`�{�\Y��POS1�U2�U�3�Q���2�@�Ш ��{�PtD�����&q)��0�d��VSTӐR�YU�\@ `� �$E.fC .k�p<p=fPf	��4��� LRТ� ��x� c�p��<�Fp�d̐?"^�_ ������Kq&���cT�MC�7� ���CL�DPӐ��TRQLaI#ѽ�ytFL��,r�5s8�D�5wS��LD5ut5uORG���91HrCRESE�RV���t���t��p��c�� � 	`u95t5u��PTp���	xq�t�vRCLMC������D�q/M��k�������$DEBUGMCAS��ް��?U8$�T@��Ee�g����MFRQՔ�� � j�HRS�_RU7��a��A<��k5FREQ� ��$/@x�OVER���n��V#�P�!EFI�%�a��g�8,S���t� \R�ԁ�d�$U�P��?��p�PS�P��	�߃C��͢a��U�\�l�?( 	����ISC� Yd@�QRQ��	��3TB � Ȗ0A�՘AX����ؗ�E�XCESjҔЪ�M��\��������=����SC�P � 	H��̔_��Ƙǰ]������MKHԳ�K�J� m�B_K�F�LIC�dB�QU�IREG3MO��O�˫3��L�`MGմ �`��T����aNDU�]���>��k�G�Df��I�NAUT���RSM>�a��@N)b]3x-��p5�PSTL\�w� 4X�LOC�V�RI%��UEXɶA�NGuBu�R�ODA����������MFO����Y�b@p�e4�2k�SUP�fv��FX��IGG� � ��p�c ���cQ6�dD�%�b|� !`��!`��|��3w�ZW�a�TI��p;� M���[�� t��MD
��I�)֟@����HݰM��DIA�����W,!�wQ�1*�D�)��O���n]�� 0�CU��VP��pu��O!_V��ѻ ���S�LX�5������P��h0N���P��KES2���-$B� �����ND2����2_{TX�dXTRA�C�?�/��M�|q�`�Pv��XҰ�Pt �SBq`�USWCS��T��	���PULYS��A�NSޔ��<R��JOIN��H��~`j�=��b��b�����P=��$��b$���TA����S���hS�HS�E��SCF�b��J��R��PLQ�o ���LO�b�н.���^� ���8�������0�RR}2��� 1��zeA�q d$��IIΐ+�G�A2+�/� �PRI�N�<$R S�W0"�a/�ABC�D_J%�¡u���_J3�
�1S�Pܠe�u�P��3P��р`u��J/�(��r�qO8QIF��CSKP"z{�{�J���QL28LBҰ_AZ�r��~ELQ��OC�MPೕ�T���RT�����1�+���P�1��>@�Z�ScMG0��=�JG�`�SCL�͵SPH�_�@��%V�u� RTER`  �< A_�@G1"�A0�@c��\$DI�
"�23UDF�v}!LW�(VELq�IN�b)@� _BL �@u��$G�q�$�'�'p�%`<�� ECHZR�/�TSA_`�%���E}`<����5��Bu�H1}`_�� �)5D2d%��A4I�1�N9t&��DH�A�:��ÀP$V `�#>A$��ł�+$Q�R}ӆ���H �$BE�Lvᵆ<!_ACC�E�!c��7/��0IR�C_] ��pNT<T��S$PS�rL�d�/Es��F{�@F
��9gGCgG36B���_�Q�2�@�A����1_MGăD1D�A]"łFW�`��`�3�EC�2�HDE�K�PPABN>G��SPEE�B�Q%_pB��QY�Y��11$US�E_��,`Pk�CTEReTYP�0�q P�YN��Ae�V)�B�QM���ѷ��@O� YA�TINCo�ڱ�B��DՒ�WG֑ENC�����u�.A�2Ӕ+@INPOQ�I6Be���$NT�#�%NT2c3_�"łIcLO� ł_`��I�_�if� @_�k�? �` ej�C400fMOSI�A������A䃔�PERCH#  �c��B" �g� �c��lb=�����oUHu@�@	A6B(uLeT 	~�1eT�ljgv�fgTRK@%�AY�� "sY��q6B�u�s۰�8]��RU�MOMq�Ւ�Y�MP�^��C0�s�CJR��DUF �B�S_BCKLSH_C6B)����f���S�t�H��RR��QDCLALM-d���pm0���CHK���GLRTY���d��Y�8��)Üd_UM]�ԉ�C��A!�=PLMT� _L�0��9��E�.� ��#E)��#H� =��Q3po�xP	C�axHW�頿Eׅ�CMCE��@�GCN�_,ND�Ζ�SF�1�iVoR��g<!���0r���CATގSH)�,�DfY��f`��7A���܀PAބ&�R_P݅�s_ ��v���s����JG��T]���Y�����TORQUaP��c�yPOU��b��P%�_W�u�t��1D��3�C��3C�IK�IY�I�3F�6�����@�VC�00RQ�t��1࿾�@ӿ��ȳJRK������UpDB Ml��UpMC� DL�1BrGRVJ�Cĭ3C��3$�H_��"�j@q��COS~˱~�LN ���µ�ĭ0����� u����̓��Z���f$�MY��؊��˾>�THET0reN�K23�3hҧ3��C�Bm�CB�3C! AS� ��u��ѭ3��m��SB�3��x�GTS$=QC�������<����$DU��Kw��B�%(��%Qq_ ��a��x�{�K���b(��\�A`Չ��p�{�{�LPH~�g�Aeg�Sµ��������g������֚�V��V���0��V��V��V���V��V	�V�V%�H��������G������H��H��H	�H��H%�O��O��OTV	��O��O��O��UO��O	�O�OցFg���	�����S�PBALANCE�_-�LE��H_`�SP!1��A��A>��PFULCEl�Tl��.:1��U�TO_����T1T2��22N���29` �!�qnL�=B�3�q�TXpO�0
A4�IN�SEG�2�aREV8��`aDIF�uS9�1�8't"1�6`O!B.!t�M��w2�9`���,�LCHWARLRCBAB�� ��#��`-ФQ 5�X�qP�R��&��2�� 
p�""��1eROB͠�CR0r5�����C��1_��T � �x $WEIGH�P`$��?3à�I�Qg`IFYQ�@LAG�Rq�S�R �R7BILx5OD�p�`&V2ST�0V2P!t�BW0��01�&1/0�30�
�P�2�QA  2yřd[6DEBUg3�L_@�2�MMY�9&E Nz�D`3$D_A�a$�0���O�  �D�O_@A.1� <@B0�6�m�Q�B�2��0N-cdH_p`�P��2O�� ��� %��T`"a��Tx/!�4)@TICKh3| T11@%�C ��@!N͠�XC͠R?��Q��"�E�"�E8@PRO�MP�SE~� $IR��Q��R;pZRMAI)��Q�R4U_r02S; �q�P�R8�COD�3FU�Pd6ID_[�vU �R!G_SUFF�u� l3�Q;Q�BDO�G �E�0�FGRr3�"�T�C�T�"��U�"�Uׁ�T8D�0ǺB0Hb _FI�1�9*cORD�1 50�236V�+b�Q1@�$ZDT}U����1;E�4 *:!L_NAmA�@�b>�EDEF_I�h�b �F�d�E�2�F�4�F�c�E�e�FISP��PAKp�Ds�C�d��44בi��2D�"�It��3D�O#OBLOCKEz��S�O�O�Gq�R�PUM�U�b�T �c�T�e�T!r�R�s�U �c�T�d�R�6�q�S � ���U�b�U�c�S�Z��X�@P` t�@qDe�)@W�x���s����TE�<D�(� l1LOMB_t��ɇ0V2VIS;�WITYV2A��O�3A_FRI��a #SIq�QR�@���@�3�3V2W��W��4����_e��QEAS^3�Rϡ��_�[pT:R�4�5�6_3�ORMULA_I�z���THR^2���Gtg�30f��<8��5COEFF_O �A	 ��A��GR�^3Sg0BCAnO/Ca$��]3n�1GRP�� � � $h�p�YBX�@TM~w����u�B�s��bCER�, Tttsd$`�  ��LL�TSpS~�_�SVNt�ߐ��$`ʸ��$`� ��SwETUsMEA*P��P��W0�1+b/0� g� h��  @�ڐo�l�o�cqz��bH�@cqq`tP�G��R�� Q\p*q[p��t>�c NPREC>azt�5@MSK_$�|�� PB11_USER����{ 8���VEL����{ 0�$Ō!I]`���MT�ACFG���O  �@@ O�"NORE-0l@o�V��SI.1�d��6�"UaXK�fP!��DE��� $KEY_��3�$JOG�� SV������!��}�SW�"�a\aS�ՐT|�GI�!0| ~^�� 4 h�8�'d2�!XYZc����3�  �_ERR#�� 8Ԡ�AfP�V�d��1����$BUF��X�����wMOR|�� HB0CUd�lA�!��GQ\axB�,"!a$� r���a����_��?�G~�� � �$SIՐ���VOx��T� OBJE_���ADJU)B��EGLAY���%�DR�OU.`=ղВQ0b=��T���0���;BDIR���; I�"0DYNW�2��	T��"R���@�0�"�OPWORK����,%@SYSB9Uy�SOP��$ޑ�U�; P�pN�<�PA�t�>�"��+OP�PUd!0�`!z��l�IMAGw�1B0y�2IM�Õ��INe�d��RGO�VRD��-��o�P q��0��J�Os���"�L�pBa���o�PMGC_Ee`���1Ny �M A�21�2  ����SL_��� �� $OVSL �ǫ�?q�`��2�" -�_��k�P��k�P u���2�C� �`��Ź���_ZERr�D��$G��� 2=���� �@*���%O~PRI��� 
JP8+�S�=!/�L��ح�T�� �0ATUS��T�RC_T���sB ��}fs�9s�1Re`��� DFAm����L���"��0a� ޱ��XEw{����1�C0vUP��+p�	qPXP�j�43� � �PG\��>�$SUBe�%��qe9JMPWAcIT z}%LO��yF�A�RCVFBQ��@x"�!R�� �x"A�CC� R&�B�'I�GNR_PL9D�BTB�0Pqy!B�WbP�$w�Uy@�%I�GT�PI��TNL�N�&2R��rL�N<P��PEED \HADOW�06�w���E[q4jO!�`S�PDV!� LbA�z�`�07�3UNI�r��0"!R��L�YZ`� o��PH�_PK��e�RETRIE9{�q�����0'PFI"�� �xG`�0D 2�g��DBGLV�#LO�GSIZ��EqKT��!U��VDD�#$0_)T�G�MՐCݱ���|@eMRvC}�3�CH�ECK0��	�P�O�V!�k�I��LYE(!��PArpT�2�K�W��@P2V!� h $ARIB iR� c�a/�O�P8�ӐATT��2�IF`|@z�Aq4S�3UX�����PLI2V!�� $g���ITCH�x"[�W �AS9���vTLLBV!��� $BA�DYs��BAM!���Y9�PJ5��Q��R�6�V�Q_KNOWh�Cb��U��AD�X�V��0D�+iPAYGLOAt��Ic_��(Rg�RgZOcL�q���PLCL_�� !7��b�QB��d���fF�iC֠�js��d�I�hRؠ�g�Ғ�dB����J��q_�J�a#���AND���Ĳ.t�b�aS�r�P�L0AL_ �@�P�0���QրC��uDNcE���J3Cp�Wv� TPPDC�K�����ĳ�_AL3PHgs�sBE���gy|��K�1�� �� ���HoD_�1Oj2ydD��AR��*��;�&���TI�A4U�5U�6��MOM��a���n���{�Y�B� ADa���n�\��{�PUB��R�� ҅n�҅{���2�Wp�ѾW �  PMsbT� �BxQ����� e$PI ��81��TgJ��ni*J�IV�Id�Ir�� [��3!��>!��rp�Ӫ�U3HIG�S U3�%�4얎4�%� ����"����!
��!�%SAMP���^��_�8�%�P4s ю� ��[ 	ӝ�3 ���0� ��&�C�����^��Sp2��H&0	�IN�Sp B����뤕"��6���6�V�GAMM�SyI�� ETْ��;��D�tA�
$ZpIB�R!62IT�$HIBِ_���C�˶E��bظAҾ���LWͽ �
���7���rЖ,0:�qC�%CHK��"o �~I_A� ����Rr�Rqܥ�Ǚ���ԥ���Ws �$�x 1���I�7RCH_DAƺ RN{��#�LE@��ǒ!,��x���90�MSWFL�$�S;CR((100��R@��3]B��ç��a���x�َ0��PI3A9�METHO����%V��AXH�XX0�԰62ERI��^�3���R�0$u	��pFH{�_���?ⲣ1��L�L�_�a�OOP࣡��wᲡ��APP:���F���@{���&أRT�V�OBp�0�T����;��� 1��I��� ��r���RAv�@MGA1AS�T�SV-��P�CsURg�;�GRO[0S_SA�Q��Y�#NO�pC!"�t Y��Zolox�����`��!b����&�DO�1A���A����Х��A����A"�WS�c ��Bh�*�� � ���YLH�qܧ���SrZ�]B�o��=�q�õq_�C�1��M_W���g���c�M� �`Vq�$p�x1o�3"r�PMJ�,�� �'Aȡ 9�!Wi:�$�LWQ|ai�tg�t@g�tg{t� �N`P���S��SpX�0O�s�RqZ��P� *�� ���M���������������X��� ��5L:�q_~R� |�q#( Y����&n��&{�Y�Z� �'�&t��Q��qQ#��"J0��qP}`�$PQ��PMON_QU�c� � 8�@Q�COU��%PQTH��HO�^0HYSf:PES�R^0UEI0tO��@O|T�  �0�PGõz�RUN_+TO��POْ.�'� PE`�5C��A�<�INDE�ROGGRAnP� 2g��NE_NO�4�5I�T��0�0INFO�1� �Q�:A�uȉ2IB� (��SLEQݖFAѕF@��6eOSy�T�{ 4�@ENAB�>�0PTION.S%0ERVE���G��A0�zCGCF�A� @bR0J$Rq�2����R�H�O�G "�EwDIT�1� �vR�K�ޓʱE�sNU0W*XAUTu�-UCOPY�ِN\����MѱNXP\[qƯPRUT9� _RN��@OUC�$G��2�T���$$CL<`?0����Q��M�� �P�S�@��X�PXK�QIRTU��_�P�A� _WRK 2� e�@ ?0  �5�QMorYhJo|m |lA	�`�m�o��`��o�o�f�e�l}�a`I[ct'`BS��*� 1�Y� <7��� ����&�8�J�\� n���������ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T�f�x����� ����ү�����,� >�P�b�t���������vsrCC��LMT?0v���s  dѴ�INڿ�дPRE/_EXE��)����0jP��za'`DVʽ�S�@e)�%�select_macro����k�|��qtIOCNVVB��� ��P��US�ňw���0V 1.4kP $$p��a�|�`?���߰>� P�b�t߆ߘߪ߼��� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������� ��$�ѰLARM�RECOV �^�����LMDG� �Ь�LM_IF ���d  YST-�323 Coll�aborativ�e speed �limit (T�CP) led �it.(L:6) ������)�;�M�_��q��, 
 ����#�>TELE�OP ǘLINE� 6ǑAUTO �PA��DǙJOI�NT 100 %�����$���1��@�$�@��C�TL-003 s�ystem is� in erro�r status� 0  clea�r뀪���ί��NG�TOL  @� 	 A\���Ѱ�PPINFO �� f�L�^�p����  ������ k���ۿſ�����5���Y�C�iϏ�%��� ٯ����������'߀9�K�]�o߁ߓߙ�P�PLICATIO�N ?t���|�Ha�ndlingTo�olǖ 
V9.40P/17\�
88340�����F0�	�549���������7DF�5�О�ǓNone���FRA�� �ؒ��,�_ACoTIVE1�  ��� �  ��ސMO�D��������CH�GAPONL�� ��OUPLEDw 1	��� >��B�T�f���CURE�Q 1
��  T*p�p�p�	���� ����l��������������i3l��p���^�H��A�t
HTTHKY�FXv| ��*<N` �������� //&/8/J/\/�/�/ �/�/�/�/�/�/�/? "?4?F?X?�?|?�?�? �?�?�?�?�?OO0O BOTO�OxO�O�O�O�O �O�O�O__,_>_P_ �_t_�_�_�_�_�_�_ �_oo(o:oLo�opo �o�o�o�o�o�o�o  $6H�l~� ������� � 2�D���h�z������� ԏ���
��.�@� ��d�v������������TO�����DO_CLEAN���E��NM  �� p�������ɯۯv�DSPDRYRL�&��HI��o�@��G� Y�k�}�������ſ׿�����ϻ�MAX@��,�����=�X,���9����PLUG�G,�-�9���PRC*��Bm�q�6�(���O����SEGF�K���� �m���G�Y�k�}ߏ�����LAP$�7ޡ����� �+�=�O�a�s������� �TOTAL�_ƈ� �USENU
$�1� �������RGDISPMM�C�d�C�O�@I@�1�O"�D���-�_STRING� 1��
�kM��S��
��_ITEM1��  n���������  $6HZl~���������I/O SIG�NAL��Tr�yout Mod�e��InpNS�imulatedޡ�Out`�OVERR!� =� 100��In� cyclT���Prog Abo�rj��JSta�tus��	Hea�rtbeat��MH Faul��Aler�!/ !/3/E/W/i/{/�/�/�/ (���(��� �/??&?8?J?\?n? �?�?�?�?�?�?�?�?�O"O4OFO�/WOR И�~A�/XO�O�O�O �O�O __$_6_H_Z_ l_~_�_�_�_�_�_�_�^PO���"`�K oEoWoio{o�o�o�o �o�o�o�o/A�Sew��bDEV%n�p9o���� #�5�G�Y�k�}����� ��ŏ׏�����1�>C�PALT�-j� �OD�������ȟڟ� ���"�4�F�X�j�|��������į֯X�GRIB�������6�H� Z�l�~�������ƿؿ ���� �2�D�V�h�z�����R�-��&��� �������"�4�F�X� j�|ߎߠ߲�������������PREG n�W���0�~���� ��������� �2�D� V�h�z���������$��$ARG_~@D ?	�����  �	$$	[�]�$:	��S�BN_CONFIQG�XWq�RCII_SAVE  $zm���TCELLSET�UP 
%  OME_IO$�$%MOV_H8� ��REP��#���UTOBACK� 	tF�RA:\D� X.D�z '`�D��w� �s  �25/11�/29 20:2/6:16D�;D�`��#//h��C/�j/|/�/�/�/�/D� X/�/??(?:?L?�/ p?�?�?�?�?�?�?g?  OO$O6OHOZO�?~O��O�O�O�O�O�O����  c_F_\A�TBCKCTL.TM�)_;_M___q_.8INIm��j�~CMESSAG�� �Qz �[ODE�_D� �j�XOx�p�_@PAUS6`� !� , �	�9/Do��,		2afotgZo �o~o�o�o�o�o�o �oH2lzyd`?TSK  mwxz�9UPDT�P�Wd�p�VXWZD_ENB�Tf
�v�STA�U�u��X�ISX UNT 2��vwy � 	 �v�uu�h�V��� ���a<D�R����P -��3�����9m������R��n�t�<���MCP� �s��ŀ�����!���4�M[ET��2@��y �PQ�A�J�A�@�A�ܸB�FiA�!)BS����>�01>��,�>��"?�]w�?-��?���N5�SCRD�CFG 1]Y ��� ���%�7�I�pD�Q��ݟ������Я� ��[���<�N�`�r��������7���FGR`9��p�_ԳPNA� �	FѶ_E�D�P1��� 
� �%-PED�T��H��R�v����Es� -FE�D��;3o�>���  ����2�����B�  ����{�����j�����3��#� �G�Y���@G�ߠ�6�����4�W������Zݨ�� Z�l������5K��� ���Y�t���&�8���\���6��d��Yހ@����(��7 �S0wY�w��f���8����{�IZ��C/��2/����9{/��//L Zݤ/?V/h/�/�/��CR���?�?Tn?��? ?2?�?V?԰!�N�O_DEL�ҲGE_UNUSE޿�дIGALLOW� 1�   �(*SYST�EM*��	$S?ERV_GR[�@n`REG�E$�C���@NUM�J�C�M�PMU?@���LAYK����PMPAL�PUCOYC10 N3^P<!^YSULSU_�M�5Ra�CLo_�TB�OXORI�ECU�R_�P�MPMC�NVV�P10|I^�PT4DLI�p��_�I	*PROG�RA�DPG_cMI!^Ko]`AL+e�joTe]`B�o�N�$FLUI_RE�SU9W�o�O�o�dMR�N�@�<�?�; M_q����� ����%�7�I�[� m��������Ǐُ돀���!�3�E�W�2BL�AL_OUT ��K���WD_A�BOR:PcO��IT�R_RTN  ��$�빸�NONS�TO�� lHC�CFS_UTIL� �̷CC_�AUXAXIS ;3$� h}�j��|�����ƽCE_R�IA_I`@��נ��FCFGG $�/�#��o_LIM�B2+�w �� � 	��SB\���$� 
Ԡ���)�Z���/�ĺ���[����� ����!�����L��(
�5�����PA�`GoP 1H���@��A�S�e�w�6�C�C� C7��J��]��p������� �C����������������é�̩�ժ��ߩ������2��;���PCk����U����������������ɱ����������� D� �D!�!�!��!� ��&?��H=E@ONFIpnC�G_P�P1H� +EH��ߟ߱�����������C�KP7AUS�Q1H�ף IR�S�H�A�� e����������� ���E�+�i�{�a���DA?Iץ�Mؐ�NFO 1��� �3��$�4����EA�m�m�2&�����K�wC�}��* D/q�� Ce���3��´J\��O� � ��L_LECT_�!�����EN+`�ʒܮ��NDE�#��/�1234567890@�"�A��/ҵHw��#)j��<i{� �;��/��/`/ +/=/O/�/s/�/�/�/ �/�/�/8???'?�? K?]?o?�?�?�?�?O��?��$� |��IO &��"S▒O�O�O�O�`GTR�2'DM(`��^�?�NN�(oMx Z��_MOR)q3)H��7ىU3��Y �_�_�_�_�_�[bR�*kQ*H�,S�?<�<щ�<cz�KFd���P,��;ϒo�o��o˿�o�oœh�U�Y@E�oS ߀sja�PD�B.���4cpmidbg3���&�s:��>uqpz���v  ��>x��}.��}�`�6�|�<�mgP���t��~f������@ud1:�?��~XqDEF -���zC)*�cO�buf.txtJ��|K��[`�/DM��>c���R�A��MCiR20_{RCd���hS�21����G���C�zA�d4�EI�j�A��	C-]��G/X"B�e;�F]�H�j��Df�F�%�J��iE�qu�I؂�Lڒ�YG�UI�!�oN��mID��MSo����=�c�j��f23DL�D�	>z�!� 2���}��yc
�@�x9� C��e D�4G�E��� � E%q�F�֟ E�p�u�F��P E��fF�3H ��G�M����?5�>��33��?�xnt9�q@�Q5�����RpA?aեL��<#�QU�@,�C�ϒ���RSMOFST +i����P_T1Ɠ4DM�A =ք�MODEg 5dm�@��	Q,�i;��%���?���<�M�>��Ͷ�TES�Tc�2i�`�R�6(�O�K�CN�AB����n� 8��\�n�C6dB���Cpp�s����p:d�QS ��� ����T��4�I7>����>B8m5$�RT�_c�PROG �%j%��d�1�h@N�USER��x�KE�Y_TBL  �e�����	
��� !"#$�%&'()*+,�-./(:;<=�>?@ABCc�G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~����������������������������������������������������������������������������>��͓���������������������������������耇����������������������4A8�LC�K��F�y��STA�T��2�X�_AL�M�����_AUT/O_DO�E��FDR 3:i�2�h&q[~�� �BUOSYS�T-322 Au�to statu�s check �time out� ���i�$T�ELEO8�i�� ��)qA����@Ĭ������?�ڛM�sB�õ�?�*?��?M�f=�o�T�R��-���D�.�B���C?���B�N�*po�4�N4�J5Hj5H��>��i�BJ�d�BF��pZ��[~�bbt�����5/�M*F��B�GA+$����@R���J�}BQ��H����������2>���@�@����&�CBx�HCKH<B��6>Tbt��/��u�US�H?Z?l?i�$7?�?:�� mϸ?�? p���?�?OO�?,O fOxO�M6?�O�O�O~? �O	_�?*_$_BOD_6_ p_~_T_�_�_�_�_�O o)o;o�OLoqo_�o �o�_�o�o�o�o�o�o FXo��No ���o���� @�N�$�b�x�����n ������A��b� \�z�|�n�������ʟ ���(�֏O�a�s�� ����T�ʯį��֯ ����2�H�~���>� ��ɿۿ���ϼ�2� ,�J�L�>�xφ�\Ϛ� �����Ϧ��1�C�� T�y�$Ϛߔ߲ϴߦ� ��������N�`�� ����V߼����� �����H�V�,�j� ������v����� $I��jd���v �����0�� Wi{&��\� ����/&/�:/ P/�/�/F�/�/�/� �/?�:?4?R/T?F? �?�?d?�?�?�? O�/ 'O9OKO�/\O�O,?�O �O�?�O�O�O�O�O
_  _V_h_O�_�_�_^O �_�_�O
oo"_$oo Po^o4oro�o�o�o~_ �o	�_,Q�_r l�o�~���� �&�8��o_�q���. ����dڏԏ���  �.��B�X�����N� ǟٟ럖���!�̏B� <�Z�\�N�����l��� �������/�A�S��� d���4�����¯Ŀ�� ���Կ�(�^�p�� �ϩϻ�f����Ϝ�� �*�,��X�f�<�z� �����߆����#��� 4�Y��z�t�ߔ�� ���������.�@��� g�y���6����l��� ��������(6J `��V������ )��JDbdV ��t���/� 7/I/[/l/�/<�/ �/��/�/�/?�/? 0?f?x?&/�?�?�?n/ �?�?�/OO2?4O&O `OnODO�O�O�O�O�? __+_�?<_a_O�_ |_�O�_�_�_�_�_�_  o6oHo�Ooo�o�o>_ �o�ot_�o�oo�o 0>Rh��^o ����o�1��oR� L�jl�^�����|��� Џ���?�Q�c�� t���D�����ҏԟƟ  ���"�8�n���.� ����˯v�ܯ���"� �:�<�.�h�v�L��� ��ֿ迖��!�3�ޯ D�i���τϢ��ϖ� ���ϴ����>�P��� w߉ߛ�FϬ���|��� ��
����8�F��Z� p���f�������� �9���Z�T�r�t�f� ���������� �� GYk�|�L�� ������* @v�6���~ �	/�*/$/BD/6/ p/~/T/�/�/�/�/� ?)?;?�L?q?/�? �?�/�?�?�?�?�?�? OFOXO?O�O�ON? �O�O�?�O�OO__ @_N_$_b_x_�_�_nO �_�_o�OoAo�Obo \oz_|ono�o�o�o�o �o(�_Oaso ��To���o�� ���2�H�~���> ��ɏۏ����2� ,�J�L�>�x���\��� ��������1�C�� T�y�$����������� ��į��N�`�� ������V���ῌ�� �����H�V�,�j� �϶���v����߾� $�I���j�d߂τ�v� �߾ߔ������0��� W�i�{�&ߌ��\��� ���������&���:� P�����F�������� ����:4R�TF ��d��� �� '9K��\�,� �������
/  /V/h/�/�/�/^ �/�/�
??"/$?? P?^?4?r?�?�?�?~/ �?	OO�/,OQO�/rO lO�?�O~O�O�O�O�O �O&_8_�?__q_�_.O �_�_dO�_�_�O�_�_� o.ooBoXo�otc��$CR_FDR_�CFG ;re��Q
UGD1:�W�P�aJ�d�  �`�\�bHI�ST 3<rf  ��`  ?��R@tAtB��bC�P7pD�tEtItg�P�potw�_��bI�NDT_EN6p~�T�q��bT1_DO  1�U�u�sT2��w�VAR 2=�g�p hq  �ʈ�ʈ4�R��4����m[�z�RZ�`STOP���rTRL_DEL�ETNp�t ��_�SCREEN �re�rkcs�c�rUw�MMEN�U 1>��  <�\%�_��T ��R��S/�U���e� w�ğ������џ�	� B��+�x�O�a����� ������ͯ߯,��� b�9�K�q�������� ��ɿ����%�^�5� Gϔ�k�}��ϡϳ��� �����H��1�~�U� gߍ��ߝ߯������� 2�	��A�z�Q�c�� ����������.�� �d�;�M���q�������������YӃ_M�ANUAL{��rZCD�a?�y�rG� ���R�fx"
�"
?|(��P�dTGRP 2@:�y�B� � �s��� �$DwBCO�pRIG����v�G_ERRL�OG A��Q��I[m �N_UMLIM�s���u
�PXWOR/K 1B�8����//�}DBT;B_�� C%����S"� �aDB__AWAY��Q�GCP �r=���m"_AL�F�_�Yz����p�vk � 1D� , 
��/"�/%?/(c_M�pqw,@�=5�ONTIM���f�t�_6�)
�0~�'MOTNENFp�F�;RECORDw 2J� �-?�SG�O��1�?" x"!O3OEOWO�8_O�O �?�OO�O�O�O�O�O (_�OL_�Op_�_�_�_ A_�_9_�_]_o$o6o Ho�_lo�_�o�_�o�o �o�oYo}o2�oV hz��o��C �
��.��R��K� �������Џ?��ߏ �*�����+�b�t�� ������Ο=�O��� ��:�%���p�ߟ񟦯 ��O�ǯ�]������ H�Z���������#��5����ϩ�i"TO�LERENCv$B�ȿ"� L��� C�SS_CCSCB� 2K�\0" ?"{ϰϟ���7�� 
����@�R�d�3߈���"�x�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C�Ugy��� �������R�LL]�La�m1T#2� C�C�p�F�^ A�C�%pC���#�0�? 	 A����B���?�  ��$����\0����0��B��`#sߠK/]/o/�ϓ/��/�/s/�/�/�K2�i2L�٧���L�;b�x��?�UȦ��/�Q�/`?;�@���O?�?�?�?Ȏ0A0F��?{F�A OO��7�1���9M	AB 
AZOdBAE�9$O�O�O��Oi:P��`�@0��DJCA� @5��
X-.
[$h=�� M?�>O�ڴ �q_�_�_�_:W�A<o:[<ǲ/o�/�_+oPobotoǦeACHC�V�WB$�Dz�cD�`�a=/��o�oo�oW�a.+!��2=t,y�J?� .s�s�js�w�yj� ������Q�Qs�@`��$�����A ����Bމ�o��'� 9��_]�o�N���r��� ɟ۟_�B�ʄ���YZ>`6�B��]�AΝ��c��������Z�l�~����`_м¯���
� ��̯9�,�]�o��� � H�����ٿ뿊��ƿ 3�E�W�iϬ���$ϱ� ���� Ϟ����/�A� S߶�w�V�h߭ߌ��S���ߐ�_�f	� �H�?�Q�~�u��� ����������D� �-�g�q��������� ����
@7I�cm��߾�  �����)M @qdv���� ���//I/P�m/ �v/�/�/�/�/�/�/ �/?3?*?<?i?`?r? �?^/�?�?�?�?�?O /O&O8OJO\O�O�O�O�O�O�O�O�g	 [ Q�P�su �PC4p�*p�p6U6P\�C9p/p�� �]V^PM]�6P�:P�X>P�VJ_�^P�bPa�fP�Vr]v���p Q
k���_oo�i1d1Q&oNo ;o_�co�oˏUUA   x�o�k1Q@�  �o��k�b����B��p �� 1��6�1�1C���C�cPf�L��?#�c>��{���`�cP�@a@�d��r�`B�cP�>�s�qC��p�����b�t<�o?��PH�)S�B��tq�q�p�r�`B!���eIC�&�Q��4( �oz�UU5:���AΜQ�c���򊽻��4�Q�-RB�t���������2B���-�b��`ځ`  ?�p���U�[?���}t��$����$DCSS_CLLB2 2M��p�P�^?��NSTCY 2N����  �������ʟ؟ ���� �2�D�Z�h� z�������¯ԯ��S�A�DEVICE K2O��!�$�� 4&V�h�������˿¿ Կ���
�7�.�[�R� ϑϣϵ�����4(A��HNDGD P̅�*�Cz�A�LS 2Q��_�Q�c߀u߇ߙ߽߫���?�PARAM RP���1�`�&�RBT �2T�� 8�P<C�'pÀ�pi�2l��s@"�R��(q�I�X��0�pB C7W  ��B\x�N�0�`Z����%��)���X�j��p����zq������B �(s,� F�p�V��q���b�,��B ��4&c �S� e�l�4+����H1�~����D�C�$Z��b����A,� 4�u@��X@��^@w����]B���B��cP%��C4��C3:^C4Ս�nЬ ��p8��-B{B���A���� l���C�C3��JC4jC3���yn+�3 D�ff 2�A PB W4+@:�]o� W�����/� /P/'/9/K/]/o/�/ �/�/�/?�/�/�/? #?5?�?Y?k?�?�?�o �?�?O�?6O!OZOlO WO�O�Es�?�?�?�O �O_�O�OL_#_5_G_ Y_k_}_�_�_�_ o�_ �_�_oo1o~oUogo �o�o�o�o�owO  D/Aze��� �O�o�o
��o��R� )�;���_�q������� ���ݏ�<��%�r� I�[�m��������ǟ ٟ&�8��\�G���k� ������گů���� �F��/�A�S�e�w� Ŀ������ѿ���� �+�x�O�aϮυϗ� �ϻ�����,���b� t�ﯘ߃߼ߧ����� ����:��C�U߂� Y�k��������� ��6���l�C�U�g� y����������� �� 	-?Q��� ����@+ dvQ����� ���*///%/r/ I/[/�//�/�/�/�/ �/&?�/?\?3?E?�? i?{?�?�?U�?�?"O 4OOXOCO|OgO�O{ ��?�O�?�O�O0__ _f_=_O_a_s_�_�_ �_�_�_o�_oo'o 9oKo�ooo�o�o�o�o �o�O:%^I�������H�$�DCSS_SLA�VE U��}�	���z?_4D  	���AR_MENU V	� �j�|�������ď�BY�� ���~?�SHOW 2}W	� � �b �aG�Q�X�v�������@��П֏���� @� :�d�a�s��������� �߯��*�$�N�K� ]�o�������̯ɿۿ ���8�5�G�Y�k� }Ϗ϶����������� "��1�C�U�g�yߠ� �߯��������	�� -�?�Q�c��s��� ����������)�;� M�t������������ ����%7Ip� m��������� �!3ZWi� ��J����/ /DA/S/e/��/� �/�/�/�/�/?./+? =?O?v/p?�/�?�?�? �?�?�??O'O9O`? ZO�?�O�O�O�O�O�O O�O_#_JOD_nOk_ }_�_�_�_�_�O�_�_ o4_.oX_Uogoyo�o �o�o�_�o�o�oo Bo?Qcu���o�:���CFG �X)�3�3q�5p�FRA:�\!�L+�%04d�.CSV|	p}�� �qA g�CHo�zv�	����
3q�����́܏�� ���4��JP�(���qp1� ��RC_OUT -Y��C���_C_FSI ?�i�  .�������͟���� �>�9�K�]������� ��ίɯۯ���#� 5�^�Y�k�}������� ſ�����6�1�C� U�~�yϋϝ������� ���	��-�V�Q�c� uߞߙ߽߫������� �.�)�;�M�v�q�� ����������� %�N�I�[�m������� ����������&!3 Eni{���� ���FAS e������� �//+/=/f/a/s/ �/�/�/�/�/�/�/? ?>?9?K?]?�?�?�? �?�?�?�?�?OO#O 5O^OYOkO}O�O�O�O �O�O�O�O_6_1_C_ U_~_y_�_�_�_�_�_ �_o	oo-oVoQoco uo�o�o�o�o�o�o�o .);Mvq� �������� %�N�I�[�m������� ��ޏُ���&�!�3� E�n�i�{�������ß ՟������F�A�S� e���������֯ѯ� ����+�=�f�a�s� ��������Ϳ���� �>�9�K�]φρϓ� ������������#� 5�^�Y�k�}ߦߡ߳� ���������6�1�C� U�~�y��������� ���	��-�V�Q�c� u��������������� .);Mvq� ����� %NI[m��� �����&/!/3/ E/n/i/{/�/�/�/�/��/�/�/3�$DC�S_C_FSO �?���71� P  ??T?}?x?�?�?�? �?�?�?OOO,OUO PObOtO�O�O�O�O�O �O�O_-_(_:_L_u_ p_�_�_�_�_�_�_o  oo$oMoHoZolo�o �o�o�o�o�o�o�o%  2Dmhz�� �����
��E� @�R�d���������Տ Џ����*�<�e� `�r���������̟�� ���=�8�J�\��������?C_RPI4>F?��������3?�&�o����� >SLү@d������ %�7�`�[�m�Ϩϣ� �����������8�3� E�W߀�{ߍߟ����� �������/�X�S� e�w��������� ���0�+�=�O�x�s� ������������ 'PK]o�� ������(# 5Gpk}��� ��Q���/6/1/C/ U/~/y/�/�/�/�/�/ �/?	??-?V?Q?c? u?�?�?�?�?�?�?�? O.O)O;OMOvOqO�O �O�O�O�O�O___ %_N_I_[_m_�_�_�_ �_�_�_�_�_&o!o3o Eonoio{o�o�o�o�o �o�o�oFAS e������>��NOCODE }ZU��?��PRE_CHK �\U��pA �p�< ��p�U�]�o�U� 	 < Q��������ۏ�Ǐ �#����Y�k�E��� ��{�şן��ß�� ��C�U�/�y�����s� ��ӯm���	���?� �+�u���a������� ɿ�Ϳ߿)�;��_� q�K�}ϧϝ������� ����%����[�m�G� �ߣ�}߯��߳���� !���E�W�1�c��g� y������������� A�S�-�w���c����� ��������+= asM_���� ��'�]o 	������ /#/�G/Y/3/e/�/ i/{/�/�/�/�/?�/ ?C?9Ky?�?%?�? �?�?�?�?	O�?-O?O OKOuOOOaO�O�O�O �O�O�O�O)_____ q_K_�_�_a?�_�_�_ �_o%o�_Io[o5oGo �o�o}o�o�o�o�o �o�oEW1{�g ���_����/� A��M�w�Q�c����� �����Ϗ�+��� a�s�M���������ߟ ���'���3�]�7� I������ɯۯ��� ����G�Y�3�}��� i���ſ�������� 1�C���+�yϋ�eϯ� �ϛ���������-�?� �c�u�Oߙ߫߅ߗ� �������)��M�_� U�G���A������ �������I�[�5�� ��k����������� ��3EQ{q�� ��]����/ AewQ��� ����/+//7/ a/;/M/�/�/�/�/�/ ��/?'??K?]?7? �?�?m??�?�?�?�? O�?5OGO!O3O}O�O iO�O�O�O�O�O�/�O 1_C_�Og_y_S_�_�_ �_�_�_�_�_o-oo 9oco=oOo�o�o�o�o �o�o�o__M_ �ok�o���� ����I�#�5�� ��k���Ǐ��ӏ��׏ �3�E��i�{�5c� ��ß�����ӟ�/� 	��e�w�Q������� ѯ㯽�ϯ�+��O� a�;��������Ϳ߿ y����!�K�%�7� �ϓ�mϷ��ϣ����� ����5�G�!�k�}�W� �߳ߩ������ߕ�� 1���g�y�S��� ���������-�� Q�c�=�o���s����� ��������M_ 9��o���� �7I#m Yk������ !/3/)/i/{//�/ �/�/�/�/�/�/?/? 	?S?e???q?�?u?�? �?�?�?OO�?%OOO E/W/�O�O1O�O�O�O �O__�O9_K_%_W_ �_[_m_�_�_�_�_�_ �_o5oo!oko}oWo �o�omO�o�o�o�o 1UgAS�� ����	���� Q�c�=�����s���Ϗ �o������;�M�'� Y���]�o���˟��� �۟�7��#�m�� Y������������ !�3�ͯ?�i�C�U��� ����տ������� 	�S�e�?ωϛ�uϧ���ϫϽ�������$DCS_SGN� ]	�E��-����30-�NOV-25 2�1:20 ��{29R�0:27_��x�x� [}�t��q�т�xҚ����JѨ�EƼÿ�� ��ǖ� � 1�HOW ^�	� �x�/�VERSIO�N =�V�4.5.2��EF�LOGIC 1_~���  	������C��R�%�PR�OG_ENB  ���:�{�s�UL�SE  X���%�_ACCLIM^�����d��WRSTJNT��vE��-�EMO|��zя�$���INIT� `2����O�PT_SL ?	�	�	�
 	Rg575��]�74b��6c�7c�50��1����C���@�TO�  L��� �V.�DEX��dE�x��PATH A=�A\k}���HCP_CLN�TID ?�:�� D�ռ��I�AG_GRP 2�e	�����z�	 @�  �
ff?aG�x��B�  2Ě�/�8[I@c��ς!�7@��z�@^�@
��!��mp2�m15 8901?234567�����  ?����?�=q?���
?޸R?��Q�?��?������(�?��z���x�@�  A_�Ap !7�A�88_�B4��� ��L�x�
��@�@���\@~�R@xQ��@q�@j��H@c�
@\���@U�@Mp��//'$�; ��O)H��@Ct >�d 9��@4�/�\)@)� #t ?{@��/�/�/�/�/P'?����?���_ ?}�p�?u?n�{?s ?\�Q�? ?2?D?V?h8_�
=?����0�w5�z�H?p��h��?^�R��?�?�?�?�?h8��*t0���@�?��0�;@&O8O JO\OnOP'�$_�_ Y_k_�O?_�_�_�_�_ �_s_�_�_1oCo!ogo yoo�o��Bj"� �2x{1�@"?���f�t0�d"5!�
u4V��u"�BP3t�A>u��?@[q���@`,=q��=b��=�E1�>�J�>�n��>��H"<�o� �z�s�q��� �x�C�@<(�]Uz� 4�� Z����A@x�?* �o��m*�P�b���t n���2���Ώ����ޮi>J��&�byN2�"��G�N�R�o@�@v���0��^��@ffr!l Ο�33���(���"C�� ƒI��CH�)C.?dBت"8"����'���"~�A�?�&"K����pf�B��@�p�������p�����oO3�2x>Zq3bQ@�ǡå��� 1�oAD�/  � CeR�> ������0���N�T�����3���o#����� ȿ���׿����?,��<�o��CT_C�ONFIG f���|�e�gY��STBF_TTS��
�������}���1�MAU�������MSW_C5F��g�  # �ڿOCVIEW��h!�-���s߅� �ߩ߻��ߟ�a���� �,�>�P���t��� �����]�����(� :�L�^���������� ����k� $6H Z��~����� �y 2DVh �������v�KRC�i���!� ��/S/B/w/f/�/�/��/��SBL_FA?ULT j*6�>�!GPMSK���'���TDIAG ik��-�������UD1: 6�78901234A5I2��=1�Ǥ�P\� �?�?�?�?�?�?�?O O'O9OKO]OoO�O�O �Od696���r
t?�O>|�TRECP"?4:
B44_[7��s?p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�O��O�O�o7�UMP__OPTIO=��.F�aTR����)u�PME��Y_T�EMP  ÈW�3BC�gp�B�QtUNI����gq��YN_BRK �lL�7�EDITO�R�a�a@�r_
PE�NT 1m) � ,&TELGEOP^P ����p�PSNA�:�&MTPG�p+�=� �/��I�z�����ۏ ����5��Y�k�R� ��v���ş���П� ���C�*�g�N�v��� ���������ޯ���?�Q���EMGDI_STAzuV�gq��uNC_INFO� 1n!��b����X���������n�1o!� ��o���
�
�d�oU�g�y� �ϝϯ���������	� �-�?�Q�c�u߇ߙ� �߽��� u����
�� *�B�*�P�b�t��� �����������(� :�L�^�p��������� 2�������9�C Ugy����� ��	-?Qc u�������� //1;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?��?�?�?O)/O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�?�?�_ �_o�_3O=oOoaoso �o�o�o�o�o�o�o '9K]o�� ��_�_����+o 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y��������ӟ ���	�#�-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� �7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߹��� �������%�/�A�S� e�w��������� ����+�=�O�a�s� �������������� �'9K]o�� ������# 5GYk}�	�� ����/1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?��?�?�?�? /O)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�? �_�_�_�_O�_!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew��_�_��� �o�+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o���� ���ɟ۟���#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� ���߹���������� %�7�I�[�m���� �����������!�3� E�W�i�{��߇����� �����/AS ew������ �+=Oas ����������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?���?�? �?�?��?OO1OCO UOgOyO�O�O�O�O�O �O�O	__-_?_Q_c_ u_�?�_�_�_�_�?�_ oo)o;oMo_oqo�o �o�o�o�o�o�o %7I[m�_u� ���_���!�3� E�W�i�{�������Ï Տ�����/�A�S� e��������u�� ����+�=�O�a�s� ��������ͯ߯�� �'�9�K�]�w����� ����ɿ�����#� 5�G�Y�k�}Ϗϡϳ� ����������1�C� U�g߁��ߝ߯���ۿ ����	��-�?�Q�c� u����������� ��)�;�M�_�y߃� ������������ %7I[m�� �����!3 EWq�c����� ����////A/S/ e/w/�/�/�/�/�/�/ �/??+?=?O?i{ �?�?�?�?��?�?O O'O9OKO]OoO�O�O �O�O�O�O�O�O_#_ 5_G_�?s?}_�_�_�_ �?�_�_�_oo1oCo Uogoyo�o�o�o�o�o �o�o	-?Qk_ u����_��� ��)�;�M�_�q��� ������ˏݏ��� %�7�I�cQ������ ���ٟ����!�3� E�W�i�{�������ï կ�����/�A�[�� �$ENETM�ODE 1p����  
k�k�f�����j��OATCFG �q�����Ѵ��C���DAT�A 1rw�Ӱ�.��*	�*��'�9�K�]�l�dlύ�e��ϻ�������� �'ߡϳ�]�o߁ߓ� �߷�1���U����#� 5�G�Y����ߏ��� ��������u��1�C� U�g�y������)��� ����	-����c�u�����j�RPOST_LO��	t�[
׶#5�Gi�RROR_P-R� %w�%L��XTABLE  w�ȟ�����RSEV_NUM� ��  ����  �_AUT�O_ENB  ����X_NO5! �uw���" W *�x �x �x 	�x + +w �/�/�/�Q$FLTR=/O&H�IS#]�J+_A�LM 1vw� e�[x,e�+�/�Q?c?u?�?�?�?�/_\"W   w�v!����:j�TCP_V_ER !w�!x޻?$EXT� _R�EQ�&�H)BCSsIZKO=DSTKhI�f%�?BTOL�  ]Dz�"��A =D_BWD��0�@�&�A���CDI�A wķ���]�KSTEP�O�Oj�>POP_DO�Oh��FDR_GRP s1xw��!d 	�?x�_��yPs�Y�Q�'�M"����l��T� ����VyS�_�]��TBIZA���Aqn�@  A火N�_�P���A��A=d� bd�]Go�_Wo}oho�o�o�o�]@g%2�@&��?��>��>�n
 �Lay] a�a]?��L"#~�3:�o^�I��XA@`�t@'S33�uh}@�q��g��yPF@ x��|yPG�  @��Fg�fC�8R�L��}?�pi��~6��X����875�t��5���5�`+��}�O�����~���j����%��:�3����[�FEATURE y����@��Ha�ndlingTo�ol �]E�nglish D�ictionar}y�4D St���ard��Analog I/O>��G�gle Shi�ftZ�uto S�oftware �Update�m�atic Bac�kup���gro�und Edit� ��Camera�U�FY�CnrRn�dIm���omm�on calib' UI��nˑ�Monitor$��tr�Reliaybn��DHCP ��[�ata Acq�uis3�\�iag�nos��R�v�is�playΑLic�ensZ�`�ocu�ment Vie�we?�^�ual �Check Sa�fety��ha�nced���s��Frܐ�xt.� DIO /�fiܬ�@�end�ErEr>�L��\�4�s[��rP�K� �@
�FCTN Menu���vZ���TP InΝ�facĵ�Gi�gE־�Đp Mask Exc��g=�HT԰Pro�xy Sv��i�gh-Spe�S�ki�� Ť�O�mm�unic��onsV�ur����q�V�ײ�connect �2��ncrְst#ru!��ʴ�eۡ���J��X�KAREL Cmd. L��ua���Run-;Ti<�Env�Ȟ��el +��s��S�/W�ƥ���r�B�ook(Syst�em)
�MACR�Os,M�/Offseu�p�HO���o��u�MR8�4���Me�chStop+�t�����p�im�q���x��R�����odo�w�itch�ӟ�.<��4�OptmF��N,�fil䬳�g��~p�ulti-T��Γ�PCM fu	n�Ǽ�o��������/Regie�rq���riݠF���S�N?um Sel��/�>:� Adjua�*�xW�q�h�tatu����ߪ�RDM R�obot�sco3ve'���ea��<��Freq Anl�yq�Rem��O�n�5�����Servo�O�!��SNPX �b-�v�SN԰Cl�iܡ?r�Libr�&�_�� ��q +ozJ�t��ssag��X�@ ����	�@/�Iս�MILIB���P Firmt���P��AccŐ�͛TPTXk��eln���������orquo�imu�la=��|u(�PAa&��ĐX�B�&+�gev.���ri���TUSB po�rt �iPf�a�ݠ&R EVNT�� nexcep�t�����%5��VEC�rl�c���V����"�%q�+SR S9CN�/SGE�/�%�UI	�Web Pl��>��A43���ۡ��ZDT Ap�plj�
�{1EOA�T����&0?�7G�rid�񾡬=�?iR�".5� F���/�גRX-10iA�/L�?Alarm Cause/���ed(�All Smooth5���C��scii+�V�Losad䠌JUpl�@�w�toS ��ri�tyAvoidM�(�s7�t�@�y�cn�����_�C9S+���. c��XJo���-T3_H�.R�X��U���Xcol�labo����RA`�:�.9D��in����NRTHI
�O}n��e Hel�����ֿ�����1tr�U�ROS Eth $��A������;,�Ga �B�,|HUpV�%�W�t ԰�_i�RS�ݐ�64MB� DRAM�o�cF�RO���L8F F!lD�����2M �A:�opm�ԕex@V�
�#sh�q��wce�u���p��|tyn�sA�
�%�r����J��b^�.v� P)Q/sbS��`���O�N��ma�i��U���R�q6�T1�^FC+Ԍ%̋Fs9�ˌk̋��Typ߽FC%�h�ױV�N Sp�For0ްK��Ԭ�lu!���<�cp�PG j�֡��RJ�[L`Sup�"}��֐f��cr�FP��lu� ��al�����r��i�
q��4@а�uest~,IMPLE ׀ 6*|HZ���c0�B�Tea(�|���$r�tu���V�9HMI��¤��UIFc�pono2D�BC�:� L�y�p���������ʿ ܿ	� ��?�6�H�u� l�~ϫϢϴ������ ���;�2�D�q�h�z� �ߞ߰��������
� 7�.�@�m�d�v��� ����������3�*� <�i�`�r��������� ������/&8e \n������ ��+"4aXj �������� '//0/]/T/f/�/�/ �/�/�/�/�/�/#?? ,?Y?P?b?�?�?�?�? �?�?�?�?OO(OUO LO^O�O�O�O�O�O�O �O�O__$_Q_H_Z_ �_~_�_�_�_�_�_�_ oo oMoDoVo�ozo �o�o�o�o�o�o
 I@Rv�� �������E� <�N�{�r�������Տ ̏ޏ���A�8�J� w�n�������џȟڟ ����=�4�F�s�j� |�����ͯį֯��� �9�0�B�o�f�x��� ��ɿ��ҿ�����5� ,�>�k�b�tφϘ��� ���������1�(�:� g�^�p߂ߔ��߸��� ���� �-�$�6�c�Z� l�~���������� ��)� �2�_�V�h�z� ��������������% .[Rdv�� �����!* WN`r���� ���//&/S/J/ \/n/�/�/�/�/�/�/ �/??"?O?F?X?j? |?�?�?�?�?�?�?O OOKOBOTOfOxO�O �O�O�O�O�O___ G_>_P_b_t_�_�_�_ �_�_�_oooCo:o Lo^opo�o�o�o�o�o �o	 ?6HZ l������� ��;�2�D�V�h��� ����ˏԏ���
� 7�.�@�R�d������� ǟ��П�����3�*� <�N�`�������ï�� ̯����/�&�8�J� \�����������ȿ�� ���+�"�4�F�Xυ� |ώϻϲ��������� '��0�B�T߁�xߊ� �߮���������#�� ,�>�P�}�t���� ����������(�:� L�y�p����������� ����$6Hu�l~������  H55�2��21R7�850J61�4ATUP'5�45'6VCA�MCRIbUI�F'28cNREv52VR63wSCHLIC��DOCV�CSU�869'02E�IOC�4R6=9VESET?U�J7UR68M�ASKPRXY�{7OCO#(3�?+ &3j&J6�%53�H�(LC�HR&OPLG?0^�&MHCRS&S�'�MCS>0.'55�2MDSW+7u'OPu'MPRv&��(�0&PCMzR0`q7+ 2� �'51J�51�80JPRSv"'69j&FRDb�FREQMCN�93&SNBA���'SHLBFM�1G�82&HTC�>TMIL�T{PA�TPTXcF#ELF� �8�J95�TUTvv'95j&UEV"&wUECR&UFRb�VCC
XO�&VI�PnFCSC�FCS�G��IWEBn>HTT>R6�شH;RVCGiWIG�QWIPGS�VRC�nFDGu'H7�7RK66J5'R�8WR51
(6�(2�(I5V�J8�86��L=I% �84g6�62R64NV�D"&R6�'R84ֺg79�(4�S5ni'J76j&D0�g�F xRTSFCR�gCRXv&CLIZ8ICMS�Sp>�STYnG6)7CT�O>��7�NN�j&ORS�&C &F�CB�FCF�7C�H>FCR"&FC-I�VFC�'J�PO7�GBfM�8OLaxE�NDS&LU�&CPUR�7LWS�xC��STxTE�gS60nFVR�IN�7IHaF�я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{������ �/ASew �������/ /+/=/O/a/s/�/�/ �/�/�/�/�/??'? 9?K?]?o?�?�?�?�? �?�?�?�?O#O5OGO YOkO}O�O�O�O�O�O �O�O__1_C_U_g_ y_�_�_�_�_�_�_�_ 	oo-o?oQocouo�o �o�o�o�o�o�o );M_q��� ������%�7� I�[�m��������Ǐ�ُ�  �H552��21n�R78�50��J614�ATU]P7�5457�6��VCAM�CRIn��UIF7�28���NRE�52v�R�63�SCH�L{ICƚDOCV�wCSU�8697��0F�EIOCǛ4��R69v�ESE�TW�u�J7u�R6�8�MASK�P�RXY��7�OC�O��3W����6�3��J65�536�H�$�LCHƪOPL�GW�0�MHCR�ǪS��MCSV�0���55F�MDSW����OP��MPR����6�06�PCM��R0E˓�F���6�[51f�51��0f��PRS��69�F{RD��FREQ��MCN�936�S�NBAכ%�SHLEB�ME��ּ26��HTCV�TMIL��6�TPAV�TPTX��ELړ�6�q8%�#��J95���TUT��95�U�EV��UECƪU�FR��VCCf�OVIP��CSCN��CSGƚ$�I�wWEBV�HTTV��R6՜��S���CG���IG��IPGS�'�RC��DG��H]7��R66f�5��u�R��R51f�6J�2�5v�#�J׼
��6��LU�5�s�v��4��66F�R64n�NVD��R6���R84�79�4v��S5�J76��D0uFRTSv&�CR�CRX���CLI&�e�CMS�V�sV�STY��6��CTOV�#�V�7v5�NN�ORS��ܳ�6�FCBV�FC�F��CHV�FCRn��FCIF�FC���J#��G
M��O�L�ENDǪLU���CPR��Lu�Sj�C$�StTE�wS60�FVRV�IN��IH���m? ?�?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�O__ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o'9K] o������� ��#�5�G�Y�k�}� ������ŏ׏���� �1�C�U�g�y����� ����ӟ���	��-� ?�Q�c�u��������� ϯ����)�;�M� _�q���������˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �!�3�E�W�i�{ߍ� �߱����������� /�A�S�e�w���� ����������+�=� O�a�s����������� ����'9K] o������� �#5GYk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏�ߏ�STD~�LANG� ��0�B�T�f�x��� ������ҟ����� ,�>�P�b�t������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��� �2�D�V�h�z�p�ߞ߰���RBT
�OPTN������ '�9�K�]�o����p��������DPN	� ��)�;�M�_�q��� ������������ %7I[m�� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�? OO'O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_oo1o CoUogoyo�o�o�o�o �o�o�o	-?Q cu������ ���)�;�M�_�q� ��������ˏݏ�� �%�7�I�[�m���� ����ǟٟ����!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩϻ������� ��'�9�K�]�o߁� �ߥ߷���������� #�5�G�Y�k�}��� ������������1� C�U�g�y��������� ������	-?Qc�f�������99��$F�EAT_ADD �?	���~  	� #5GYk}�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ���������DEMO �y   �L�B�T߁�xߊ� �߮����������� G�>�P�}�t���� ����������C�:� L�y�p����������� ����?6Hu l~������ ;2Dqhz ������ /
/ 7/./@/m/d/v/�/�/ �/�/�/�/�/?3?*? <?i?`?r?�?�?�?�? �?�?�?O/O&O8OeO \OnO�O�O�O�O�O�O �O�O+_"_4_a_X_j_ �_�_�_�_�_�_�_�_ 'oo0o]oTofo�o�o �o�o�o�o�o�o# ,YPb���� ������(�U� L�^�����������ʏ ����$�Q�H�Z� ��~�������Ɵ��� �� �M�D�V���z� ������¯ܯ��
� �I�@�R��v����� ����ؿ����E� <�N�{�rτϱϨϺ� �������A�8�J� w�n߀߭ߤ߶����� ����=�4�F�s�j� |����������� �9�0�B�o�f�x��� ������������5 ,>kbt��� ����1(: g^p����� �� /-/$/6/c/Z/ l/�/�/�/�/�/�/�/ �/)? ?2?_?V?h?�? �?�?�?�?�?�?�?%O O.O[OROdO�O�O�O �O�O�O�O�O!__*_ W_N_`_�_�_�_�_�_ �_�_�_oo&oSoJo \o�o�o�o�o�o�o�o �o"OFX� |������� ��K�B�T���x��� ����ۏҏ���� G�>�P�}�t������� ןΟ�����C�:� L�y�p�������ӯʯ ܯ	� ��?�6�H�u� l�~�����Ͽƿؿ� ���;�2�D�q�h�z� �Ϟ����������
� 7�.�@�m�d�vߐߚ� �߾��������3�*� <�i�`�r������ �������/�&�8�e� \�n������������� ����+"4aXj �������� '0]Tf�� ������#// ,/Y/P/b/|/�/�/�/ �/�/�/�/??(?U? L?^?x?�?�?�?�?�? �?�?OO$OQOHOZO tO~O�O�O�O�O�O�O __ _M_D_V_p_z_ �_�_�_�_�_�_o
o oIo@oRolovo�o�o �o�o�o�oE <Nhr���� �����A�8�J� d�n�������яȏڏ ����=�4�F�`�j� ������͟ğ֟��� �9�0�B�\�f����� ��ɯ��ү�����5� ,�>�X�b�������ſ ��ο����1�(�:� T�^ϋςϔ��ϸ��� ���� �-�$�6�P�Z� ��~ߐ߽ߴ������� ��)� �2�L�V��z� ������������%� �.�H�R��v����� ����������!* DN{r���� ���&@J wn������ �//"/</F/s/j/ |/�/�/�/�/�/�/? ??8?B?o?f?x?�? �?�?�?�?�?OOO 4O>OkObOtO�O�O�O��O�O�O__0]  'XF_X_j_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o �o�o�o�o�o, >Pbt���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п�����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ���(:L ^p������ � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?V?h?z?�? �?�?�?�?�?�?
OO .O@OROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo\o no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x����� ����ҏ�����,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
��>.�  /�)� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX j|������ ���0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ��������� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� ����������&�8� J�\�n����������� ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸπ������ ��$�4�8�+�N�`�r߄ߖ� �ߺ���������&� 8�J�\�n����� ���������"�4�F� X�j�|����������� ����0BTf x������� ,>Pbt� ������// (/:/L/^/p/�/�/�/ �/�/�/�/ ??$?6? H?Z?l?~?�?�?�?�? �?�?�?O O2ODOVO hOzO�O�O�O�O�O�O �O
__._@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�o �o�o�o�o�o& 8J\n���� �����"�4�F� X�j�|�������ď֏ �����0�B�T�f� x���������ҟ��� ��,�>�P�b�t��� ������ί���� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢϴ��� ������� �2�D�V� h�zߌߞ߰������� ��
��.�@�R�d�v� ������������ �*�<�N�`�r����� ����������& 8J\n���� ����"4F Xj|����� ��//0/B/T/f/ x/�/�/�/�/�/�/�/ ??,?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�O �O�O�O�O __$_6Y��$FEAT_D�EMOIN  V;T�fP�<PNT_INDEX[[jQ��NPILECOM�P z�����QiRIU�PS�ETUP2 {��U�R�  �N �Q�S_AP2�BCK 1|�Y  �)7Xok%�_8o<P�P&oco 9U�_�oo�oBo�o�o xo�o1C�og�o ��,�P��� ��?��L�u���� (���Ϗ^�󏂏�)� ��M�܏q������6� ˟Z�؟���%���I� [��������D�ٯ h������3�¯W�� d������@�տ�v� Ϛ�/�A�пe����� ��*Ͽ�N���r���� ��=���a�s�ߗ�&� ����\��߀��'�� K���o���|��4��� X������#���G�Y� ��}������B���f�@����1�Y�PP�_� 2�P*.V1R8���*��`�����l PC�|��FR6:�"2�V�TzPz �w�]PG����*.Fo/��	��:,�^/�STMi/�/ /�-M/�/�H�/?�'�?�/�/g?�GIF q?�?�%�?D?V?�?�JPG�?O�%O�?�?oO�
JSyO�O���5C�OMO%
Ja�vaScript�O�?CS�O&_�&_��O %Casc�ading St�yle Shee�tsR_��
ARGNAME.DT�_
��� \�_S_�A�T��_�_�PDISP	*�_���To�_�Q�LaZooCLLB�.ZIwo2o$ :\ҝa\�o�i�ACo�llabo�o�o
�TPEINS.X3ML�_:\![o��QCustom Toolbarb�iPASSWOR�DQo��FRS:�\�dB`Pass�word Config���/��(� e��������N�� r�����=�̏a��� ���&���J���񟀟 ���9�K�ڟo����� ��4�ɯX��|���#� ��G�֯@�}����0� ſ׿f������1��� U��y��ϯ�>��� b���	ߘ�-߼�Q�c� �χ�߽߫�L���p� �ߦ�;���_���X� ��$��H�����~�� ��7�I���m���� � 2���V���z���!�� E��i{
�.� �d����S �wp�<�` �/�+/�O/a/� �//�/8/J/�/n/? �/�/9?�/]?�/�?�? "?�?F?�?�?|?O�? 5O�?�?kO�?�OO�O �OTO�OxO__�OC_ �Og_y__�_,_�_P_ b_�_�_o�_oQo�_ uoo�o�o:o�o^o�o �o)�oM�o�o� �6��l�� %�7��[����� � ��D�ُh�z����3� ,�i��������ß�R��v������$�FILE_DGB�CK 1|������� < �)
SU�MMARY.DG<!�͜MD:U����ِDiag Summary�����
CONSLO�G��n���ٯ����Console �log���	TPOACCN�t�%\������TP Accountin;����FR6:IP�KDMP.ZIP�Ϳј
�ϥ���E�xception�"�ӻ��MEMCH�ECK���������-�Memory �Data����J�n )��RIPE��~ϐ�%ߴ�%��� Packet� L:���L�$�<c���STAT��|߭� %A�?Status��^�	FTP����	����/�mment� TBD2�^� >�I)ETHERNEw�
�d�u�﨡EthernJ�~1�figuraA�����DCSVRF�&���7����� �verify a�ll:��� 4��DIFF/��'�x��;�Q�diff���r�d���CHG01 ������A����it�2���270���fx3����I �p��VTRNDIAG.LSu&8���=� Ope��L�� ��nostic���c�)VD;EV�DAT��x����Vis�?Device�+IMG��,/>/�/z:�i$Imagu/n+UP ES/~�/FRS:\?�Z=��Updates ListZ?���� FLEXEVEN��/�/�?����1 UIF E�vM�M���-vZ�)CRSENSSPK�/˞�\!Oܸ��CR_TAOR�_PEAKbOͩP�SRBWLD.C	M�O͜E2�O\?.��PS_ROBOW�ELS���:GIG���@_�?d_��Gi�gE�(O��N�@��)UQHADO�W__D_V_�_��S�hadow Ch�ange����@d�t�RRCMERR��_�_�_oo��4`C�FG Error�o tailo M�A�k�CMSGLIBgoNo`o�o|R��e��z0ic�o�a7�)�`ZD0_O��os��ZD�Pa�d�l �RNO�TI�Rd���Notific��<���,�AG��P� ӟt���������Ώ]� ����(���L�^�� �������G�ܟk� � ���6�şZ��~��� ���C�د�y���� 2�D�ӯh�������� ¿Q��u�
�ϫ�@� Ͽd�v�Ϛ�)Ͼ��� _��σ�ߧ�%�N��� r�ߖߨ�7���[��� ��&��J�\��߀� ��3����i���� "�4���X���|���� ��A�����w���0 ��=f����� O�s�>� bt�'�K� ��/�:/L/�p/ ��/�/5/�/Y/�/ ? �/$?�/H?�/U?~?? �?1?�?�?g?�?�? O 2O�?VO�?zO�OO�O ?O�OcO�O
_�O._�O R_d_�O�__�_�_M_ �_q_oo�_<o�_`o �_mo�o%o�oIo�o�o o�o8J�on�o ��3�W�{� "��F��j�|���� /�ď֏e������0���$FILE_F�RSPRT  ��������?�MDON�LY 1|S��� 
 �)M�D:_VDAEX?TP.ZZZ1�����ț6%N�O Back f�ile ���S�6P�����>��K� t�����'���ί]�� ���(���L�ۯp��� ���5�ʿY�׿ Ϗ� $ϳ�H�Z��~�Ϣ� ��C���g���ߝ�2� ��V���cߌ�߰�?� ����u�
��.�@����d��߈��C�VIS�BCKq�[���*�.VD����S�F�R:\��ION\�DATA\��v��S�Vision VD���Y�k� ���y��B�����x� ��1C��g��� ,�P��� �?�Pu�( ��^��/�� M/�q/�/>/�/6/�/ Z/�/?�/%?�/I?[? �/??�?2?D?�?9��LUI_CONF�IG }S�|���; $ �3v�{S�;OMO_OqO�O�O�I#@|x�?�O�O �O__%\�OH_Z_l_ ~_�_'_�_�_�_�_�_ o�_2oDoVohozo�o #o�o�o�o�o�o
�o .@Rdv�� ������*�<� N�`�r��������̏ ޏ�����&�8�J�\� n��������ȟڟ� ����"�4�F�X�j�� ������į֯��� �0�B�T�f������� ����ҿ�{���,� >�P�b����ϘϪϼ� ����w���(�:�L� ^��ςߔߦ߸����� s� ��$�6�H���Y� ~������]����� � �2�D���h�z��� ������Y�����
 .@��dv��� �U��*< �`r����Q ��//&/8/�\/ n/�/�/�/;/�/�/�/ �/?"?�/F?X?j?|? �?�?7?�?�?�?�?O O�?BOTOfOxO�O�O 3O�O�O�O�O__�O >_P_b_t_�_�_/_�_ �_�_�_oo�_:oLo�^opo�o�o$h  �x�o�c�$FL�UI_DATA �~����a�(a�dRESULT 3�e�p �T��/wizard�/guided/�steps/Expert�o=Oa s���������z�Conti�nue with{ Gpance� :�L�^�p����������ʏ܏� � �b-��a�e�0 �`0`��c�a?��ps���������ҟ �����,�>�P�� 0ow���������ѯ� ����+�=�O�a�?��1�C�U�e�cllbs�ֿ�����0� B�T�f�xϊϜ�[��� ��������,�>�P� b�t߆ߘߪ�i�{���t��]�e�rip(p ſ-�?�Q�c�u��� �����������)� ;�M�_�q��������� �������������`�e�#pTime?US/DST	� ������!�3E�Enabl(�y��������	//-/?/Q/�b�)�/M_q24|�/�/??)? ;?M?_?q?�?�?Tf �?�?�?OO%O7OIO [OmOO�O�Ob/t/�/�/Z�"qRegion�O5_G_Y_k_}_��_�_�_�_�_�_�America!� #o5oGoYoko}o�o�o@�o�o�o�o��Ay�O��O3�O_qEditor�o���� �����+�=� �� Touch P�anel rs (�recommenp�)K�������Ə؏����� �2�D�|��%��I[qaccesoܟ� �� $�6�H�Z�l�~������Connect� to Network��֯���� �0�B�T�f�x�����
x��@��}����,�!��s Introduct!_4�F�X� j�|ώϠϲ������� ���0�B�T�f�x߀�ߜ߮��������� ɿ��"�i� {������������ ��/�A� �e�w��� �������������+=�H�3�� +�O�����  2DVhz� K������
// ./@/R/d/v/�/�/Y k}�/�??*?<? N?`?r?�?�?�?�?�? �?��?O&O8OJO\O nO�O�O�O�O�O�O�O �/_�/1_�/X_j_|_ �_�_�_�_�_�_�_o o0oBoS_foxo�o�o �o�o�o�o�o, >�O_!_�E_�� �����(�:�L� ^�p�����So��ʏ܏ � ��$�6�H�Z�l� ~���O��s՟��� � �2�D�V�h�z��� ����¯ԯ毥�
�� .�@�R�d�v������� ��п⿡��ş'�9� ��`�rτϖϨϺ��� ������&�8���\� n߀ߒߤ߶������� ���"�4��=��a� ��Mϲ���������� �0�B�T�f�x���I� ����������, >Pbt�E��i� ����(:L ^p������ �� //$/6/H/Z/l/ ~/�/�/�/�/�/�� ��/?�V?h?z?�? �?�?�?�?�?�?
OO .O�ROdOvO�O�O�O �O�O�O�O__*_<_ �/??�_C?�_�_�_ �_�_oo&o8oJo\o no�o?O�o�o�o�o�o �o"4FXj| �M___q_��_�� �0�B�T�f�x����� ����ҏ�o���,� >�P�b�t��������� Ο�����%��L� ^�p���������ʯܯ � ��$�6�G�Z�l� ~�������ƿؿ��� � �2��S��w�9� �ϰ���������
�� .�@�R�d�v߈�G��� ����������*�<� N�`�r��Cϥ�g��� �ύ���&�8�J�\� n��������������� ��"4FXj| ���������� -��Tfx�� �����//,/ ��P/b/t/�/�/�/�/ �/�/�/??(?�1 U??A�?�?�?�? �? OO$O6OHOZOlO ~O=/�O�O�O�O�O�O _ _2_D_V_h_z_9? �?]?�_�_�?�_
oo .o@oRodovo�o�o�o �o�o�O�o*< N`r����� �_�_�_�_#��_J�\� n���������ȏڏ� ���"��oF�X�j�|� ������ğ֟���� �0����u�7��� ����ү�����,� >�P�b�t�3������� ο����(�:�L� ^�pς�A�S�e��ω� �� ��$�6�H�Z�l� ~ߐߢߴ��߅����� � �2�D�V�h�z�� ������������ ��@�R�d�v������� ��������*;� N`r����� ��&��G	� k-������� �/"/4/F/X/j/|/ ;�/�/�/�/�/�/? ?0?B?T?f?x?7�? [�?�?�?OO,O >OPObOtO�O�O�O�O �O�/�O__(_:_L_ ^_p_�_�_�_�_�_�? �_�?o!o�OHoZolo ~o�o�o�o�o�o�o�o  �ODVhz� ������
�� �_%o�_I�s�5o���� ��Џ����*�<� N�`�r�1������̟ ޟ���&�8�J�\� n�-�w�Q���ů��� ���"�4�F�X�j�|� ������Ŀ������ �0�B�T�f�xϊϜ� ������������ٯ >�P�b�t߆ߘߪ߼� ��������տ:�L� ^�p��������� �� ��$������i� +ߐ�������������  2DVh'� ������
 .@Rdv5�G�Y� �}���//*/</ N/`/r/�/�/�/�/y �/�/??&?8?J?\? n?�?�?�?�?�?��? �O�4OFOXOjO|O �O�O�O�O�O�O�O_ _/OB_T_f_x_�_�_ �_�_�_�_�_oo�? ;o�?_o!O�o�o�o�o �o�o�o(:L ^p/_����� � ��$�6�H�Z�l� +o��Oo��sou���� � �2�D�V�h�z��� ��������
�� .�@�R�d�v������� ��}�߯����ٟ<� N�`�r���������̿ ޿���ӟ8�J�\� nπϒϤ϶������� ���ϯ��=�g�)� �ߠ߲���������� �0�B�T�f�%ϊ�� ������������,� >�P�b�!�k�Eߏ��� {�����(:L ^p����w�� � $6HZl ~���s������� /��2/D/V/h/z/�/ �/�/�/�/�/�/
?� .?@?R?d?v?�?�?�? �?�?�?�?OO�� �]O/�O�O�O�O�O �O�O__&_8_J_\_ ?�_�_�_�_�_�_�_ �_o"o4oFoXojo)O ;OMO�oqO�o�o�o 0BTfx�� �m_�����,� >�P�b�t��������� {oݏ�o��o(�:�L� ^�p���������ʟܟ � ��#�6�H�Z�l� ~�������Ưد��� �͏/��S��z��� ����¿Կ���
�� .�@�R�d�#��ϚϬ� ����������*�<� N�`����C���g�i� ������&�8�J�\� n�����u����� ���"�4�F�X�j�|� ������q�������	 ��0BTfx�� �������, >Pbt���� ���/����1/ [/�/�/�/�/�/�/ �/ ??$?6?H?Z? ~?�?�?�?�?�?�?�? O O2ODOVO/_/9/ �O�Oo/�O�O�O
__ ._@_R_d_v_�_�_�_ k?�_�_�_oo*o<o No`oro�o�o�ogOyO �O�O�o�O&8J\ n������� ��_"�4�F�X�j�|� ������ď֏���� �o�o�oQ�x����� ����ҟ�����,� >�P��t��������� ί����(�:�L� ^��/�A���e�ʿܿ � ��$�6�H�Z�l� ~ϐϢ�a��������� � �2�D�V�h�zߌ� �߰�o��ߓ��߷�� .�@�R�d�v���� ����������*�<� N�`�r����������� ������#��G	� n������� �"4FX�| �������/ /0/B/T/u/7�/ []/�/�/�/??,? >?P?b?t?�?�?�?i �?�?�?OO(O:OLO ^OpO�O�O�Oe/�O�/ �O�O�?$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ �? o2oDoVohozo�o �o�o�o�o�o�o�O_ �O%O_v��� ������*�<� N�or���������̏ ޏ����&�8�J�	 S-w���cȟڟ� ���"�4�F�X�j�|� ����_�į֯���� �0�B�T�f�x����� [�m����󿵟�,� >�P�b�tφϘϪϼ� �����ϱ��(�:�L� ^�p߂ߔߦ߸����� �� ￿ѿ�E��l� ~������������ � �2�D��h�z��� ������������
 .@R�#�5�Y� ����*< N`r��U��� ��//&/8/J/\/ n/�/�/�/c�/��/ �?"?4?F?X?j?|? �?�?�?�?�?�?�?? O0OBOTOfOxO�O�O �O�O�O�O�O�/_�/ ;_�/b_t_�_�_�_�_ �_�_�_oo(o:oLo Opo�o�o�o�o�o�o �o $6H_i +_�O_Q���� � �2�D�V�h�z��� ��]oԏ���
�� .�@�R�d�v�����Y ��}ߟ񟵏�*�<� N�`�r���������̯ ޯ𯯏�&�8�J�\� n���������ȿڿ� ����ϟ�C��j�|� �Ϡϲ���������� �0�B��f�xߊߜ� ������������,� >���G�!�k��Wϼ� ��������(�:�L� ^�p�����S߸����� �� $6HZl ~�O�a�s�����  2DVhz� �������
// ./@/R/d/v/�/�/�/ �/�/�/�/���9? �`?r?�?�?�?�?�? �?�?OO&O8O�\O nO�O�O�O�O�O�O�O �O_"_4_F_??)? �_M?�_�_�_�_�_o o0oBoTofoxo�oIO �o�o�o�o�o, >Pbt��W_� {_��_��(�:�L� ^�p���������ʏ܏ ���$�6�H�Z�l� ~�������Ɵ؟꟩ ��/��V�h�z��� ����¯ԯ���
�� .�@���d�v������� ��п�����*�<� ��]����C�EϺ��� ������&�8�J�\� n߀ߒ�Q��������� ���"�4�F�X�j�|� ��Mϯ�q������� �0�B�T�f�x����� ����������, >Pbt���� ��������7�� ^p������ � //$/6/��Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?�;_?�? K�?�?�?�?�?
OO .O@OROdOvO�OG/�O �O�O�O�O__*_<_ N_`_r_�_C?U?g?y? �_�?oo&o8oJo\o no�o�o�o�o�o�o�O �o"4FXj| �������_�_ �_-��_T�f�x����� ����ҏ�����,� �oP�b�t��������� Ο�����(�:�� ���A�����ʯܯ � ��$�6�H�Z�l� ~�=�����ƿؿ��� � �2�D�V�h�zό� K���o��ϓ���
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� �������#���J�\� n��������������� ��"4��Xj| ������� 0��Q�u7�9 �����//,/ >/P/b/t/�/E�/�/ �/�/�/??(?:?L? ^?p?�?A�?e�?�? �/ OO$O6OHOZOlO ~O�O�O�O�O�O�/�O _ _2_D_V_h_z_�_ �_�_�_�_�?�?�?o +o�?Rodovo�o�o�o �o�o�o�o*�O N`r����� ����&��_/o	o S�}�?o����ȏڏ� ���"�4�F�X�j�|� ;����ğ֟���� �0�B�T�f�x�7�I� [�m�ϯ������,� >�P�b�t��������� ο�����(�:�L� ^�pςϔϦϸ����� ������!��H�Z�l� ~ߐߢߴ��������� � �߿D�V�h�z�� �����������
�� .������s�5ߚ��� ��������*< N`r1���� ��&8J\ n�?��c����� �/"/4/F/X/j/|/ �/�/�/�/�/��/? ?0?B?T?f?x?�?�? �?�?�?��?�O� >OPObOtO�O�O�O�O �O�O�O__(_�/L_ ^_p_�_�_�_�_�_�_ �_ oo$o�?EoOio +O-o�o�o�o�o�o�o  2DVhz9_ ������
�� .�@�R�d�v�5o��Yo ��͏����*�<� N�`�r���������̟ ����&�8�J�\� n���������ȯ��я ������F�X�j�|� ������Ŀֿ���� �ݟB�T�f�xϊϜ� ������������ٯ #���G�q�3��ߪ߼� ��������(�:�L� ^�p�/ϔ������� �� ��$�6�H�Z�l� +�=�O�a���������  2DVhz� �������
 .@Rdv��� ��������/��</ N/`/r/�/�/�/�/�/ �/�/??�8?J?\? n?�?�?�?�?�?�?�? �?O"O��/gO)/ �O�O�O�O�O�O�O_ _0_B_T_f_%?w_�_ �_�_�_�_�_oo,o >oPoboto3O�oWO�o {O�o�o(:L ^p������o � ��$�6�H�Z�l� ~�������Ə�o珩o ��o2�D�V�h�z��� ����ԟ���
�� �@�R�d�v������� ��Я�����׏9� ��]��!�������̿ ޿���&�8�J�\� n�-��Ϥ϶������� ���"�4�F�X�j�)� ��M����߅������ �0�B�T�f�x��� �����������,� >�P�b�t��������� {��ߟ�����:L ^p������ � ��6HZl ~������� /����;/e/'�/ �/�/�/�/�/�/
?? .?@?R?d?#�?�?�? �?�?�?�?OO*O<O NO`O/1/C/U/�Oy/ �O�O__&_8_J_\_ n_�_�_�_�_u?�_�_ �_o"o4oFoXojo|o �o�o�o�o�O�O�O	 �O0BTfx�� �������_,� >�P�b�t��������� Ώ������o�o�o [���������ʟܟ � ��$�6�H�Z�� k�������Ưد��� � �2�D�V�h�'��� K���o�Կ���
�� .�@�R�d�vψϚϬ� ��Ͽ������*�<� N�`�r߄ߖߨߺ�y� �ߝ�����&�8�J�\� n����������� �����4�F�X�j�|� �������������� ��-��Q��� �����, >Pb!����� ���//(/:/L/ ^//A�/�/y�/ �/ ??$?6?H?Z?l? ~?�?�?�?s�?�?�? O O2ODOVOhOzO�O �O�Oo/�/�/�O_�/ ._@_R_d_v_�_�_�_ �_�_�_�_o�?*o<o No`oro�o�o�o�o�o �o�o�O_�O/Y _������� ��"�4�F�X�o|� ������ď֏���� �0�B�T�%7I ��mҟ�����,� >�P�b�t�������i� ί����(�:�L� ^�p���������w��� ������$�6�H�Z�l� ~ϐϢϴ��������� �� �2�D�V�h�zߌ� �߰���������
�ɿ ۿ�O��v���� ����������*�<� N��_����������� ����&8J\ �}?�c���� �"4FXj| �������/ /0/B/T/f/x/�/�/ �/m�/��/�?,? >?P?b?t?�?�?�?�? �?�?�?O�(O:OLO ^OpO�O�O�O�O�O�O �O _�/!_�/E_?	_ ~_�_�_�_�_�_�_�_ o o2oDoVoOzo�o �o�o�o�o�o�o
 .@R_s5_�� mo�����*�<� N�`�r�������gȍ ޏ����&�8�J�\� n�������c��џ ���"�4�F�X�j�|� ������į֯����� �0�B�T�f�x����� ����ҿ�������ٟ #�M��tφϘϪϼ� ��������(�:�L� �p߂ߔߦ߸����� �� ��$�6�H��� +�=ϟ�a��������� � �2�D�V�h�z��� ��]���������
 .@Rdv����k�}�����$F�MR2_GRP �1���� �C4  �B��	 ��x9K6F@ ay@�6G�  ��Fg�fC�8R<�y?�  ���66�X���8�75t��5��ߛ5`+�yA�3  /+BH�w�-%@S339%�5[/l-6@6!�/x l/�/�/�/�/?�/&? ?J?5?G?�?k?�?���_CFG �TK�?�? OO�9�NO 
�F0FA K@�<RM�_CHKTYP  ��$&� �ROMa@_MIN\g@�����@�R ]XSSB�3�� 7��O���C�O�O�5TP�_DEF_OW � ��$WIR�COMf@_�$G�ENOVRD_DeO�F��E]TH�֊D dbUdKT_E�NB7_ KPRA�VC��G�@ �Y�O�_�?oyqo&oI* �Q�OU�NA8IRI<�@���oGo�o�o�o��C�p3��O:��B�+sL�i�O�PSMT��Y(�@�
t�$HOSTC��21��@�\5 MC��R{����  2�7.00�1�  e�]�o������� K�ď֏���������	anonymous!�O�a�s����� �4������ ��D�!�3�E�W�i��� ������ï柀�.�� �/�A�S���课�П ����Ŀ����+� r�O�a�sυϗϺ�� �������'�n��� �����ϓ�ڿ������ ����F�#�5�G�Y�k� ���υ���������� B�T�f�C�z�g��ߋ� �����������	 -P�����u��� ���(�:�<)p� M_q������ ��/$ZlI/[/ m//�/����// �/D!?3?E?W?/? �?�?�?�?�/�?./O O/OAOSO�/�/�/�/ �?�O?�O�O__+_ r?O_a_s_�_�_�O�? O�_�_oo'o�t�q�ENT 1�hk� P!�_no  �p\o�o�o�o�o�o �o�o�o:_" �F�j���� �%��I��m�0��� T�f�Ǐ��돮��ҏ 3���,�i�X���P��� t�՟��៼�
�/�� S��w�:���^�������������ܯ=� �?QUICC0J�&��!192.16?8.1.10c�X�A1��v�8��\�2��ƿؿ9�!ROUgTER:��!���a��PCJOG|��e�!* ���0��U�CAMPRT�϶�!������RTS���x� !�Softwar�e Operat�or Panel�U߇���7kNAME� !Kj!RO�BO����S_CF�G 1�Ki ��Auto�-started^�DFTP�Oa� �O�_���O�������� ��E_�.�@�R�u�c� 	�����������cN:� L�^�;r���R�� ������% H�[m��� jO|O�O�O4!/hE/ W/i/{/�/T�/�/�/ �/�//�//?A?S?e? w?�?����??�? </O+O=OOO?sO�O �O�O�O�?`O�O__ '_9_K_�?�?�?�?�O �_�?�_�_�_o#o�O GoYoko}o�o�_4o�o �o�o�of_x_�_ g�o��_���� �o��-�?�Q�tu� �������Ϗ�(: L^`�2��q����� ������ݟ���%� H�ʟ[�m�������� ��� �ί4�!�h�E� W�i�{���T���ÿտ �
�Ϟ�/�A�S�e��w����_ERR ���ڇϗ�PDU�SIZ  �^�6����>��WR�D ?(���� � guest���+�=�O��a���SCD_GR�OUP 3�(� u,�"�IFT��w$PA��OMP��w ��_SH�޻ED�� $C��C�OM��TTP_A�UTH 1���� <!iPen�danm�x�#�+!�KAREL:*8x���KC�������VISION SET��(�����?�-�W�R���v� �����������������G�CTRL �Ҧ�a�
��FFF9E3���FRS:DE�FAULT��FANUC We�b Server �
tdG����/�� 2DV��WR�_CONFIG ����������IDL_CP�U_PC� �B����� BH�M�IN����GNR_IO������Ȱ�HMI_EDIT� ���
 ($ /C/��2/k/V/�/z/ �/�/�/�/�/?�/1? ?U?@?y?d?�?�?./ �?�?�?�?OO?OQO <OuO`O�O�O�O�O�O��O�O__;_�NP�T_SIM_DO��*NSTAL�_SCRN� ��\UQTPMODN�TOL�Wl[�RT�YbX�qV�K�EN�B�W�ӭOLN/K 1�����o�%o7oIo[omoo�RM/ASTE��Y%�OSLAVE ���ϮeRAMCA�CHE�o�ROM�O�_CFG�o�S�cU�O'��bCMT_�OP�  "��5sYC�L�ou� _ASG� 1����
  �o������� "�4�F�X�j�|����k�wrNUM����
��bIP�o�gRTR�Y_CN@uQ_�UPD��a��� �bp�b��n��M���аP}T?��k ��._������ɟ ۟퟈S���)�;�M� _�q� �������˯ݯ �~��%�7�I�[�m� �������ǿٿ��� ��!�3�E�W�i�{�
� �ϱ��������ψϚ� /�A�S�e�w߉�߭� ����������+�=� O�a�s���&���� ��������9�K�]� o�����"��������� ������GYk} ��0���� �CUgy�� ,>���	//-/ �Q/c/u/�/�/�/:/ �/�/�/??)?�/�/ _?q?�?�?�?�?H?�? �?OO%O7O�?[OmO O�O�O�ODOVO�O�O _!_3_E_�Oi_{_�_ �_�_�_R_�_�_oo /oAo�_�_wo�o�o�o �o�o`o�o+= O�os����� \n��'�9�K�]� ���������ɏۏi��c�_MEMBER�S 2�:��   $:� ���v���1����RCA_ACC� 2���   [�ߚ ��:l�6�����  ��  ����������3�� �a�BUF001� 2�n�= ���u0  u0�����
�
�)�
�7
�F
�T
�cz
�q�  pPP�YJ�� *J�8J�UGJ�UJ�dJ�rJ�U�J��J��J��J�U�J��J��J��J����ڤڤ�ڤ,ڤ9ڤIڤVRڤeڤ�������������Ȫڤ�ڤ�ڤ���M�n�j�j�i��)�1�9�A�Upj�}j��j��j�{�H��H����	��ߙ2����� �����!��)� �1��9��A��I� �P�R�X�U�"�h�U� q�U�y�U�U�U� ��U�U¡�U©�U� ��U¹�U���U�ɠU� ѠU�٠������� ����������	��� ������(��ª� 8��º�H���Q���Y� ��a���i��p�u�y� uҁ�u�rĐ�u�:Ġ� u�Jİ�uҹ�u���u� ɰu�Ѱұر���ߙ3�����l��� �!�/��1�?��A� O�l�]�`�l�+�h�w� l�y���l�����l��� ��l�����l�����l� ɢ��l�٢�Ú���� ����Ӛ�	�Ӛ�� 'Ӛ���0�?Ӛ���H� WӚ�Y�gӚ�i�w�~� y���~�{䐳��~�K� ����~���~�ɲ����ٲ����d�CFGw 2�n� 4��Tl�l�<l�4�7��HIS钜�n� �� 2025-12-�l� ��5�� �����!3�l�[~�qq1-�3]�   �# &f  �' "7��  Te�7 X�`�hl�|O�l�$  x {��8 �l�;  ��   7 �����9 ��9, ���  !  8��� d�q4[}�RM29}	�R/d/�v/�/�/�/�/�-(� %   � -�R  *g_��,B��=/*?<? N?`?r?�?�?�?�?�? ??OO&O8OJO\O nO�O�O�O�?�?�O�O �O_"_4_F_X_j_|_ �O�O�_�_�_�_�_o o0oBoTo�O��[m
7d_o�o�o�o �o!3EWEW8 cm8��� ���c��b��b�_+  X� ��X�"�!c�,�: J�"�0 � Q�1 
 R� " : b(: �q%/7/m���������Ǐُ��(5�c 2�� ,�� 1  \�_�_I�[�m�� ������ǟٟ럑_4� !�3�E�W�i�{����� ��ï���Я��/� A�S�e�w�����ү� �������+�=�O� a�s�aoN�Ѐo�o
3��������0�B�@T�f�x�fxe
��m�����ߧ�ҵ@�ҽ���������G���� 2�	��������"J� .�� Z� �� J�\���������������*T�[�6��  �澿пr��������� ������K�]�J \n������ �#5"4FXj |������ //0/B/T/f/x/�/��/��_I_CFG� 2��� H�
Cycle T�ime�Bus=y�Idl�"��min�+1�Up�&�Re�ad�'Dow�8?F� 1�#Co�unt�	Num	 �"����<��>�qaPROG�"힦����)/�softpart�/genlink�?current�=menupage,1133,�g�OO&O8O<b5leS�DT_ISOLCW  ����p�/�J23_DSP_�ENB(�vK0�@INC ��M�ӄ@�A   ?�=�?��<#�
�A�I:�o&��N_��X�O<_�GOB�0C�C�"�1�FVQG_GR�OUP 1�vK�r<��C���_D_?���?�_��Q�_o.o@o�_dovoȈo�o��,_NYG_IN_AUTO �>�MPOSRE^_pV�KANJI_MA�SK v�HqREL?MON ��˔?��y_ox����(�.6r�3��7�C����u�o�DKCL_�L�`NUM(��E�YLOGGING� ����Q�E�0LA�NGUAGE ���~��DEFAULT ��6��LG�!��:2k��3�80�H  ���'�� _ � 
��ћ���GOUF ;��
~��(UT1:%�� � �-�?�Q�h� u���������ϟ����(g4�8i�N_DISP ��O�8�_�_��LOCT3OL����Dz<�A��A��GBOOK ���d�1
�
�۠������#�5��G�Y�i���3{�W�	��쉞QQJ¿Կ1���_BUFF ;2�vK ��Ё25
�ڢVB&�7� Collaborativ�=�O� �ώϠϲ��������� '��0�]�T�fߓߊ�����DCS � �9�B�Ax���Rh�%��-�?�Q���IO 2��� ���Q��������� ����*�<�N�b�r� ���������������&:e�ER_ITMsNd�o��� ����#5G Yk}�����p����hSEV�`��MdTYPsN��c/u/�/
-�aRS�T5���SCRN__FL 2�s��0����/??1?C?U?�g?�/TPK�sOR">��NGNAM�D���~�N�UPS_AC�R� �4DIGI��8+)U_LOA�D[PG %�:%�T_NOVIC�Et?��MAXUA�LRM2��a���2�E
ZB�1_P�5�`� ��y�Z@CY���˭�O+���ۡ�D|PPw 2�˫ �Uf	R/_
_C_._g_y_ \_�_�_�_�_�_�_�_ oo?oQo4ouo`o�o |o�o�o�o�o�o) M8qTf�� �����%��I� ,�>��j�����Ǐُ �����!���W�B� {�f�������՟���� ܟ�/��S�>�w��� l�����ѯ��Ư�� +��O�a�D���p����RHDBGDEF ���E�ѱO��_L?DXDISA�0�;�c�MEMO_AP޻0E ?�;
 ױ��3�E�W�i��{ύϟϱ�Z@FRQ_CFG ��Gm۳A ��@�����<��d%�� ���t���B��K���*i�/k� **:tҔ�g�y�� ���߱��������� �J�Es�J d������,(H���[� ����@�'�Q�v�]� ���������������*NPJISC 31��9Z� ���� ��ܿ�����	Z�l_MSTR ��#-,SCD 1�"͠{��� �����//A/ ,/e/P/�/t/�/�/�/ �/�/?�/+??O?:? L?�?p?�?�?�?�?�? �?O'OOKO6OoOZO �O~O�O�O�O�O�O_ �O5_ _Y_D_i_�_z_ �_�_�_�_�_�_o
o oUo@oyodo�o�o�o �o�o�o�o?*�cN�MK���;љ$MLT�ARM���N��r ��հ��>İMETPU��zr���CNDSP?_ADCOL%�ٰ�0�CMNTF� �9�FNb�f�7�FS�TLI��x�4 �;ڎ�s����9�_POSCF��q��PRPMe��STvD�1�; 4�#�
v��qv����� r��������̟ޟ � ��V�8�J���n����¯�������9�SI�NG_CHK  }��$MODA����t�{�~2�DE�V 	�	M�C:f�HSIZE���zp�2�TASK� %�%$12�3456789 �ӿ�0�TRIG ;1�; lĵ��2ϻ�!�bϻ�YP蠱��H�1�EM_�INF 1�N��`)AT&F�V0E0g���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ��2�ԁH6�^���Rφ��A��߶�q��������  ��5������ߏ�B� ������������1� C�*�g��,��P�b� t������R�?�� �u0������ ���������M q ���Z���/ �%/��[/ 2 �/�/h�//�/�/� 3?�/W?>?{?�?@/�? d/v/�/�/O�//OAO x?eO?�ODO�O�O�O|�O_�NITORÀ�G ?z�   	EXEC1~s�&R2,X3,X4,X5�,X��.V7,X8,X9~s'R�2�T+R�T7R �TCR�TOR�T[R�TgR��TsR�TR�T�R�S2��X2�X2�X2�X2��X2�X2�X2�X2��X2h3�X3�X3�7R2�R_GRP_�SV 1��� �(꡾� �>��ˈ�F�y����c��@,3�da���_D�B��~�cION_DB<���@�zq  �Jzp�zp�Y�1u�zp͆>w�$�E�M�Y��@N   J(�rp)>|�〛Y�-ud1������8�PG_JOG S�ʏ�{
�2��:�o�=���?����0� B��~\�n������`��H�?��C�@�ŏ8׏���  ������qL_NAME� !ĵ8��!�Default� Persona�lity (fr?om FD)qp0��RMK_ENON�LY�_�R2�a �1�L�XL��8�gpl d ����şן����� 1�C�U�g�y������� ��ӯ���	����
� <�N�`�r���������8̿޿� :�� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� ��������������+��<�Sew ����������A�a�� B�Bw��Pf� �����/!/3/ E/W/i/{/�/�/�/� ��/�/??/?A?S? e?w?�?�?�?�?�?�? �?�/�/+O=OOOaOsO �O�O�O�O�O�O�O_�_'_9_&O�S���x_�]�rdtS���_ �]�_�_�W�����S"ope_oXoa �� qogoyo�o�o�o�o�o�uP�p"|����	�`[oUgy8qK�A�\����s� A� ��y@h�Q�Q��"����Tk\$�_�  ��P�P�E�xC�  � I�@oa�<o��p��������ߏ
f�Q*������0��PCr� �� 3r �.� @oD�  A�?�G��-�?.I�.@I��A����  ;��	lY�	 ��X  ������� �, � �����uP�K�o�����]�K��K]�/K	�.��w�r_x	����@
�)��b�1�����I��Y�����T;f�Y�{S���3�	���I�>J���;Î?v�>��=@�O����E��Rѯ�עZ���wp��u�� kD!�3��7p�g  �  ��9�͏W���	'�� � u�I� �  ��u���:�È��È�=��ͱ���@��ǰ�3��\�3��E�&���N�pC�  'Y�&�Z�i�b�1@f�i�n�C���¢I�C����b���r����ڟ.�B �p�Ŕq���}ر�.DzƏ<ߛ�`�K�p�ܖ����������А 4�P����.z��d � �Pؠ?��ff�_��	�� 2p>�P���8.f�t�C>L���U���(.��P���٨���������� x��;e��m��KZ;�=�g;�4�<<a����%�G��3�|���p?fff?ذ�?&S���@=0e�?��q�+�r N�Z���I���G���7� ��(�����!E0 iT����+��F�p���#�� D��w��� ����//=/(/ a/L/�/p/��/�p� 6�/Z#?�/ ?Y?k? }?��?�?>?�?�?�? �?�?1O�����KD�y�^KCO�OO�O��ɃذO�O�O�Oai����J��}�DD1���.�D��@�AmQa���9N,ȴA;��^@��T@|j�@$�?�V��>�z�ý���=#�
>\�)?��
=�G}�-]�{=����,��C+�ןBp���P��6���C98R����?N@��(���5-]G�p��Gsb�F�}��G�>.E�V�D�Kn����I�� F�W��E��'E����D��;n����I��`E����G��cE�vmD���-_�oQ_ �o�o�o �o$H 3X~i���� �����D�/�h� S���w��������я 
���.��R�=�v�a� s�����П����ߟ� �(�N�9�r�]����� ����ޯɯۯ���8� #�\�G���k������� ڿſ���"��F�1� C�|�gϠϋ��ϯ����������P(�Q343�] �����Q�	�x9�Oߵ53~�mm��aҀ5Q�߫�a�Ǔ����ߵ1��������1��U�C�(y�g��%P�P���!�/��'���
���.������4�;�t� _��������������� :%��/�/d������� �7%[I�m���027� � B�S@J@�CH#PzS@�0@ZO/1/@C/U/g/y/�-�#���/�/�/�/�/�3?��3�� @�3��0�0�13��5
 ?f?x?�?�? �?�?�?�?�?OO,Op>OPO�Z@1 �������c/�$MR�_CABLE 2�ƕ� ��TT�����ڰO���O �)�@���C_���_ O_u_7_I__�_�_�_ �_�_o�_�_oKoqo 3oEo{o�o�o�o�o�o �o�o�oGm/�K!�"���O�����ذ�$�6����*Y�** �COM� ȖI�����:0� ��G%�% 234567O8901���� ��HÏ��� � !� ��!
���M�not sent� b��W���TESTFECS�ALGR  egD�*!d[�41�
k�������$pB����������� 9U�D1:\main�tenances�.xmlğ�  �C:�DEF�AULT�,�BGR�P 2�z�  嬓 ,��%  ��%!1st cl�eaning o�f cont. �v�ilatio�n 56��ڧ�!0�����+B��*�`����+��"%���mech��cal� check1�  �k�0u�|��ԯ����Ϳ߿��@���rollerS�e�w�ū��m���ϣϵ�@�Bas�ic quarterly�*�<�ƪ,\�)�;�M�_�q�8�cMJ��ߓ "8��!� ���ߕ ��� ��+�=��C�g��ߋ�ʦ�߹���������@�Overghau�ߔ��?�C x� I�P����@}���������� $n� ������)l�ASe w������ � +=O�s� ������/R �9/�(/��/�/�/ �/�//�/�/N/#?r/ G?Y?k?}?�?�/�?? ?�?8?OO1OCOUO �?yO�?�?�O�?�O�O �O	__jO?_�O�Ou_ �O�_�_�_�_�_0_o T_f_;o�__oqo�o�o �o�_�oo,oPo% 7I[m�o��o�o ����!�3�� W��������ÏՏ �6����l����e� w���������џ�2� �V�+�=�O�a�s� �����ͯ���� '�9���]�������� ��ɿۿ���N�#�r� ��YϨ�}Ϗϡϳ��� ���8�J��n�C�U� g�yߋ��ϯ������ 4�	��-�?�Q��u� �����ߞ�������� �f�;�������� ���������P��� t�I[m���� ��:!3E W�{��� � ��//lA/�� w/��/�/�/�/�/X*�"	 X�/?.?@?�)B a/o?m/o%w? �?�?}?�?�?OO�? �?OOaOsO1OCO�O�O �O�O�O__'_�O�O ]_o_�_?_Q_�_�_�_��_�_�\ Џ!?�  @�!  M?HoZolo�&4o�o�oܽo�(*�o** F�@ �Q�V�` o'9�o]o�����/^&�o� ����/�A�S�e� ��#�����я��� ��+�q�����7��� ����k�͟ߟ��I� [���K�]�o���C������ɯ��o$�!��$MR_HIST� 2��U#�� �
 \7"$ 23�45678901P3�;���b2�90/ ����[���./���� ǿٿF�X�j�!�3ρ� ����{��ϟ����� B���f�x�/ߜ�S��� �߉��߭��,���P��t��=��$�S�KCFMAP  ]�U&��b�
�� ����ON?REL  �$#�������EXCFE�NB�
����&�F�NC-��JOGO/VLIM�d#�v���KEY�y���_PAN������RUNi�y����SFSPDTY�PM����SIGN|��T1MOTk�����_CE_G�RP 1��U ��+�0�ow�#d� �����& �6\�7y� m���/�4/F/ -/j/!/t/�/�/�/{/��/�/�/?�+��QZ_EDIT
�����TCOM_CFG 1���0�}?�?��? 
^1SI 	�N����?�?��!�?$O����?XO~78T_ARC_*��X�T_MN_oMODE
�U:�_SPL{O;�UA�P_CPL�O<�N�OCHECK ?��� ��  _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo���NO_WAITc_L	S7> NTf1�����%��qa_7ERRH2��������?o�o�o�o��POGj�@O�cӦm�| ��:GA����EA�mm�2�&����K��wC����<���?���)��|�n�bPARAM�b]����tGO��8
�.�@� =  n�]�o�w�Q������� ����Ϗ�)��7��[�m� �����ODRDSP�C8��OFFSET_C�ARI0�OǖDIS�ԟœS_A�@AR�K
T9OPEN_FILE��1T6��0OPTION_�IO����K�M_P�RG %��%$�*����'�WO�-�Ns�ǥ� ��5�9���	 �������>d���RG�_DSBL  �����jN���RI_ENTTO���C�����A ��U^�@IM_DS����r��V��LCT �{mP2ڢ�3̹���d��%���_PEqX�@���RAT�G� d8��̐UP� װ�:����`S�e�Kωϗ��$�r�2G�L�XLwȚ�l� ��������'�9�K� ]�o߁ߓߥ߷����߀�����#�5�G���2 ��v�������������e�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?�q1�~?�?�?�?�? �?�?�?O O2ODO�yA�a�tn?~M��~O�O�P�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�O�Oo $o6oHoZolo~o�o�o �o�o�o�o�o �_ oVhz���� ���
��.�@�R�0d�QOES������
B�d�ӏ�ʏ� �������Y�D�}�0��r���������ԟ ڟ���p���=�M��q�	`��������c�:�o�¯ԯ�����A�  P�k�C�C�ڰ"ڰ����O��/  ���-���~)�C�  �t� k���g�����Կ��ѿ�
�5���_:�ĳ�OU����A��A��H��n�� o� ^�\�� @D�  p�?��v�\�?:px�:qC�4r�p�(��  ;��	l��	 ��X  ������� �,? � ��������Hʪ�����H���Hw�_zH�����8�B���B�  �Xѐ�`�o�*��3�	���t�>u���fC{�����:pB\�
��Ѵ9:qK�t�� ����$����*��� DP��^��b�g  �  �h������)�	'� � ���I� � � ��'�=��q�����t�@��@��!�b��^;b�t��U�(�N��r�  '���E�C�И�t�C��И��ߗ���jA�@!�����%�B�� ���,���H:qDz �k�ߏz���w�����А 4P��D�:uz:���	f�~�?�ff'�&8� ]�mb�8:p��>L��H���$�(:p�P���	������:� �x�;e�m"��KZ;�=g;�?4�<<���E/�Tv��b���?offf?�?&� �)�@=0�%?��%_9��}!��$� x��/v��/f'��W,? ?P?;?t?_?�?�?�? �?�?�?O�?(OOLO �/�/�/EO�OAO�O�O �O�O_�O_H_3_l_ W_�_{_�_�_1��_A� ��eO+o�ORooOo�o �o�oK/�o�omo�o@*'`+�,�zt���CL�H��}?�����
������u����#D1�/n�t��p�qޜ�@I�h~,���A;�^@���T@|j@$��?�V�n�z��ý��=#��
>\)?���
=�G�����{=��,���C+��Bp�����6��C98R���?}p���(��5���G�p�Gsb��F�}�G�>�.E�VD�K�L����I��� F�W�E���'E���D���;L����I���`E�G���cE�vmD���\�՟��ҟ���/� �S�>�w�b������� ѯ�������=�(� :�s�^���������߿ ʿ�� �9�$�]�H� ��lϥϐϢ������� ��#��G�2�W�}�h� �ߌ��߰�������� 
�C�.�g�R��v�� �������	���-�� Q�<�u�`�r������� ������'M�=(�34�]O!����8h~�%3�~�m����5qQ������<�!���  �`N�r��	eP@"P��Q�_/V�/9/$/]/H)����c/j/�/�/�/�/�/ �/�/!??E?0?i?T?�"&�_�_�?�?�8� �?�?O�?OBO0OfO TO�OxO�O�O�O�Oy2f?_  B��p,yp$QCHR�z�p@�N_`_r_�_�_�_�]c�O�_�_oo�+o?�Bc� @*d4�QqJc�D
 2o �o�o�o�o�o�o %7I[m��oa� �����c/��$PARAM_MENU ? ��  �DEFPU�LSE��	WAITTMOUT�{�RCV� �SHELL_WR�K.$CUR_S�TYL�p"�OsPT8Q8�PTBM��G�C�R_DECSN�p��������� �����-�(�:�L��u�p��������qSS�REL_ID  ���̕USE�_PROG %��z%���͓CCR��pޒ��s1�_HO�ST !�z!6�s�+�T�=���V��h���˯*�_TI�ME�rޖF��pGDEBUGܐ�{͓�GINP_FLM3SK��#�TR2�#�WPGAP� ��_�b�CH1�"�TYPE�|�P����� ���0�Y�T�f�x� �ϜϮ���������� 1�,�>�P�y�t߆ߘ� �߼�����	���(��Q�L�^�p��%�WO�RD ?	�{
 �	PR�p#�MAI��q"SU�d���TE��p#��	91���COLn%��!���L�� !���F�d�TRA�CECTL 1�v �q �_� �#��|��_�DT Q� ���z�D � ��^a�� ��c`���������� 1CUgy�� �����	- ?Qcu���� ���//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?�?�?�?�? O!O3OEOWOiO{O�O��O�O�O�O�G� �@�P�BM`�Bk` �B���O�O�ON_`_r_ �_�_�_�_�_�Y��
U oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n��� ������"�4� F�X�j�|�������ď ֏�����0�B�T� f�x���������ҟ� ����,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� .�oP�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/Dϒ/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z�����������$PG�TRACELEN�  ��  �_����Ά�_UP ������������΁_CFG M���烸�
���*�:�D�O���O��  �O��D�EFSPD ܲ������΀H�_CONFIG s���� �����dĔ�݂ ���ǑP^�a�㑹���΀IN�TRL' ��=�8^����PE��೗����*�ÑO�΀LI�D���	T�LL�B 1ⳙ k��BӐB4��O� 䘼�����Q� << ��?������� M�3�U���i����������ӿ��	�7�T� Ϣk�b�tϡ�诚���������S�GRP �1爬���@A!���4I����A �Cu��C�OCjVF
�/��Ȕa�zي�ÑÐ�t��ޯs�F��´�ӿߨ�B�� ���������A�S�&�B34�_�0������j��� ������	�B�-����Q���M�������  Dz����.����� &L7p[�� �����6!�Zh)w
V7�.10beta1�*�Ɛ@�*��@�) @�+�A Ē?��
�?fff>���~�B33A�Q��0�B(��A�?��AK��h� ���//'/9/P�p*�W�ӑ�n/�/��%���R�fh����*���P 2�LR��/�/�/�/�/HH?�Ĕ�I�u� &:���?��x?�?A����P!\3 Bu�B�L�?�5BH�3[4��1o��4��[45�)�/B\3x3Dx�?YO �?aOkO}O�<<�R @��O�C�O�O�O�O�D�A�X�KNOW_M�  Z�%�X�SV7 賚ڒ�� �_�_�_?�_�_�_Po����W�M+�鳛� ��	@�3#���_�o�\A���
]bV4�@u��u��e�o�l,�VX�MR+��JmT3?���W�1C{�OAD?BANFWDL_V�{ST+�1 1����P4C���[� �i/�����?� 1�C���g�y������� �ӏ�*�	��`�?�Q�c��w2�|Va�upG�<ʟ���p3��Ɵ؟Ꟃw4��+�=��w5Z�l�~����wA6����ѯ㯂w7 ��$�6��w8S�e�w�����wMAmp�������OVLD  ���yo߄rPARNUM  �{p+þ�?υqSCH�� �
��X���{s��UPDX�)ź���>��_CMP_@`��̑p|P'yu�ER�_CHK���`yqbb3��.�RSp�p?Q_MOm��_�}ߥ�_RES_G
�p쩻
�e����� 0�#�T�G�x�k�}�� �������������׳���������:�Y� ^���Y�y������Ӭ� ������������ ��R�6UZ�ӥ�ux����V 1�F|vpVa@k�p��THR_INRp���(byudMASmS Z)MN�GMON_QUEUE �uyvup�\!��N�UZ�N8W��END��ߎ�EXE����B�E���OPTI�O��ۚPROG�RAM %z%���~ϘTAS�K_I��.OCFG �z+�n/� �DATACc�+�@ '9up? 2 �??`/?A?S?]51 s? �?�?�?�?�6p1�?�?��?O"O,F�!INFOCc��-��bdlO ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_��_�_�_�_�/A@FD���, 	��!��K_Ƥ!�)fN!fEN!B��0m��Pf2Yokh�G�!2�0k X�,		d�=��M·o���e�a$�p�d��i�i�g_EDIT ��/%7�����*SYST�EM*upV9.4�0107 cr7/�23/2021 �A��Pw��PRGADJ_p  h $X[Ѿp $Y�xZ��xW�xқtZқtS�PEED_�p�p�$NEXT_CYwCLE�p �q��FG�p �~�pALGO_V ��pNYQ_FR�EQ�WIN_T�YP�q)�SIZ:1�O�LAP�r!��[��M+����qCR�EATED�r�IsFY�r@!NAM�p�%h�_GJ�ST�ATU��J�DEB�UG�rMAILTuI����EVEU��LAST�����t�ELEM� � $ENAB�r�N�EASI򁼁AwXIS�p$P߄�����qROT_sRA" �rMAX �ԞqE��LC�AB�
���C D_LVՁ`�BAS��`�1��{���_� ��$,x���RM� RB�;��DIS����X_SqPo�΁�� ��t|�P� | 	�� 2 \�AN�� �;����8�Ӓ�� �0�PAYLO��3�V�_DOU�qS���p��tPREF� �( $GRID*�E
���R���uY����OTOƀ>�q  �p��q!�p��k�OXY� � $L��_PO|�נVa�SRV��)���DIRECT_1�� �2(�3(�4(�5*(�6(�7(�8����F��A�� $�VALu�GRO3UP��� ���_� !���@!�������RAN泲���R��/���TOTA��F���PW�I=!%�REGEN#�8����� ��/���ڶnTzЉ���#�_S����8�(��V[�'���4���GRE��w���H��D������V_H��DAY:3�V��S_Y�Œ~;�SUMMAR���2 $CON?FIG_SEȃ����ʅ_RUN�m�C|�С�$CMPR��P�DEV���_�I�ZP�*��q��ENHANCE�	�
���1���'INT��qM)b�q��2K����OVR6o�PGu�IX��;����OVCT����qF>u�
 4 ����|a˟��PSLG"�>� \ �;��?�1���SƁϕc�U�����Ò��4�U��]�Tp�G (`�-��rJ<��O� CK�IL_M�J���VN�+��TQ�n{�N5���C�U�LȀD�V(�C6�P�_�຀@�MW�V1VV�V1d�2s�2d�U3s�3d�4s�4d� �'�	�������p	�{IN	VIB1qp�1� 2!pq/,3* 3,4 4,�p ?��;��A���N��������PL��TO�Rr3�	��[�S{AV��d�MC_FOLD ?	$SL�����M,�I��L�� �pL�b��KE�EP_HNADD�	!Ke�UCCOMc�k��
�lOP���pl\��lREM�k���΢���U��enkHPW� K�SBM��ŠCOLLAB|�Ӱn��n��+�IT�O���$NOL�FCALX� �DON�r�p��� ,��FL|���$SYN�y,M�C=����U_P_DLY�qs"�DELA� ����Y�(�AD��$TA�BTP_R�#���QSKIPj% ����OR� �E�� P_��� �)�� �p7��%9��%9A�$: N�$:[�$:h�$:u�$:t��$:9�q�RA��� X�����M}B�NFLIC]���0"�U!�o���NO�_H� �\�< _S�WITCHk�RA_PARAMG�O ��p��U���WJ��:Cӣ�NGRLT� OO�U���p��X�<A��T_Ja1�F�rAPS�WEI{GH]�J4CH��aDOR��aD��OO��)�2�_FJװ���saA�AV��C�HOB.��.�`�J2�0�q�$�EX��T$�'QIT��'Q�pG'Q-�GΨ�RDC�m" G� ��<��
R]���
H���RGEAp��4��U�FLG`�g��H��ER	�SsPC6R�rUM_'P>��2TH2No��@�Q 1  ���0����  �D �وIi�2_P�25cS�ᰁ+�_L10_CI��pe� �pk�� ��UՖD��zaxT�p�Q(�;a��c���޲+�i���e��`� P`DESIG\Rb$�VL1:i1Gf��c�g10�_DS���D�Xp
`FPOS;11�q l�pr0��x1C/#AT�B���U
WusIND ��}�mqCp�mq`B	��HOME�r��?t2GrM_q����!@s3Gr���X ��$� >u4GrG�Y�k�}�����`!
@s5Grď֏���(����6GrA�S�0e�w����� @Ar7Gr��П�����6�8Gr;�M�_��q�����*�S �q ` �@sM��PQ�<K@��! T`M�L�M�IO��m�I��:2�OK _OPy���x »Q�cPOWE�" 7�x EQ:AE � #s%Ȳ�$DSBo�GNAH�b� C�P2�)WQ�S232S�$ ��iP��xc�ICE�<@%�PE`2� @I9T��P�OPB7 1�oFLOW�TRa@42��U$�CUN��`��AUXT��2Ѷ�EORFAC3İUU��	�CH��% t<_9�EЎA�$FREEFROMЦ�A�PX qЎUPD"YbA�PT.�pEEX0���Í!�FA%b�5���RV�aG� & W C�E�" 1�AL�  �+�jc'���D�  2& ��S\PcP(
  �$7P�%�R�2SP���T�`AXU���DSP���@�W���:`$��RNP�%�@����=K��_MIR����f�MT��AP�`��P"�qD�QSYz�������QPG7�BR�KH���ƅ AXI�  ^��i����1 ����BSOC����N��DUMM�Y16�1$SV�DE��I�FSP_D_OVR79�2 D����OR��֠�N"`��F_����@O�V��SF�RUN���"F0�����UF�"@G�TOd�LCH|�"�%RECOV��9@�@W�`&�ӂH���:`_0�  @>�RTINVE��ѡ�OFS��CK�KbFWD������1B喻�TR�a�B �FAD� ��1= B1pBL� �6� A1L�V��Kb����#��@+<�AM:��0��j��_M@ ~�@h����T$X`x ��T$HBK���F��A�S����PPA �
��	������?DVC_DB�3@@pA�A"��X1`�X3`��Se@�`��0��Uꣳ�h�CABPP
R�S #��c�B�@���GUBCP	U�"��S�P�`R���11)ARŲ�!$HW_CGpl�11�� F&A1Ԡ@8p�_$UNITr�l >e ATTRIr@y"���CYC#b�CA���FLTR_2_FI������2b�P��CHK_��S�CT��F_e'F_o,�"�*FS�Jj"CHA�Q�'91Is�82RSD����1���_Tg�`� �i�EM�NPMf�T�&2 8p&2- �6D�IAGpERAIL�ACNTBMw�LOh@�Q��7��PS��b� � ��PRB)SZ`�`BC4&�]	��FUN5s��RIN�PZaߠ�07DFh�RAH@���`� �`C�@�`C�Q�CBOLCURuH�DA�K�!�H�HDAp�aA�H�C�ELD������Cd��jA�1�CTIB�Uu�8p$CE_gRIA�QJ�AF �P�>S�`DUT2b�0C��};OI0DF_LC�H����k�LMLF�aHRgDYO���RG�@�HZ0��ߠ�@�UMUGLSE�P�'3iB$J��J����FAN_ALM�d�bWRNeHAR�D��ƽ�P��k@2�aN�r�J�_}�A�UJ R+4�TO_SBR��~b�Іje �6?A�cMPINF´�{!�d�A�cRE�G�NV��ɣZ�D���NFLW%6r$M�@� ��f� �0� h'uCM4NF�!�ON	 e!e#�p(b*r3F�3 �	 ����q)5�$�3$Y�r�� u�_Ѿ�p*$ �/�EaGE�����qAR�Єi���2�3�u�@<�A�XE��ROB��R�ED��WR��c�_���SY`��q� ?�SI�WRI���vE �STհ�ӭ d���Eg!���t8��^a�БB����9�3� O�TO�a����AR�Y��ǂ�1�����F�IE���$LIN]K�QGTH���T_������30���XYZ���!N*�OFF����J�ˀB��,Bl�0��e���m�FI� ���C@Iû�,B��_J $�F�����S`����3-!$1�w0���R2��C��,�DU���3�P�3TUR`XS.�Ձ�bXX�� ݗFL�d���pL�0�按34���� 1�)�K��M�5��5%B'��ORQ��6��fC㘴��0B�O ;�D�,������a�'OVE��rM���� �s2��s2��r1���0�0��0�g /�AN=!� 2�DQ�q���q�}R� *��6����s��V���SER��jA	�2E��H.�C��A���0���XE�2Ӈ�A��AAX ��F��A�N!�SŴ1 _��Q_Ɇ�^ʬ�^ʴ��^��0^ʙ�^ʷ�^�1 &�^ƒP[ɒPkɒP{� �P�ɒP�ɒP�ɒP�� �P�ɒP�����ɪ �R�>�DEBU=#$�8ADc�2����
�AB��7����V� <" 
��i�q��-!�� %��׆��׬��״��� �1�י��׷�JT��DR\�m�LAB��ݥ9 FGRO� ݒ=l� B_�1�u��� }��`����ޥ��qa��AND�����qa� �Eq��1�0�A@�� �NT$`��c�VEL�1��m��1`u���QP��m�NA[w�(�CN1� ��3�����SERV9Ec�p+ $@@d@n��!��PO
�� _�0T !��򗱬p,  �$TRQ�b
�(� -DR2,�+"P�0_ . ql"@!�&ERR���"I� q���~TO	Q����L�p]�e��
�0G��%���p�RE�@ / ,h��/I -��RA�? 2. d�&s��"  0�pC$&��2tPM� ��OC�A8 1  }pCOUNT��� ��SFZ�N_CFG2 4B �f�"T�:#�0�Ӝ�  ^�s/3 ���M:0�R��qC@��/�:0�FA1P��?V�X������r���� �P�:b]HELpe�4 5��B_wBAS�cRSR�f� @�S�!QY 1T�Y 2|*3|*4|*U5|*6|*7|*8��L!RO�����NL�q �AB���0Z �ACK��INT�_uUS`�Pta9_cPU�>b%ROU��PH@�h9#�u`w�9��TPFWD_KA1R��ar RE���PqP��A]@QUE�i@&��	�f�>`QaI`���9#�j3r��f�SCEME��6��PA�7STY4SO�0�DI'1�`���18�rQ�_TM�cMANR�QXF�END��$KEYSWIT�CHj31:A�4HE�	�BEATM�3PE�pLE��1��H�U~3F�42S?DD_O_HOMBPO:a60EF��PRr��(*�v�uC�@O�Qo ��OV_Mϒ��E�q�OCM���7����
:#HK�q5# D��g�Uj�2�M�p�4R��FOR]C�cWAR�����:#OM�p 6 Q@�Ԣ�v`U|�P�pQ1�V'p�T3�V4��V ��S#O�0L�Ry7��hUNLOE0�hdEDVa  8���@d8 <pAQ�9�l1MSUPG��UaCALC_P�LANcc1��AY�S1�19c�9 � 	X`��P �q;a@�թ�w��2��j�M$P��㣒�fyt$��rSC�M�pm�q ���aq���0�tYzZzE!U�Q�b�� T!�Hr�pPv�]NPXw_ASf: 0g �ADD��$S{IZ%a$VA��~�MULTIP�"�ns�PA�Q; � $T9op�B����rS��j!C~ �vF'RIF�2S�0�Y�T�pNF[DODB�UX�B��u&�!���CMtA�Е����������lqZ ��< �3 �p�TEg���^��$SGL��T���X�&{���㰀��S�TMTe�ЃPSE�G�2��BW���S�HOW؅�1BAN�`TPO���gᣥ��Ԣ��� V�_Gv�= ��$PC��X�O�FB�QP\��SP�0A&0^�, V�DG��>� �cA00�����P����P���P���P��5���6��7��8��9��A��b`���P��w���S`��F����h����1��v�h�י1�1��1��1�1�1�%�12�1?�1L�1�Y�1f�2��2��2���2ʙ2י2�2��2��2�2�2�%�22�2?�2L�2�Y�2f�3��3��3���3ʙ3י3�3P�����3�3%�U32�3߹3L�3Y�U3f�4��4��4��U4ʙ4י4�4�U4��4�4�4%�U42�4߹4L�4Y�U4f�5��5��5��U5ʙ5י5�5�U5��5�5�5%�U52�5߹5L�5Y�U5f�6��6��6��U6ʙ6��6��6�U6��6�6(�6%�U62�6߹6L�6Y�U6f�7��7��7��U7ʙ7��7��7�U7��7�7(�7%�U72�7߹7L�7Y��7f��V�`_UP�D��? �c� 
]V���@ x $TOR�1T�  �cOP �, 6ZQ_7RE^��(� J��SsC�A���_U�p��Y�SLOA"A � �u$�v��w�@��x�@��bVALUv�10�6�F�ID�_L[C:HI5I~�R$FILE_X3�eu4$�C�P�S;AV��B hM �?E_BLCK�3�|ȁ�D_CPU���p��p5hzQPY���R3R C � PW��� 	�!;LAށSR�#\.!'$RUN�`G@% $D!'$�@G%e!$e!�'%HR03$� '$�QT�2Pa_LI�RD w � G_O�2}�0P_EDI�R�8`T2SPD�#�E�"i0ȁ�p	���DCS9@G)�F � 
$JPQC71q�� S:C;}C9$MDL73$5P>9TC�`@7�UF�@?8S� ?8C�OBu ��!|�L�G��P;;� 9�:;kqTABUI�_�!L�HGb�% sFB3G$�3�A�sR�LLB_AVAI�B�q�3�!��wI $� SEL� sNẼ�@RG_D aN��Ta���3SC�POJ �1/AB�P1T�R?�w@_M]`L��K \M f/QL_���FMj��PGi�Ut9R�6��PS_��P\� �p�EE7B��TBC2�eL ����``�`b$�!F�T�P'T�`TDCg�� BPLp�sNU;WTH��qhTgtW�R�2$�pERV�E.S�T;S�Tw�R_�ACkP MX -$�Q�`.S�T;S��PU@�`IC�`LOMW�GF1�QR2g��`��p�S�ERTIA�d^0iP�PEk�DEUe�LACEMMzCC#c�V�B�rpTf�edg�aTCV8�l�adgTRQ�l�e��j|�Scu��edcu�J7_ 4J!��Se)@qde�Q2�0����1�PRcuPJKlvV�K<�~qcQ~qw�spJ�0��q�sJJ�sJJ�sAAL�s�p�s�pȲv���r5sS�`N1@�l�p�k�`5dXA_́�PCF�BN =`M GROU ���bh�NPC0sD�R�EQUIR�R� E�BU�C�Q�6g0 �2Mz��Pd�QS�GUO�@�)AP�PR0C7@� 
$:� N��CLO� ǉ�S^U܉Se
Q�@A.�"P �$PM]P�`8�`sR�_MGa!��C���+��0�@,�B{RK*�NOLD*�SHORTMO�!Hm�Z��JWA�SP�t p`�sp`�sp`�sp`�s(p`�A��7��8sQ�0|�RTQ� m���R.Q�cQ�PATH�*� �*��X&����P�NT|@A��"p��� �IN�RU�C4`a��C�`UM��Y
`�)p��>��Q��cP���p��PA�YLOAh�J2LN& R_Am@�L ������+�R_F�2LSHR�T/�L�O���0���>���ACRL0z�p�y�ޤsR9H5b$H+����FLEX��#�JVR P��_._�_�_����US :�_�Vd`0�G��_tQ0d`�_�_lF1G��� ��o0oBoTofoxo��E�o�o�o�o�o�o�o  ����wz3lt��@��3EWF�^zT!��X�'qju��uu ~�W؁���p�u�u@�u�u���� ��(�T �P5�G�Y��' AT��l�pE�L0�_B��s�J�Svz�JEW�CTR7B�`NA��d�HAN/D_VB�����TUO@`+�`T�SW8F�A�V� $$M��e  G�AV�Qs�De�o�AA��@�	$�A(5�G�AU�Ad�� �6��G�DU�Dd�P2D�G/ -STI�54V�5Ng�DYF �� +�x����P&�G�&��A��lw�o�Q�k�P ������ʕӕܕ��9�UW 7 ��� ��3%�?!AS�YMT��m�T�Vp�o�A�t�_SH� ~������$����Ưد�J񬢐�#39\"���_VI��`8|�q0V_UNIrS�4��.�Jmu�2��2 A��4X��4�6a�pt� ������&E_������!�E��CH( X� ̱���T-Oc�PP�VsSvD�US�RU�P�����z@�D�A}@_5�U��P�EyAa��RPROG�_NA��$�$�LAST���CA�Ns�ISz@XYZ_SPu�DW]R@Ͱb,VSV@�E1QENc���DCUR�H�P��H7R_T��YtQ"9S�d��O�T���uP?�Z ��I�!A�D���Q���#�S������2�vP �[ � MEB�O��R#B�!T�PPT0F@1�a��A̰� h1a%iT0�� $DUM�MY1��$PSm_��RF��  1��lfװFLA*�Y�P�bc$GLB_TI �U�e`gA���LIF(!\����g`OW�P��e�VOL#qb �a_	2��[d2�[`����b�P�cZ`TC���$BAUDv��cS�T��B�2g`ARI{TY0sD_WAIt�AIyCJ2�OU�6�ZqyyTLAN1S�`�{S�SZc��BUF_�r�fиx��PyyCHK_�@CkES��� JO`�E�aA�x�bUBYT�����r�.��.� ��aA��M���8����Q] Xʰ��֚�ST����SB=R@M21_@��T$SV_ER�bL����CL�`��A1��O�BpPGLh0EW~(!^ 4 $a�$Uq$�q$AW�9�A�@R��tt`ӃUم_ "���D$GI��}=$ف ^҄��(!` L�.��"}�$F�"E6�NEA9R��B$F}�йTQ# �J�@R� a7�$JOINTa�)���Ձ�MSET(!b  "+�Ec�2�^�Se�' �J�_�(!c�  ھ�U�?���LOCK_FO@� �PoBGLV��GL'��TE�@XM���EMP��:�K��b��$U�؂a�2_���q�`<� �q��^��CE/�?��� �$KARb�M�ST�PDRA܀����VcECX�����IUq��av�HE�TOOiL���V��REǠ'IS3��6��A�CH̐m b^QON$e[d3���IdB�`�@$RAIL_B�OXEa���RO�B�@D�?���HOWWAR0Aa�i`-�ROLMtb��$�*����T��`����O_F�U�!��HTML58QS�� ����(!d��N@�@�(!e���������}p(!'f t��m�^a��Xt��B�PO��A	IPE�N���O�����q��AORDEaD�m �z�XT`���A)mSP�O�P �g D �`OB �����ǯ�Uc�`���� ��SYS��AD�R��pP`U@^  �h ,"��f$A���E��E�QPV�WVA�Qi �c �@ق�UPR�B>�$EDI�Ad�_VSHWRU�z�ƀ�IS�Uq�pND��P7���G�HEAD��! @���!i�KE�UqO`CP)P��JM�P��L�UN�TR�ACE�Tj����IL�S��C��N�E���TICK�!MKQ"��HNr�k @���HW�C��P�FF��`STYeB+�LO�a��Ҕ[�C�l3�
�@�F%�$A��D=��S�!$�1�p a�e�q�e9Pv �FSQU��#�LO�b_1TERC�`!�TS?�m 5���R�m@3����ܡ��O`	c IZ�d�A�eha�qtb�}�hA}pP~r��_D)O�B�X�pSSQ�S'AXI�q��v�bS��U�@TL���RE3Q_ܠ��ET���`��CY%��FY'��A,f\!\d9x�P� g�SR$$nl-�w �����c
�uV
Qh(�AA���dC`�A�@�	�Y��D���p�E"�	CC�C`��/�/�/	4VA ��SC�` o h�5�DSmడ[`SPL�@�AT� 
R��xL��XbADDR�s3$Hp� IF�Ch�O_2CH���pO��\��- �TUk�Ir7 p��CUCp*F�V��I�Rq�4����c��
K�
V8*���Pr \z�D�A���|,K� P�"C�N��*CƮ��!�T�XSCREE��s8�Pp@�INA˃<��4�D���Q9_��`t Tᫀ �b����O Y6���º�U4h�RR������дR1�T<0UE��u# �j �qz`Ś��'RSML��U����V�1tPS_��6\� �1�9G\���C��2�@4 2��0O�v�R��&F�AMTN_FL*�`Q��W�~�� �BBL_/�9WB`�Pw ����B5O ��BLE"�Cxg�R"�DRIGHt�RD��!CKGR�B`�ET���G�AWIDTHs���R	��a��r�UI��EYհRx d�ʰ�����`y�BACKЍ�tb>U���PFO܉�QWLAB�?(��PI��$UR�m�~P��P�PHy1 y 8 $�PCT_��,"�R�PRUp �s5�C�RO%!t�%zV�ȇ�pU�@�S9R ���LUM�S��� ERVJ�h�PP|��T{ � " �GE�Rh� �¯�LIPAeE��)^g@�lh�lh�ki5ik6ik7ikpP`�Z�x����$u1��p�Q� zQUSR�ل| <z��PU�2�a#2�FOO 2�P�RI*m9�[�@pT�RIPK�m�U�NDO��})�`��Yp��y����h����p ~�Rp�qG ��T���-!&�rOS2��vR��2�s�CA�����rHo�Qi�UIaCA�����3Ib_�sOFFTA�D@���Ob��r�5�L�t��GU��Ps��������+Q�SUBo� ��E/_EXE��V
�s�WO� �#���w��WAl�p΁zfP
 V_DB�H��pT�pO�V☖����3OR/�5�RAU@6�TK���y__���� |j ��OWNj�34$GSRC�0`���DA�<��_MPFI����ESP��T�$0��c��g�An�z�E!G� `%�ۂ34J�n��COP��$���p_���/�+�6����CT�Cہ�ہ��C��DCS��P;4�COMp�@�;��Oo�=����K�^�/�VT��q'���Y٤Z���2���@p�w#SAB����2�\0˰_��qM��%!]�DIC#池AY�3G�PEE2�@T�QS�VR1���"eQL�� a��P� D ��f�z��f�> ����6�Z!A�t�b# ��L2SHADOW���#ʱ_UNSC�Ad�׳OWD�˰D�GDE#LEGAyC)�q' �VC\ }C��� v����だm�RF07����7d`C2`7�DRI%Vo���ϠC�A]��(�` ���MY_UBY�d?Ĳ��s��1@��$0�����_ఴ����L��BM�A�$�DEY	�EXXp@C�/�MU��X���,��0US����;p_�R"1�0p#�2�G>PACIN*���RG��c�y�:�y��sy�C/�RE�R"!�q�sB�y�D@� L !�G�P�"��P�R�pD@�&P�Px1dQ��	.���RE���SWq�_Ar�u@$+�{�Oq�AA/�3��hEZ�U���� Yy@�HK���P�J��_/�Q0{�EAN��ۀ2�2�X���MRCVCA� ��:`ORG��Q�dR	p��L�����REFoG �����!�+`	�p ��������<���q�A_����r��� S�`�C��Ú�q�@D� ��0�!��#q�š��OU����?� ��Վ2�J@0� 1�*p����0� UL�@��C�O�0)��� NT�[��Z�Qf�af% L飏��Q|��a�VIAچ7� �ÀHD7 6P�$JO�`oB?�$Z_UPo��2Z_LOW��$�QiBn��1$EP �s�y�� 1!f� � 1¦4�� 5�PA�A ��CACH&�LO �w�ВQB����Cn�I#F^��T8m����$HO2�32!{��Uÿ2O�@����Ro��=a��ƐV�P���@A"_SIZ&�K$Z$�F(�G'��v�CMPk*FAIo�5G��AD�)/��MRE���"P'GP��0е�9�ASYNwBUFǧRTD�%��$P!�COLE_2D_4�5W�sw�~��UӍQO��%EC;CU��VEM��v<]2�VIRC�!5�#�2�!_>�*&�pWp���AG	9R�XYZ@�3�W���8���4+Qz0T"��IM�16�2P�GRA�BB�q��;�LERrD�C ;�F_D��F�f50MH�PE�R���0�����JRL�AS�@��[_GEb� �H൑~23�ET����"���b���I�D�ҙ6m�BG_gLEVnQ{�PK|�X�6\q��GI�@N\P�4����P��!g�$dr�S� �NRT�	Lʁc�Ų��#a�4�c"!D�qDE�����Xа�X��	 ���2��d��p�zZ���d�c���DR4qȾ�2pT��U&��� $�ITPr�9p[Q��ՓV�VSF$�d�  fp/�ff�UR����SMZus�dr��ADJ`�C�� ZDVf� D�XAL� � 4 �PERIKB$MoSG_Q3$Q! o%[���p'��dr:g�qQ� �XVR2\t��B�pT_\��R��ZABC"�����Sr���
��aA�CTVS' � � $|u�0�c�CTIV�Q!IO0u¥s&D�IT�x�DVϐ
x�P��i�!���pPS���� �#��!���q!LSTD�!�  �_ST��a�aq�;CHx�� L-�@���u�Ɛ*���P G�NA#�C�!q�_�FUN�� mo�ZIPu��HR��$L���XZ/MPCF"��`bƀp�rX�ف��LNK���
Ł�0#��� $ !��ބCM+CMk�C8�C"�����P{q $	J8�2�D6!>�O�H� p@T�p@2�����M���sUX�1݅UXE1� ���1C���Y�������8��˗7�FTFG>������_�Z���s �k�� �Ā꜀YD'@ �� 8n�R� Uӱ?$HEIGH��:h#?(! 'v��@�>��� � Gd��qp$B% � E��SgHIF��hRVn�!F�`�HpC� 3� (�8H`O�ѡ�C���+%D	�"�CE�pV��1�SPHER>s� � ,! M��c�u��$POWERFL  �p�|����|�p�RG��`  �������AЋ  ��?�p���pdv��NSb ����?� � Bz|� l�  �<@�|�Z�|�%� ��˃����ŵ��� 2ӷ�� 	UH��l&��౿>���A |�ɻt$��*��/�� **:���p��ȥ��͘���������ɘ��|����� 5�������%ߟ�I� [߉�ߑ������� ����w�!�3�a�W�i� ����������O��� �9�/�A���e�w��� ����'���� �=O}s��� ����k'U K]������ C/��-/#/5/�/Y/ k/�/�/�/?�/�/? �/?�?1?C?q?g?y? �?�?�?�?�?�?_O	O�OIO?OQO�� 	 �O�O�O_�E��3_����O`_�O�_�_÷P?REF Ӻ�p��p
��IORI�TY q|����p����pSPL`z����W�UT�VqÈ�ODU,~�����_?�OG��Gx��R��,f�HIBqOy�|kTOENT 1��~yP(!AF_b��`�o�g!tc�p�o}!ud��o)~!icmX�0bXY̳�kw �|�)� �����p����u ������N�5� r�Y�������̏�����*/c̳ӹ���8E�W�|�>�wx��D���/��4���|���,�7�A��,  ��P����%�|�'���Z��h�z�茯��|��ENHANCE 	#��7�A9�d����� ' �,f�T
�_�Sz����PORTe��rb�@�U��_CARTREP�P|r|brSKSTAgޛkSLGS�`�k����@Un?othing�� ����Ϳ>�P�b�To���TEMP �?isϨE/�_a_?seibanm_�� i_�����0��T�?� x�cߜ߇ߙ��߽��� ����>�)�N�t�_� ������������ �:�%�^�I���m��� �������� ��$ H3lWi��� ����D/ hS�w���u�>��VERSI�P=g�  dis�able��SA�VE ?j	�2670H705��k/!�m//*�/ 	�(%b�O�+	�/�Se?6?H?Z?l?z:%<�/�?4�*']_j` 1�kX �0ubuE�?OqG�P/URGE��Bp`�ncqWF<@�a�TӒ*f�W�`]Daa�WRU�P_DELAY �z�f�B_HOT %?e'b��O�nER_NORMA�L�HGb�O%_�GSE�MI_*_i_�QQS�KIP�3.��3x ��_��_�_�_�]?e o+goKo]ooo5o�o �o�o�o�o�o�o�o 5GYi�}� ������1�C� U��y�g����������я����-�?�7%��$RACFG ��[ќ�3�]�__PARAM�Q3y��S @И@`\�G�42C۠��2M��CbFB�B]��BTIF���J]�C_VTMOU������]�DCR�3��Y ��Q?��9B�2cB��w@�dQ>� �:�lr�]��+�5�Ю�ſ��~�U�_��o ;e��m���KZ;��=g;�4�<�<���f@����� �5�G�Y�k�}� ������ſ׿���xU�RDIO_TYP�E  �V�5��E�DPROT_a��&>��4BHbbCEސSǆQ2c�7 ��B�ꐪ� ����ϐ����&�� ��W�V_~�o����� ����������A�O� m�r���9����� ���������=�_�d� �������������� ��'I�Nm�� ������� #EJi+k� �����//4/ F//g//�/y/�/�/ �/�/�/	?+/0?O/? c?Q?�?u?�?�?�?�?��??;?,O��S�INOT 2�I���l�G;� jO|K���<�O�f�0 �O�K �?�O�?___N_<_ r_X_�_�_�_�_�_�_ �_�_&ooJo8ono�o fo�o�o�o�o�o�o�o "F4j|b� ���������B�O�EFPOS1� 1"�  xO��o×O���� ݏ鈃���Ϗ0��T� �x����7���ҟm� �������>�P���� 7�������W��{�� ���:�կ^������ ����S�e��� ��$� ��H��l��iϢ�=� ��a��υ�� ߻��� �h�Sߌ�'߰�K��� o���
��.���R��� v��#�5�o������ �����<���9�r�� ��1���U��������� ��8#\���� ?��u��"� FX�?��� _��/�	/B/� f//�/%/�/�/[/m/ �/?�/,?�/P?�/t? ?q?�?E?�?i?�?�? O(O�?�?OpO[O�O /O�OSO�OwO�O_�O 6_�OZ_�O~_�_+_=_ w_�_�_�_�_ o�_Do��_Aozocf�2 1r�o.oho�o�o
 o.�oR�oO�# �G�k���� �N�9�r����1��� U����������8�ӏ \���	��U�����ڟ u�����"����X�� |����;�į_�q��� ���	�B�ݯf���� %�����[���ϣ� ,�ǿٿ�%φ�qϪ� E���i��ύ���(��� L���p�ߔ�/�A�S� ��������6���Z� ��W��+��O���s� �������V�A�z� ���9���]������� ��@��d��# ]���}�* �'`���C �gy��&//J/ �n/	/�/-/�/�/c/ �/�/?�/4?�/�/�/ -?�?y?�?M?�?q?�? �?�?0O�?TO�?xOOx�O�o�d3 1�o IO[O�O_�O7_=O[_ �O__|_�_P_�_t_ �_�_!o�_�_�_o{o fo�o:o�o^o�o�o�o �oA�oe �$ 6H�����+� �O��L��� ���D� ͏h�񏌏�����K� 6�o�
���.���R��� ퟈����5�ПY��� ��R�����ׯr��� ������U��y�� ��8���\�n������ �?�ڿc�����"τ� ��X���|�ߠ�)��� ����"߃�nߧ�B��� f��ߊ���%���I��� m���,�>�P���� �����3���W���T� ��(���L���p����� ������S>w� 6�Z���� =�a� Z� ��z/�'/�$/ ]/��//�/@/�/�O�D4 1�Ov/�/ �/@?+?d?j/�?#?�? G?�?�?}?O�?*O�? NO�?�?OGO�O�O�O gO�O�O_�O_J_�O n_	_�_-_�_Q_c_u_ �_o�_4o�_Xo�_|o oyo�oMo�oqo�o�o �o�o�oxc� 7�[���� >��b����!�3�E� ���ˏ���(�ÏL� �I������A�ʟe� ������H�3�l� ���+���O���ꯅ� ���2�ͯV���� O�����Կo������ ���R��v�Ϛ�5� ��Y�k�}Ϸ���<� ��`��τ�߁ߺ�U� ��y���&������� ��k��?���c��� ����"���F���j�� ��)�;�M������� ��0��T��Q�%��I�m��/�$5 1�/���m X���P�t� /�3/�W/�{// (/:/t/�/�/�/�/? �/A?�/>?w??�?6? �?Z?�?~?�?�?�?=O (OaO�?�O O�ODO�O �OzO_�O'_�OK_�O �O
_D_�_�_�_d_�_ �_o�_oGo�_koo �o*o�oNo`oro�o �o1�oU�oyv �J�n���� ���u�`���4��� X��|�ޏ���;�֏ _������0�B�|�ݟ ȟ���%���I��F� ����>�ǯb�믆� �����E�0�i���� (���L���翂�Ϧ� /�ʿS�� ��Lϭ� ����l��ϐ�ߴ�� O���s�ߗ�2߻�V� h�zߴ�� �9���]� �߁��~��R���v�����#�	6 1&����������� ����}���<�� `����CUg ��&�J�n 	k�?�c�� /���	/j/U/�/ )/�/M/�/q/�/?�/ 0?�/T?�/x??%?7? q?�?�?�?�?O�?>O �?;OtOO�O3O�OWO �O{O�O�O�O:_%_^_ �O�__�_A_�_�_w_  o�_$o�_Ho�_�_o Ao�o�o�oao�o�o �oD�oh�' �K]o�
��.� �R��v��s���G� Џk�􏏏���ŏ׏ �r�]���1���U�ޟ y�۟���8�ӟ\��� ���-�?�y�گů�� ��"���F��C�|�� ��;�Ŀ_�迃����� �B�-�f�ϊ�%Ϯ� Iϫ����ߣ�,���xP�6�H�7 1S� ���I��߲������ ��3���0�i���(� ��L���p�����/� �S���w����6��� ��l�������=�� ����6���V� z� 9�]� ��@Rd�� �#/�G/�k//h/ �/</�/`/�/�/?�/ �/�/?g?R?�?&?�? J?�?n?�?	O�?-O�? QO�?uOO"O4OnO�O �O�O�O_�O;_�O8_ q__�_0_�_T_�_x_ �_�_�_7o"o[o�_o o�o>o�o�oto�o�o !�oE�o�o>� ��^����� A��e� ���$���H� Z�l�����+�ƏO� �s��p���D�͟h� 񟌟���ԟ�o� Z���.���R�ۯv�د ���5�ЯY���}�c�u�8 1��*�<� v���߿��<�׿`� ��]ϖ�1Ϻ�U���y� ߝϯ�����\�G߀� ߤ�?���c����ߙ� "��F���j���)� c����������0� ��-�f����%���I� ��m������,P ��t�3��i ���:��� 3��S�w / ��6/�Z/�~// �/=/O/a/�/�/�/ ? �/D?�/h??e?�?9? �?]?�?�?
O�?�?�? OdOOO�O#O�OGO�O kO�O_�O*_�ON_�O r___1_k_�_�_�_ �_o�_8o�_5ono	o �o-o�oQo�ouo�o�o �o4X�o|� ;��q���� B����;������� [�������>�ُ�b�����!�������M�ASK 1 ��⤒���ΗXNO�  ݟ���MO�TE  ���S�_?CFG !Z����N�����PL_RGANGV�N������OWER "���Ϡ��SM_DRYPRG %����%W��եTAR�T #Ǯ�UME_PRO���q����_EXEC_E�NB  ����G�SPDJ�����Ρ�TDB����RM�п��IA_OPTgION��������NGVERS���`�řI_AIRPUR��� R�+���ÛMTE_֐T X���ΐ�OBOT_ISO�LC��������^��NAME8��H��ĚOB_CATEG�ϣ,��S�[��.�ORD_NUM� ?Ǩ���H705  �N��ߨߺ�ΐPC_TIMEOUT��{ xΐS232s��1$��� L�TEACH PENDAN��o����)��V�T��Maintena�nce Cons�N�&�M�"B�P�?No Use6�r� 8��������̒��GNPO$��Ҏ�"Ž��CH_LM��Q���	a�,�!OUD1:��.�RՐ�VAILw���|��*�SR  t�� ���5�R_I�NTVAL��� ���V_DA�TA_GRP 2�'���� D��P�������	� �����B 0RTf���� ��/�/>/,/b/ P/�/t/�/�/�/�/�/ ?�/(??L?:?p?^? �?�?�?�?�?�?�?O  O"O$O6OlOZO�O~O �O�O�O�O�O_�O2_  _V_D_z_h_�_�_�_ �_�_�_�_o
o@o.o�Povodo�o��$S�AF_DO_PU�LSW�[�S���i�S'CAN��������SCà(A��B���+S�S�
����P��q�q�qN� � L^p���5���� ��$���+��r2M�qqd�Y�P�`�J�	t/� @��������ʋ|�� r ք��_ @N�T ��'��9�K�X�T D��X���������ɟ۟ ����#�5�G�Y�k��}�������䅎������Ǧ  ="�;�oR� ����p"�
�u��Di���q$q�?  � ���u q%�\�������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$�6�H�Z����珈�� �����������g� ;�D�V�h�z�������@��������(�Ӣ0� r�i�y���$�7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/?r�+? =?O?a?s?�?�?�?�? �?8��?OO'O9OKO ]OoO�O��$�r�O �O�O�O	__-_?_Q_ c_u_�_�Y�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|�c�路g����� ��0�B�T�f�x����������ҏ����p��:�Ҧ��y��3�	�	123�45678��h�!B!�� +\��p0�� ��Ο�����(�:� @��c�u��������� ϯ����)�;�M� _�q�����R���ɿۿ ����#�5�G�Y�k� }Ϗϡϳ����ϖ��� ��1�C�U�g�yߋ� �߯���������	�� -���Q�c�u���� ����������)�;� M�_�q���B������ ����%7I[ m������� �!3EWi{ �������/ ///�S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?D/�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O*����O	_�E�?5_�G_Y_�yCz  �A��z   ���x2�r }��)�
�W_�  	�*�2�O �_�_ oo"l�#\��_hozo�o�o�o�o �o�o�o
.@R dv����Mo� ���*�<�N�`�r� ��������̏ޏ��� �&�8�J��X #P$Pt�Q�R<u� k�~�Q  �������S�P���Q�Qt�  �PÙ۟�P(� `,b����]��PFl�$SCR_�GRP 1*B�+B4� �� �,a ��U	 v��~������ d���%���ɯ���h]���P�D1� D7n��3��Fl�
CRX-10�iA/L 234�567890�P�d� r��Pd�L ��,a
1o�����Z���[ ¶~� +fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@��R�d�t���H�~�Ă�m��ϴ�@�����ϼ��,a�Ϡ1���U�[�G�imXh�uP,[~����B�  BƠߞҷ�r��A�P��  @1`��՚�@����� ?	���H����ښ�F@ F�`A� I�@�m�X��|���� ��������������`:�%�7�I�[�B�i� ��������������� -Q<u`��@En�ٯ���W�P�"+f@_�5��1`4b���x����ͣ�O�,dA����$���Fa�,a �#!"/4/E-!�Z(f/x/G/ (�P�!(� �/�/�/��/�/?#9b�����S7س�M�ECLV�L  ,a���ݲ�Q@f1L_D?EFAULTn4b1_�1`�3?HOTSTR�=���2MIPOWER�Fm0pU�5�4W7FDO�6 �5L��ERVENT 1�+u1u1�3 L!�DUM_EIP�#?5H�j!AF�_INE�0SO,d!'FT)O�NIO�O9!���O ��O�O�!RPC_MAIN�O�H��O>_S'VIS_�I�-_�_?!OPCUf�_�Wy_�_!TMP�PPU�_<Id�_�"o!
PMON_�PROXY#o?Fe ono�R<o8Mf]o�o�!RDM_SR�V�o<Ig�o!�R��"=Hh�oR!%
PM�o9LiA��!RLSYNC̟�y8��!gROS(O��4��6�!
CE�PMT'COM7�?Fk%���{!	K�CONS���>Glq�Ώ!K�WOASRC�o?Fm��v�!K�USB��=Hn	�f�!STM�0��;JoU����O�֟�c����CICE�_KL ?%K� (%SVCPGRG1��G�1�2G�DL�6�3o�t�6�4��D��6�5��į6�6��6�7��6���W�R�9_�d�3��� 6�9���6�a�ܿ6��� �6���,�6�ٯT�6� �|�6�)���6�Q��� 6�y���^����^�ʿ D�^��l�^�ϔ�^� Bϼ�^�j���^���� ^���4�^���\�^�
� �2���6��/� ���V��<�'�`�K� ��o����������� ��&J5nY� ������� 4F1jU�y� ����/�0// T/?/x/c/�/�/�/�/ �/�/�/??>?)?P?�t?_?�?
�_DEV� I�M{C:�84���4?GRP 2/E�0�+�bx 	�� 
 ,@�0 �?OD8OJO1OnOUO �O�O�O�O�O�O�O�O "_	_F_-_j_|_c_�_�[E�1�_�_�_o �_'ooKo]oDo�oho �o�o�o�o�o�o�o�o 5Y�_D�u�C �����
��� @�'�d�K�]������������ۏ�o	A %�S�:�w���_���� Ο����(��L� 3�E���i�����ʯܯ �_ ����6���Z�A� ~���w�����ؿ�ѿ ���2�D�+�h�Oό�s�E����f���� ��τ��'߅�v�]� �߁߾��߷������ *�5�N��r���� �����������&�8� �\�C���g�y����� ������g�4- jQ�u���� �B)fx _����)�� /,//P/7/t/[/m/ �/�/�/�/�/?�/(?�?L?^?E?�?�7d ��[~
�6 �s 	 A;�*=� 6?�=����D�>ޟ���g�:�0���ī��|@��-�@�5_�eA5�-�=�BG+h�&����6)AB�m�����`x���=�?7O%TEL�EOP8OcN[~�y��5�o�ʾ�TF�����������|��ҝ����E��1�E@�*��A`�~�n��!��$�A����M�Y<T�������C=��J����Gc��McO��IJO/_��[~��6r� _�1<�׻���y;��	A�`�ʛ1bP��N	�V�A�&@���@���@)�E�]�1������0ד� x����Q��U?�Q��O�__ _�oDU�NU9���6>���E��bQ�2]�j_ ���rAS��AT�@���@G$�_ ���yC� �Pr�}��Q� 2i?�R�_�o�_�_�o�DU�K�5��l�������S����`
�� 3�>v�ĚM@��@�V�@��%@��Ŀ�qߝ��]V�N���N�!C(u�µ�� �®�ɒow�o��o�DU�b�5?������T�@O��P�%�*�?-��Ƒ�N�P�A����
Q�@���q��A��M�{��B&�br�'C9rt�1��^ѺfK��������pm�5>����@«���͙~�E�A�����c�N�'pA(�AC�8AD����ߧA�y�Nd��A��R����������s��`_�^��\�n��S�BW�c�v"���?/���H�?��4@� ��+79��$Ώ�A8	AAl���c`�f�@��c+�Ne?6A��z2��LQ� �f��t���`�D��2�D�)�DS �I�IV�D�z�h�������ԯ%�/���ho֯ 0��T�B�x�f���ޯ ÿ��������,�� P�>�t϶���ڿd��� �������(��Lߎ� s߲�<ߦߔ��߸��� ����$�f�K���~� l��������,�� #�������D�z�h��� �������(���
 ,.@vd����  ���(* <r���b�� ��//$/z�q/ �J/�/�/�/�/�/�/ ?R/7?v/ ?j?�/z? �?�?�?�?�?*?ON? �?BO0OfOTOvO�O�O �OO�O&O�O__>_ ,_b_P_r_�_�O�_�O �_�_�_oo:o(o^o �_�o�oNopoJo�o�o �o 6xo]�o& �~������ P5�t�h�V���z� �������(��L�֏ @�.�d�R���v���� ��$�����<�*� `�N���Ɵ���t�ޯ p����8�&�\��� ��¯L�����ڿȿ� ���4�v�[Ϛ�$ώ� |ϲϠ��������N� 3�r���f�Tߊ�x߮� �����������߾� ,�b�P��t������ �������(�^� L��������r�����  ��$Z��� ��J������ b�Y�2�z �����:/^ �R/�b/�/v/�/�/ �//�/6/�/*??N? <?^?�?r?�?�/�?? �?O�?&OOJO8OZO �O�?�O�?pO�O�O�O �O"__F_�Om__6_ X_2_�_�_�_�_�_o `_Eo�_oxofo�o�o �o�o�o�o8o\o�o P>tb���� �4�(��L�:� p�^�����͏���  ��$��H�6�l��� ��ҏ\�ƟX�֟���  ��D���k���4��� ��¯��ү����^� C����v�d������� ��ο��6��Z��N� <�r�`ϖτϺ����� �Ϫ��Ϧ��J�8�n� \ߒ��Ϲ��ς����� �����F�4�j�ߑ� ��Z������������ �B���i���2����� ����������J�p�A ��tb���� �"F�:�J p^����� �/ /6/$/F/l/Z/ �/��/��/�/�/? �/2? ?B?h?�/�?�/ X?�?�?�?�?
O�?.O p?UOgOO@OO�O�O �O�O�O_HO-_lO�O `_N_p_r_�_�_�_�_  _oD_�_8o&o\oJo lono�o�o�_�oo�o �o4"XFh�o �o��o����� 0��T��{��D��� @����ҏ���,�n� S������t������� ��Ο�F�+�j���^� L���p�������ܯ� �B�̯6�$�Z�H�~� l����ɿۿ������ ��2� �V�D�zϼ��� �j�����������.� �Rߔ�y߸�B߬ߚ� �߾�������*�l�Q� ����r������ ��2�X�)�h��\�J� ��n�������
���.� ��"��2XF|j ������� .TBx��� h����//*/ P/�w/�@/�/�/�/ �/�/�/?X/=?O?? (??p?�?�?�?�?�? 0?OT?�?HO6OXOZO lO�O�O�OO�O,O�O  __D_2_T_V_h_�_ �O�__�_�_�_o
o @o.oPo�_�_�o�_vo �o�o�o�o<~o c�o,�(��� ���V;�z�n� \�������ȏ���.� �R�܏F�4�j�X��� |���ğ��*���� �B�0�f�T���̟�� ïz���v����>� ,�b�����ȯR����� ̿ο���:�|�a� ��*ϔςϸϦ����� ���T�9�x��l�Z� ��~ߴߢ����@�� P���D�2�h�V��z� ��������
���� @�.�d�R�������� x�������<* `�����P��� ��8z_� (������� @%/7/�/�X/�/ |/�/�/�//�/</�/ 0??@?B?T?�?x?�? �/�??�?O�?,OO <O>OPO�O�?�O�?vO �O�O_�O(__8_�O �O�_�O^_�_�_�_�_� o�_$of_Ko�_` � �$SERV�_MAIL  ʖU�`��QvdOU�TPUT�h��P@vdRV �20f  �` �(a\o�ovdSAV�E�l�iTOP10� 21�i d �6 s�P6r _�P2oXj |������� ��0�B�T�f�x��� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�:��guYP�cFZ�N_CFG 2e�c�T�a�e~|�GRP 23���q ,B   �AƠ�QD;� B}Ǡ�  B4�S�RB21�fH7ELL�4ev��`�o��/�>�%RSR>�?�Q���u� ����ҿ������,π�P�;�t�_Ϙϩ�~���  � �����Ϸͻ��P��&�'�ސW��2Pd��g��HKw 15�� ,� �߫ߥ��������� @�;�M�_���������������OMM� 6��?��FT?OV_ENB�d�a�u�OW_REG�_UI_��bIMI_OFWDL*�7.��ɥ��WAIT\� `ٞ����`���d��wTIM�������VA�`����_UNcIT[�*yLCy�WTRY��uv`ME�8���aw֑dt ��9� ������<���X�Pڠ6p`?�  ��o+=Ip�VL�l�fMO�N_ALIAS k?e.��`heGo ������/)/ ;/M/�q/�/�/�/�/ d/�/�/??%?�/I? [?m??�?<?�?�?�? �?�?�?!O3OEOWOO {O�O�O�O�OnO�O�O __/_�OS_e_w_�_ �_F_�_�_�_�_�_o +o=oOoaoo�o�o�o �o�oxo�o'9 �o]o��>�� ����#�5�G�Y� k��������ŏ׏�� ����1�C��g�y� ����H���ӟ���	� ��-�?�Q�c�u� ��� ����ϯᯌ���)� ;��L�q�������R� ˿ݿ��Ͼ�7�I� [�m��*ϣϵ����� �ϖ��!�3�E���i� {ߍߟ߱�\������� ����A�S�e�w�� 4����������� +�=�O���s������� ��f�����'�� K]o��>�� ���#5GY�}����l��$SMON_DE�FPROG &������ &*SYS�TEM*���R�ECALL ?}�� ( �}7�copy frs�:orderfi�l.dat vi�rt:\tmpb�ack\=>19�2.168.56.1:2796/ؓ/�/�.}.K"mdb:*.*`/r.z/�??/?�%2xK$:1\�/U0�/6 �/�?(�?�?�!3K5aS?e? �$?O"O4O� J/\/ �/ O�O�O�O�/cO�/ ~O_!_3_F?�?�O|? �_�_�_�?U_g_�?o o/oBOTO�OxO�o�o �o�O�Omo�O+ >_P_�_t_����_��__�_��'��m
�xyzrate 11 �������䯏�eK�k�18540 j�|���1���ctpdisc 0Տ������������etpconn 0 T�f�x�	��-��g8Ko]oS���������m/�of�މ {���0��}�f�� ���������`4�\� َ���#�5�H�Z�� ���ϡϳ�Ưa��|� ��1�D�׿�z��� �߯�¿S�e���	�� -�@�R�����ߌ�� ��C�͒ԏd�v��� +�>�P���tυ����� ����i���':� L���p���8�� [m�#5H�Z� ���������a�� |//1/D��z �/�/�/�S/e/�	? ?-?@R�v�?�? �?��k?�OO)O </N/�/r/�O�O�O�/ �/]O�/�O_%_�OJ? \?�? _�_�_�_�?c_��?~_o!o3oDP�$�SNPX_ASG 2:���Va� ��DP%�7o~o  ?��GfPARAM �;Ve`a ��	lkP>TDP�>X�d� ���I`OFT_KB_?CFG  CS\e�FcOPIN_SI�M  Vk�b�+=OYsI`RVN�ORDY_DO � �eukrQS�TP_DSB~��b�>kSR <�Vi � & TELEO�e�{v�>TW`I`TOP_ON_ERRxGb��PTN Ve�P��D:�RI?NG_PRM'��r�VCNT_GP �2=Ve�ac`x 	���DP��я�����BgVD�RP 1	>�i�`�Vq؏0� B�T�f�x��������� ҟ�����,�>�e� b�t���������ί� ��+�(�:�L�^�p� ��������ʿ�� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�}�zߌߞ߰� ��������
��C�@� R�d�v������� ��	���*�<�N�`� r��������������� &8J\n� ������� "4[Xj|�� �����!//0/ B/T/f/x/�/�/�/�/ �/�/�/??,?>?P? b?t?�?�?�?�?�?�?��?O�PRG_CoOUNT�f�P�N)IENBe�+EMUC��dbO_UPD 1}?�{T  
O DR�O�O�O�O�O__ A_<_N_`_�_�_�_�_ �_�_�_�_oo&o8o ao\ono�o�o�o�o�o �o�o�o94FX �|������ ���0�Y�T�f�x� ������������� 1�,�>�P�y�t����� ����Ο��	���(� Q�L�^�p��������� �ܯ� �)�$�6�H� q�l�~�������ƿؿ ���� �I�D�V�"L�_INFO 1@��E�@��	� yϽϨ�����?���?����P`�3����� ���EA��mm�2&�����K�wC�����  @`�� ?�`i�=����� D/  �� Ce��?�3��´j�|��-@YSDEBUG�:@�@�o�d�I��S�P_PASS:E�B?��LOG uA���A  o�9i�v�  �Ao�UD1:\��<}���_MPC�ݚEHk�}�A&�� �A~K�SAV B��`IA���*�i�1��SVB�TEM_T�IME 1C����@ 0  �6n�.i�"��*����MEMBK  	�EA�����ޡ�X|�@� 	@��$����������dh�9
�� ��@�`r��������� � @Rdv�����
Le�//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H?Z?��SKV�[�EAj�К?�?�?��
7�B�]2���?i�  0H]
:O.@R��O�O�O}N�o�c ��OBD��O�_'_9_-L2��Y_�_�_�_�_�_o�U �_�_�o'o9oKo]o oo�o�o�o�o�o�o�o �o#5GYk_?�T1SVGUNS�PD�� '�����p2MODE_LIM D��Ҋt�2�p�qE�݉uA�BUI_DCS H}5���0�G� 0��D��|-�X�>���o*���� 
���e��i���r�i������uEDIT� I��xSCR/N J���rS�G K�.�(�0�߅SK_OPTI�ON��^����_D�I��ENB  �/����BC2_G_RP 2L��󘵟L�MPC�ʓ�|B�CCF/�N���� ����FV�<��� `�K���o�����̯ޯ ɯ��&��J�5�n� Y�k�����ȿ���׿ ���4�F�1�j�Uώ� ��̀�϶�������v� �
�/�U�@�yߧ�� `�iМ��߰�����
� ��.��>�@�R��v� �����������*� �N�<�r�`������� ��������̀4 FX��|j��� ����B0 fTvx���� �/�,//</b/P/ �/t/�/�/�/�/�/�/ �/(??L?d?v?�? �?�?6?�?�?�?O O 6OHOZO(O~OlO�O�O �O�O�O�O�O __D_ 2_h_V_�_z_�_�_�_ �_�_
o�_.oo>o@o Ro�ovo�ob?�o�o�o �o<*Lr` �������� &��6�8�J���n��� ��ȏ���ڏ��"�� F�4�j�X���|����� ���֟��o$�6�T� f�x���������ү�� �����>�,�b�P� ��t��������ο� �(��L�:�\ς�p� �ϔ��ϸ������� � �H�6�l�"��ߖߴ� ����V������2� � V�h�z�H������ ��������
�@�.�d� R���v����������� ��*N<^` r������� &8�\Jl�� ������"// F/4/V/X/j/�/�/�/ �/�/�/?�/?B?0? f?T?�?x?�?�?�?�? �?O�?,O�DOVOtO �O�OO�O�O�O�O�O�_ V4P�$TBC�SG_GRP 2�O U� � �4Q 
 ?�  __q_[_�_ _�_�_�_�_�_o%k�8R?SQF\d��HTa?4Q	 H�A���#e>����>$a�\#eAT��A WR�o�h|djma�G�?Lfgr�bp�o�n�ffhfG��ͼb4P|j��o�*}@��Rhf�ff>�33pa#e<q!B�o+=xrRp�qrUy�rt~��H�y0 rIpTv�pBȺt~ 	xf	x(�;���f����N�`���ˏڋ�����	V3.00~WR	crxlڃ	*��3R~t2��HH��� \�.�n]�  cC.�X����8QJ2?SRF]�����CFG -T UPQ SPܚ+��r�ܟ1��1�W�e�	Pe� ��v�����ӯ����� ���Q�<�u�`��� ������Ϳ�޿�� ;�&�_�Jσ�nπϹ� ��������WRq@� 0�B���u�`߅߫ߖ� �ߺ������)�;�M� �q�\������4Q  _���O ���J�8� n�\������������� ����4"XFh j|������ .TBxf� �nO����// >/,/b/P/�/t/�/�/ �/�/�/�/�/?:?(? ^?p?�?�?N?�?�?�? �?�?�? O6O$OZOHO ~OlO�O�O�O�O�O�O �O __D_2_T_V_h_ �_�_�_�_�_�_
o�_ o@o�Xojo|o&o�o �o�o�o�o�o* N`r�B��� ����&��6�\� J���n�����ȏ��؏ ڏ�"��F�4�j�X� ��|���ğ���֟� ��0��@�B�T���x� ����ү䯎o���̯ ʯP�>�t�b������� �������Կ&�L� :�p�^ϔϦϸ��τ� ����� �"�H�6�l� Zߐ�~ߴߢ������� ���2� �V�D�z�h� ������������� 
�,�.�@�v����� ��\�������< *`N����x ���8J\ (������ ��/4/"/X/F/|/ j/�/�/�/�/�/�/�/ ??B?0?f?T?v?�? �?�?�?�?�?OO�� 2ODO�� O�OtO�O�O �O�O�O_�O(_:_L_ 
__�_p_�_�_�_�_ �_ o�_$oo4o6oHo ~olo�o�o�o�o�o�o �o D2hV� z�����
�� .��R�@�b���v��� &OXO֏菒����� N�<�r�`�������̟ ޟ🮟��$�&�8� n�������^�ȯ��� گ��� �"�4�j�X� ��|�����ֿĿ�� ��0��T�B�x�fψ� �Ϝ����������� >�P���h�zߌ�6߼� �����������:�(� ^�p���R�����8�� ���  &�*�� *�>�*��$�TBJOP_GR�P 2U����  ?�/��C*�	V�]��Wd������X  �*��� �,� � ���*�� @&�?��	 ߐA�����C��  DD�����>~v�>\? ���aG�:�o���;ߴAT������A�<��M�X����>��\)�?���8Q�|����L��>�0 ^&�;iG.���Ap< � F�A�ff�v��� ^):VM�.�� �S>o*�@��R�Cр	���������ff�:��6/�?�33�B   ��/�������>):�S���� �/�/@��H�%&/��/��=� <#��
*��v�;/��f�!?���4B�3 ?'?2	��2?hZ?D? R?�?�?�?F?�?�?�? �?OAOO�?`OzOdO�rO�O�O*�C�*����A��	V3.0}0{�crxl��*P��%�%c5Z F� JZ�H F6� F�^ F�� F��f F� G�� G5 G�<
 G^] G�� G���G��*�G�S G��; G��ERD�u�\E[� E�� F( F�-� FU` F�}  F�N F�� F�� F�ͺ F� F��V G� G�z Ga 9'ѷ�Q�LHefJQ4�o,b*�0c�1���OH�ED_TCH Xd�+X2S��&�&�d$�'X�o�o*�1F�T�ESTPARS c ��cV�HRpABLE 1Yd� N`*�����g)$j�g�h�h)�T1��g	�h
�h�hTHu*��h�h�h�%vRDI0n��GYk}��u	�O �#�-�?�Q�c�u�)r	S�l� �z6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ��I���m�Fwͩ�� ȏڏ쏘������x)r��NUM  ���n����2� Ep�)r_CF�G Z��I���@�V�IMEBF_T�TqD��e޶VE�R�����޳R {1[8{ 8�o�*�%�Q� ��د  9�K�]�oρϓϥ� �����������#�5� G�Y�k�}��ߡ߳��� ��������1���E� W�i�{�������� ������/�A�S�e� w���������������@+=O�_����@��`LIF7 \��D`�����DR�(FP
��!p�!p� d�� ��MI_CHA�N� � DB/GLVL��f�ETHERAD S?u��0`1��_}�ROUT6�!�j!��~SNMASKY|�j255.%�S///A/S�`OOLOFS_DIp��CORQCTRL ]8{��1o�-T�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OL�/6O%O�ZOcPE_DET�AI7�*PGL_�CONFIG �c������/c�ell/$CID?$/grp1^O�O �O�O
__|���G_ Y_k_}_�_�_0_�_�_ �_�_oo�_CoUogo yo�o�o,o>o�o�o�o 	-�oQcu� ��:����� )���_�q���������׮}N����%�@7�I�a�KOq�P��M� ����ʟܟ� �G�$� 6�H�Z�l�~������ Ưد������2�D� V�h�z������¿Կ ���
ϙ�.�@�R�d� vψϚ�)Ͼ������� �ߧ�<�N�`�r߄� ��%ߺ��������� &��J�\�n���� 3����������"��� F�X�j�|��������@��User �View �I}}�1234567890����+=�Ex �e����2 ��B������`r��3�Oas@����x4> //'/9/K/]/�~/x5��/�/�/�/�/?p/2?x6�/k?}?��?�?�?�?$?�?x7 Z?O1OCOUOgOyO�?�Ox8O�O�O�O	_�_-_�ON_TR �lCamera���O�_�_�_�_�_�_˂E�_o)o;n���Uogoyo�o�o�o�)  mV�	�_�o#5 GY o}���o�@�����F_�mV =�k�}�������ŏ l����X�1�C�U� g�y���2�D��"�ן �����1�؏U�g� y�ğ������ӯ��� ��D��k��E�W�i�{� ����F�ÿտ�2�� �/�A�S�e��nUY9 ������������	߰� -�?�Qߜ�u߇ߙ߫� ����v�D�If��-� ?�Q�c�u�ߙ��� �������)�;��� D��I����������� ����)t�M_@q���N�`�93 ��0B��S x�1�����(//�J	oU0�U/ g/y/�/�/�/V�/�/ �/�?-???Q?c?u? /./tPv[?�?�?�? OO(O�/LO^OpO�? �O�O�O�O�O�O�?oU �k�O:_L_^_p_�_�_ ;O�_�_�_'_ oo$o 6oHoZo_;%N��_�o �o�o�o�o �_$6 H�ol~���� moe��]�$�6�H� Z�l��������؏ ���� �2��e&� ɏ~�������Ɵ؟� ��� �k�D�V�h�z� ����E�e��5���� � �2�D��h�z��� ׯ��¿Կ���
ϱ�  ��9�K�]� oρϓϥϷ���������   ��5� G�Y�k�}ߏߡ߳��� ��������1�C�U� g�y���������� ��	��-�?�Q�c�u� ���������������);M_q� � 
��(  �>-�( 	 �� �����#3 5G}k����
� �Y�
// ./��R/d/v/�/�/�/ ����/�/�/A/?0? B?T?f?x?�/�?�?�? ?�?�?OO,O>O�? bOtO�O�?�O�O�O�O �O_KO]O:_L_^_�O �_�_�_�_�_�_#_ o o$ok_HoZolo~o�o �o�_�o�o�o1o  2DVh�o�o�� �	��
��.�@� �d�v��������Џ ���M�*�<�N��� r���������̟�%� ��&�m�J�\�n��� �����ȯگ�3�� "�4�F�X�j������� ����ֿ�����0� w���f�xϊ�ѿ���� �������O�,�>�P� ��t߆ߘߪ߼���� ����]�:�L�^�p�p����߻@ ����������� ���"frh:\t�pgl\robo�ts\crx!�1�0ia_l.xml��D�V�h�z�����`�������������� 0BTfx�� �������, >Pbt���� ����/(/:/L/ ^/p/�/�/�/�/�/�/ ��/?$?6?H?Z?l? ~?�?�?�?�?�?�/�? O O2ODOVOhOzO�O �O�O�O�O�?�O
__ ._@_R_d_v_�_�_�_ �_�_�O�_oo*o<o No`oro�o�o�o�o�ot�n �6� ���<< 	� ?��k!�o;i Oq������ ���%�S�9�k����o�����я����(��$TPGL_O�UTPUT f������� �&�8�J�\�n��� ������ȟڟ���� "�4�F�X�j�|�����в�į�p�ր23�45678901 �����1�C�K��� �r���������̿d��п��&�8�J��} T�|ώϠϲ���\�n� ����0�B�T���b� �ߜ߮�����j���� �,�>�P����߆�� �������x����(� :�L�^���l������� ����t���$6H Zlz���� ��� 2DVh  ������ �/./@/R/d/v// �/�/�/�/�/�/�/ۂ? $$��ί <7*?\?N?�?r?�?�? �?�?�?�?OO4O&O XOJO|OnO�O�O�O�O��O�O_�O0_"_T_} �an_�_�_�_�_�_�]�@�_o	z ( 	 V_Do2oho Vo�ozo�o�o�o�o�o 
�o.R@vd �������� �(�*�<�r�`���ܦ��  << I_ˏݏ������� :�L�֪��}���)��� ş�������k��C� ݟ/�y���e������ �������-�?��c� u�ӯ]�����W��� Ϳ��)χ���_�q�� yϧρϓ�����M�� %߿��[�5�Gߑߣ� ߫���s����!��� E�W��?���9��� ������i���A�S� ��w���c�u����/� ����=)s �����U�� �'9�!o	[ �����K�#/ 5/�Y/k/E/w/�/� /�/�/�/�/?�/? U?g?�/�?�?7?�?�?�?�?	OO��)WGL1.XML�_�PM�$TPOFF_LIM ���P����^FN_�SVf@  �T�xJP_MON Mg��zD�P�P�2ZISTRTCHOK h��xFk_�aBVTCOMPA�T�HQ|FVWVA/R i�M:X�D� �O R_�P��BbA_DEFP�ROG %�I�%TELEOP�i_�O_DISPL�AYm@�N�RINST_MSK  �\� �ZINUSsER_�TLCKl��[QUICKMEyN:o�TSCREY`���Rtpsc�Tat`yixB�`�_�iSTZxIRA�CE_CFG Uj�I:T�@	[T�
?��hHNL C2k�Z���aA[ gR -?Qcu�����z�eITEM 2�l{ �%$1�23456789y0 ��  =<
�x0�B�J�  !P�X�dP���[S��� "���X�
�|���W� ��r�֏����.��0� B�\�f�����6�\�n� ҟ��������>�� �"���.�����ίR� ���Ŀֿ:��^�p� 9ϔ�Tϸ�xϊ�� �d���H��l��>� Pߴ�\�������v� � �����h�(�ߞ߰� 4�L��ߦ�����@� R��v�6���Z�l��� �������*���N���  ������������X ���J
n� ��b���� "4F�/|</N/ �Z/���//�/0/ �/?f/?�/�/e?�/ �?�/�?�?�?,?�?P? b?t?�?�?DOjO|O�? �OOO(O�O�O^O_ 0_�O<_�O�O�_�O�_ _�_�_H_�_l_~_Go��dS�bm�oLj�g  �rLj �a�o�Y
 �o�o�o��o{jUD1:\�|��^aR_GR�P 1n�{� 	 @�PRd{�N�r����~� �p���q+��O�:�?�  j�|�f� ���������ҏ��� �>�,�b�P���t���������	e���~\cSCB 2ohk U�R�d�v����������Я�RlUT�ORIAL p�hk�o-�WgV_CONFIG qhm��a�o�o��<�OUT?PUT rhi}�����ܿ� � �$�6�H�Z�l�~ϐ� �ϴ�z�ɿ���� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r �������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/��/�/??0?B? T?f?x?�?�?�?�?�/ �?�?OO,O>OPObO tO�O�O�O�O�?�O�O __(_:_L_^_p_�_ �_�_�_�_f�x�ǿo o,o>oPoboto�o�o �o�o�o�o�O( :L^p���� ���o ��$�6�H� Z�l�~�������Ə؏ ��� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я���� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t�����������������X���#��N �_r������ �&8J��n �������� /"/4/F/X/i|/�/ �/�/�/�/�/�/?? 0?B?T?e/x?�?�?�? �?�?�?�?OO,O>O POa?tO�O�O�O�O�O �O�O__(_:_L_^_ oO�_�_�_�_�_�_�_  oo$o6oHoZok_~o �o�o�o�o�o�o�o  2DVgoz�� �����
��.� @�R�d�u�������� Џ����*�<�N� `�q���������̟ޟ ���&�8�J�\�k���$TX_SCR�EEN 1s%� �}��k�����ӯ���	� ��Z��I�[�m���� ���,�ٿ����!� 3Ϫ�W�ο{ύϟϱ� ����L���p��/�A� S�e�w��� ߭߿��� �����~�+��O�a� s���� ���D��� ��'�9�K������ ����������R���v� #5GYk}�����$UALRM_�MSG ?����� �n��� 	:-^Qc������� /�SEoV  �2&��ECFG uv����  n��@�  Ab!  w B�n�
 / u����/�/�/�/�/�/�??%?7?I?W7>!G�RP 2vH+ 0n�	 /�?� �I_BBL_NO�TE wH*T?��lu����w�T �2DEFP�RO� %� (�%�Ow�	OBO-B?TELEOPGO#O �O�O�O�O�O�O�O_��O&_�?�0FKEYDATA 1x����0p W'n���?�_�_z_�_�_�Z,�(�_on�(PO?INT ERon  IRECT@o�ko�PNDUo�oOcC?HOICE]�onTOUCHU`O �o�_�o7[m T�x�������!��E��Z���/frh/gui�/whiteho?me.pngQ��������ŏ׏�h�pointz���/��A�S��  i�direc��������şןf�/iny��"��4�F�X��m�choicy�������ͯ߯��h�touchup���/�A�S�e���h�arwrg �����ÿտ�n�� �(�:�L�^�p����� �ϸ�������}��$� 6�H�Z�l��ϐߢߴ� �������ߋ� �2�D� V�h�z�	������� ������.�@�R�d� v���_����������� ���2DVhz ������
 �@Rdv�� )����//� </N/`/r/�/�/%/�/ �/�/�/??&?�/J? \?n?�?�?�?3?�?�? �?�?O"O�?4OXOjO |O�O�O�OAO�O�O�O __0_�OT_f_x_�_ �_�_=_�_�_�_oo ,o>o�_boto�o�o�o��oW��k�b�����o}�o8J$v,6�{.�� �������/� �S�:�w���p����� я�ʏ��+��O� a�H���l�������ߟ ���'�9�Ho]�o� ��������ɯX���� �#�5�G�֯k�}��� ����ſT������ 1�C�U��yϋϝϯ� ����b���	��-�?� Q���u߇ߙ߽߫��� ��p���)�;�M�_� �߃��������l� ��%�7�I�[�m��� ������������z� !3EWi���� �����П/ ASew~��� ���/�+/=/O/ a/s/�//�/�/�/�/ �/?�/'?9?K?]?o? �?�?"?�?�?�?�?�? O�?5OGOYOkO}O�O O�O�O�O�O�O__ �OC_U_g_y_�_�_,_ �_�_�_�_	oo�_?o Qocouo�o�o�o:o�o �o�o)�oM_ q���6������%�7�9�}����b�@t���^�������,�� 돞����3�E�,�i� P�������ß����� ����A�S�:�w�^� ������ѯ����ܯ� +�
O�a�s������� �Ϳ߿���'�9� ȿ]�oρϓϥϷ�F� �������#�5���Y� k�}ߏߡ߳���T��� ����1�C���g�y� ������P�����	� �-�?�Q���u����� ������^���) ;M��q���� ��l%7I [������ h�/!/3/E/W/i/ @��/�/�/�/�/�/� ??/?A?S?e?w?? �?�?�?�?�?�?�?O +O=OOOaOsOO�O�O �O�O�O�O_�O'_9_ K_]_o_�__�_�_�_ �_�_�_�_#o5oGoYo ko}o�oo�o�o�o�o �o�o1CUgy ������	� ��?�Q�c�u����� (���Ϗ������ ;�M�_�q�������~ ����~ ���ҟ���Ο�*��,�[���f��� ����ٯ�������3� �W�i�P���t���ÿ ���ο��/�A�(� e�Lωϛ�z/������ ����(�=�O�a�s� �ߗߩ�8�������� �'��K�]�o��� ��4����������#� 5���Y�k�}������� B�������1�� Ugy����P ��	-?�c u����L�� //)/;/M/�q/�/ �/�/�/�/Z/�/?? %?7?I?�/m??�?�? �?�?�?���?O!O3O EOWO^?{O�O�O�O�O �O�OvO__/_A_S_ e_�O�_�_�_�_�_�_ r_oo+o=oOoaoso o�o�o�o�o�o�o�o '9K]o�o� �������#� 5�G�Y�k�}������ ŏ׏������1�C� U�g�y��������ӟ ���	���-�?�Q�c� u��������ϯ��h���0���0���B�T�f�>�����t�,��˿~� �ֿ�%��I�0�m� �fϣϊ��������� ��!�3��W�>�{�b� �߱ߘ��߼�����? /�A�S�e�w��� ������������=� O�a�s�����&����� ������9K] o���4��� �#�GYk} ��0����/ /1/�U/g/y/�/�/ �/>/�/�/�/	??-? �/Q?c?u?�?�?�?�? L?�?�?OO)O;O�? _OqO�O�O�O�OHO�O �O__%_7_I_ �m_ _�_�_�_�_�O�_�_ o!o3oEoWo�_{o�o �o�o�o�odo�o /AS�ow��� ���r��+�=� O�a����������͏ ߏn���'�9�K�]� o���������ɟ۟� |��#�5�G�Y�k��� ������ůׯ����� �1�C�U�g�y���� ����ӿ������-�@?�Q�c�uχ�^P����^P���������ͮ���
���, ��;���_�F߃ߕ�|� �ߠ����������7� I�0�m�T������ �������!��E�,� i�{�Z_���������� ���/ASew ������ �+=Oas� �����//� 9/K/]/o/�/�/"/�/ �/�/�/�/?�/5?G? Y?k?}?�?�?0?�?�? �?�?OO�?COUOgO yO�O�O,O�O�O�O�O 	__-_�OQ_c_u_�_ �_�_:_�_�_�_oo )o�_Mo_oqo�o�o�o �o���o�o%7 >o[m���� V���!�3�E�� i�{�������ÏR�� ����/�A�S��w� ��������џ`���� �+�=�O�ޟs����� ����ͯ߯n���'� 9�K�]�쯁������� ɿۿj����#�5�G� Y�k����ϡϳ����� ��x���1�C�U�g� �ϋߝ߯�����������`����`���"�4�F��h�z�T�,f���^���� �����)��M�_�F� ��j����������� ��7[B� x�����o! 3EWixߍ�� �����///A/ S/e/w//�/�/�/�/ �/�/�/?+?=?O?a? s?�??�?�?�?�?�? O�?'O9OKO]OoO�O O�O�O�O�O�O�O_ �O5_G_Y_k_}_�__ �_�_�_�_�_o�_1o CoUogoyo�o�o,o�o �o�o�o	�o?Q cu��(��� ���)� M�_�q� �������ˏݏ�� �%�7�Ə[�m���� ����D�ٟ����!� 3�W�i�{������� ïR������/�A� Яe�w���������N� �����+�=�O�޿ sυϗϩϻ���\��� ��'�9�K���o߁� �ߥ߷�����j���� #�5�G�Y���}��� ������f�����1��C�U�g�>�i��>>�������� ����������,� �?&cu\�� �����) M4q�j��� ��/�%//I/[/ :�/�/�/�/�/�/�� �/?!?3?E?W?i?�/ �?�?�?�?�?�?v?O O/OAOSOeO�?�O�O �O�O�O�O�O�O_+_ =_O_a_s__�_�_�_ �_�_�_�_o'o9oKo ]ooo�oo�o�o�o�o �o�o�o#5GYk }������ ��1�C�U�g�y��� �����ӏ���	��� -�?�Q�c�u�����p/ ��ϟ�����;� M�_�q�������6�˯ ݯ���%���I�[� m������2�ǿٿ� ���!�3�¿W�i�{� �ϟϱ�@�������� �/߾�S�e�w߉ߛ� �߿�N�������+� =���a�s����� J�������'�9�K� ��o�����������X� ����#5G��k�}���������������&�HZ4,F/�>/���� �	/�-/?/&/c/J/ �/�/�/�/�/�/�/�/ ?�/;?"?_?q?X?�? |?�?�?���?OO%O 7OIOXmOO�O�O�O �O�OhO�O_!_3_E_ W_�O{_�_�_�_�_�_ d_�_oo/oAoSoeo �_�o�o�o�o�o�oro +=Oa�o� �������� '�9�K�]�o������ ��ɏۏ�|��#�5� G�Y�k�}������ş ן������1�C�U� g�y��������ӯ� ��	��?-�?�Q�c�u� ��������Ͽ��� Ϧ�;�M�_�qσϕ� $Ϲ��������ߢ� 7�I�[�m�ߑߣ�2� ���������!��E� W�i�{���.����� ������/���S�e� w�������<������� +��Oas� ���J�� '9�]o��� �F���/#/5/�G/�$UI_IN�USER  ����h!��  H/L/_�MENHIST �1yh% � (w  �+�/SOFTPAR�T/GENLIN�K?curren�t=editpa�ge,TELEOP,1�/�/?!?�y)�/�%menu�"1133�/}?�?�?γ? �'E?W>71@l?�?O#O5O�(�?W?5k?�O�O�O�O���O�O�O__*_<_ �O`_r_�_�_�_�_I_ �_�_oo&o8o�_Io�no�o�o�o�o�o�� \a�!\o�o/A SVow����� `���+�=�O�� ���������͏ߏn� ��'�9�K�]�쏁� ������ɟ۟j�|�� #�5�G�Y�k������� ��ůׯ��o�o�1� C�U�g�y�|������� ӿ������-�?�Q� c�uχ�ϫϽ����� ��ߔ�)�;�M�_�q� ��ߧ߹�������� ��7�I�[�m���  ������������� �E�W�i�{������� ����������A Sew���<� ��+�Oa s���8��� //'/9/�]/o/�/ �/�/�/F/�/�/�/? #?5? �2�k?}?�?�? �?�?�/�?�?OO1O CO�?�?yO�O�O�O�O �ObO�O	__-_?_Q_ �Ou_�_�_�_�_�_^_ p_oo)o;oMo_o�_ �o�o�o�o�o�olo�%7I[F?���$UI_PANE�DATA 1{�����q�  	�}  �frh/cgtp�/flexdev�.stm?_wi�dth=0&_h�eight=10��p�pice=TP�&_lines=�15&_colu�mns=4�pfo�nt=24&_p�age=whol�e�pmI6)  r3im�9�  �pP� b�t������������ Ǐ��(�:�!�^�E� ����{�����ܟ�՟��I6� � �    �TJ�O�a�s����� ����ͯ@����'� 9�K���o���h����� ɿۿ¿���#�5�πY�@�}Ϗ�vϳ�&� �Ɠs�����)�;� Mߠ�q�䯕ߧ߹��� ����V��%��I�0� m��f�������� ����!��E�W����� ������������:� ~�/ASew�� ����  =$asZ�~� ���d�v�'/9/K/ ]/o/�/��/�/*�/ �/�/?#?5?�/Y?@? }?�?v?�?�?�?�?�? O�?1OCO*OgONO�O �/�/�O�O�O	__ -_�OQ_�/u_�_�_�_ �_�_6_�_o�_)oo Mo_oFo�ojo�o�o�o �o�o�o%7�O�O m����� ^_�!�3�E�W�i�{� �����Ï������� ��A�S�:�w�^��� ����џDV��+� =�O�a�������
��� ͯ߯���|�9� � ]�o�V���z���ɿ�� �Կ�#�
�G�.�k�ޟ�}�|ϵ����������)��4ߧ�#� `�r߄ߖߨߺ�!��� �������8��\�C� ���y������������������$UI�_POSTYPE�  ��� 	 �s�B��QUICKMEN  Q�`�v�D��RESTORE �1|�� � ������������mAS ew�,���� ��+=Oa n�����/ /�9/K/]/o/�/�/ 6/�/�/�/�/�/�? ?0?�/k?}?�?�?�? V?�?�?�?OO�?CO UOgOyO�O6?@O�O�O .O�O	__-_?_Q_�O u_�_�_�_�_`_�_�_ oo)o�O6oHoZo�_ �o�o�o�o�o�o %7I[�o��x����SCRE���?��u1�sc��u2�3��4�5�6�7r�8��sTATM��� ����:�US#ER�p��rT�p�Sks���4��5���6��7��8��B�N�DO_CFG a}Q�����B�PDE����No�ne��v�_INF�O 2~��)���0%�D���2�s� V�������͟ߟ� �'�9��]�o�R����z��OFFSET' �Q�-���hs ��p�����G�>� P�}�t���Я��׿ο ����C�:�L�^� �����͘���
�����av��WORK �!�����.�@����u�UFRAME�  ���RTOL_ABRT�ߜ���ENB�ߣ�G�RP 1�����?Cz  A��� ���*�<�N�`�r�֐�U�����MSK  �)���mN��%!��%z�<���_EVN�����+�ׂ3�«
� h�UEV���!td:\e�vent_use3r\�u�C7z��ϲjpF��n�SPs��x�spotwel=d��!C6��������!���G| '��5kY��� ��>��� 1�Ug���/ ��	/^/M/�/-/?/ �/c/�/�/�/�/$?�/�H?�/:J�W�3������8C?�?�?  �?�?�?�?O+OOOO aO<O�O�OrO�O�O�O �O_�O'_9__]_o_�J_�_�_�_�$VA�LD_CPC 2=�« �_�_� w��qd�Rߠ*o_oqo��hsNbd �j�`��i�da{�oav �_�ooo3BoWi {�o�o�o�o��o� PA�0�e�w�� �������� (�=�L�a�s�
����� ��ʏ�����$�ޟ H�:�o���������ڟ ؟����� �2�G�V� k�}�������¯ԯ� ����.��R�S�y� �Ϛ����������	� �*�<�Q�`�u߇ߖ� �Ϻ���������&� 8�M�\�q���߶� ��n������"�4�F� [�j����������� �����!0�B�Wf� {����������� ,>teT� ������/ +/:La/p�/�/./ �����//'?6/ H/?l/^?�?�?�/�/ �/�/�/?#O�?D?V? kOz?�O�O�?�?�?�? �?_O1_@ORO9_vO w_�_�_�O�O�O_�_ _-o<_N_`_uo�_�o �o�_�_�_�_o&o ;Jo\oq�o��� �o�o�o� �"7�F Xj�������� ���!�0�E�T�f� {�������ßҏ��� �
�,�A�P�b����� x�����Ο����� (�*�O�^�p������� ��R�ܯ� ��Ϳ6� K�Z�l�&ϐ��Ϸ��� ؿ���"� �2�G��� h�zϏߞϳ������� ��
��1�@�U�d�v� ]�ߛ���������� ,��<�Q�`�r��� �����������&� ;J�_n������� �������$F [j|����� ��0E/Ti/ x��/��/�/�/� //,/.?P/e?t/�/ �/�?�?�?�?�/?? (?:?L?NOsO�?�?�O �?�O�OvO OO$O6O �OZOo_~O�OJ_�O�_ �_�_�O_ _F_D_V[��$VARS_C�ONFIG ���Pxao  FP]S�\l�CMR_GRP ;2�xk ha�	`�`  %1�: SC130E�F2 *�o�`]T�dVU�P�h`�5_P�a?�  A@�%pp*`�Vn No9xCVXdv�p�a��<uA�%p��q�_R��_R? B���#�_Q '��H��l�;���{� ����؏ÏՏ�e�� D�/�A�z�-�����dd�IA_WORK +�xeܐ�Pf,		�Qxe���G�P ���YǑ�RTSYNCSE/T  xi�xa-��WINURL ?=�`�������य��ȯگSIO�NTMOU9�]S�d� ��_CF�G �S۳ȿS۵P�` �FR:\��\D�ATA\� �߀ MC3�LO�G@�   UD�13�EXd�_Q'� B@ �� ��x�e_ſx�ɿ�VW� � n6  ���VV��l��q  =�̡�?�]T<�y�Y�T�RAIN���N� 
gp?�CȞ��T�K���b�xk (g�����_������� ��U�C�y�g߁ߋ���߯������_GE���xk�`_P�a
�P�RꋰRE�q�xe*�`hLEX乓xl`1-e�V�MPHASE  �xec�ecRT�D_FILTERw 2�xk �u�0����0�B�T� f�x�����VW������ �� $6HZl�_iSHIFTME�NU 1�xk
 �<�\%����������= &sJ\��������'/�	LIVE/SNA�c�%vsfliv\��9/��� 7�yU�`\"menur/�w//�/�/������]��MO��y��,5`h`ZD4�V�_Q�<��0��$WAITDINEND���a2p6OK  ��i�<���?S�?�9T�IM�����<G w?M�?*K�?
J�?
J<�?�8RELE��:G�6p3���r1_AC�TO 9Hܑ�8_<� �ԙ�%�/:_af��BRDIS�`�N��$XVR��~y��$ZABC�b;1�S; ,��j��I�2B_ZmI1�@V?SPT �y��e.G�
�*�/o�*!o7o�WDCSCHG �ԛ(��Pn\g@�PIPL2�S?i��o�o�o��ZMPCF_G 1��ii�0'¯S;HMs�S��i��p'�c�g��e2���  ��oO3��2x?�  3b�Q@��q�u�� �1�oAD/  �� Ce��1��q�� �>�����F�y����c��@,� ��������� "�Z�~���Ï�>�?�3��´ԏ� ӈ*���*�@�N�x���>���?E��B��l=ڄ��?��?R&�~?s����I�E=�uD_��zC��D5��9��6��>3ȷ�>�&�6��@�y�
y��ŭ�glp����o�_CYLINuD�� { Х� ,(  *=��N�G�:�w�^����� ��ѯ���7���� <�#�5�r��������� ��޿y�_����8�� ��nπ�㜻ã wQ �5�����S������(�ٻ�X�ז�r�A��SPHE_RE 2���ҿ ��"ϧ������P�c� >�P�̿t���ߪ�� ���'���]�o�L� ��p�W�i���������l���PZZ�F �6