��  �"�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ������CCBD_�DATA_T � <$CO�MMENT �$IMCMF_�CF  NE�NDWTWCWFkDBWCd	FGW�TOOL_NUM�W w   qN�~ _FR�w �TRQ��GAIN�$T{DC�$CJI �� T�$DSR`��	I VP�AA�CTL_�TI�$MOV�E_L�WG@D�RARHY& {�/PARM9� �N PEQE} ��K�D&��3�K�K�D_M����3�h�+ �F�STd��|SU�  � L$L�IMIT� �$INSERT_�DIhx$�AM�_F Us"SRBPҎ)P�'|I3/�bBNR x �_d�!B=�'TE0��$b�!ALr�"�AE�'FV��#T�9�v!A2U�(UNJ8V� TVh5Uq8�GRAPH�'RE�TRYS�<1�<2~WEC_DDE&x� �1�7A_PO�0��2AN� �5#��TWL�3ALLT�0�VV'@�!�$VCp27@�2�$�2Ar6@LhP�HD_RA�X`ED�sAheA�GO"�@�� I�DVA_SWG2�@��Ah�@5EhA� LE� �D�MC�ORWPH��!-ASDFW�FY_j"�CP�APz1QTN_S�#�CNGFh$M�IN�@�"?A_ML�_LM�VEL_�CNST�C$AUT_RVbUnPk@3_TL�0TH�1�T��1XSRUDAMP_��O|PS OLSTOP_THRE�1�TAV~Ub �P�D�SRAA�TM�Y��V��QATTOSC_GGDW�E*e#lR�FORCE_O�u MOF\eeI ��LSU�TJUT�fRO�T� C�1� CRE�W~#u �a�eCHG�ZQ�D�dDP@�cV��P��aR�1-AINISH�s�I�`_q�D�a^W�SoT@u|�WZPOCITYjmZP�CNm D�0�Dv�Pdv� �#]#e/w/�/�/�'� 5� ($WO�R� 2�V ' )�2U"�q�ST�P ��pCH�B�rY�#RV^��g�N�Y��FtY�ACTY�C`WA�w��3e�_M���DCPdY�V�e�V�����WQ���^�8��^Q��RTN|ac��T����a�rALGwO_Sxr$P�1��tr�REV_I�T�1�MU�D�0CaCI�!8R��XI��gGAM ![AAS��vє_O@NTR�vYF�`�TR��V�CNPFv�?P�$�.lDCNC0M[ �Z�`O�CHQ�L��Y�F'�l�5�^�OV�M)�QL����IO£�D�A��b���JTH^QPA�V䥽��PDA�pc��DS�PPCCNMONL	S�$�T�1 �T�yV�@J�KPGRC�d�RG�1o��dr�RRo�O�sa�T��O�"_�Rp2�ٽV�-���PDU2CCNAgGWA�g�TH�SǱA-�M�S?ǖS�CVRS1]���a�M۵8a�82�OVK�v���P'���5���VLX����TCI���Y��TRS?`Vo�MG �CCQi��T(�s12��INDEmA�`TM�3P�fT�CC��T�R=G=�USPF8w�p���k@��TWD����f��SR۵��1D��ի����E^PK�PP�Z��CAXCP_P0�B�L��SR���#DI1��?PZH�5��&�RTY��LU�FFIXE�CREAG�Q+u��࿣F�p�q�P+CM�r��CN3FCf��EN� 2����Vѐ��RT�V��TMU��RG`��T����DU%�B�T9�?���Sm��`�P7�`�b�`�IP�)��APf@y���V����Ne�� P�M`����砣���RCh�Pe���7�PS H��(�PYC)���C(L\�p�   }_jQ|^0�! EQ}D=�MVROU2��PERIOF31P����2D'��2�TU�_D���Hǔ���T����K�	5K��K�CL����*aADJ�Q_U^Bq�AaPT�b>�2>REP�r<�]�?Wm rq$�DL�W��M��M��0�'���lB)� ��'#*�F#<+(e#�VL��#z*���#�+(�#z*�P_)B���2
�A�-�x�,� �,OVER�D&�"IB]PGFQ�L9D L9���0PCZb�CFR~7�@D�@C5P��MN1�6�q�12�>UF�p�;TOO�U@�0_T�1�5N'�H?QOR��t2p ALsoG��&�KE��e�&S��AUX�BD� 4?$IMCM�P�r���;� q�@��AUXo_AXS�� ��{C�p` 	 h�@PEx`���D ^c�Cޣ�C^a�C�X�GDXz`����
�j �XAXI@ 
 Td��Db�E�eyA~@{@ pQ�PvR	$IrX�P�V�
�S��GRN��H $�1E_U�p��T�2�Q�05��;��rE���Vk oD�ON�QVa� R_�PKG�RqP � |R`pQS`��Qb�Qb�P%d`�D`%`$�iKa^��`FL~��&pLT�P��ea���c�b���a$�DYN�E$J ugGB�g	�d��d��	PQ<CQxP
 �$Ґ  ���q�d &d  &�`:0S�IONx�  XKqIR�TUALq�SC�OM ?&x&� 2 qv|t �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�J�Uu�P�11 3c{�xd 1pJ���G����  ���� �?�  ŵ��A�   յ��ĺŹ@@ǻ��
��=�C��� B�߲Cʮ����-χ�Y�����F@y ����=�������Dz  ������P��C�`����P�m�"�~�������ǿ ٿ���������E�W� i�{��ߟ��������� ��?��/�A߂�&��� ����+�����	���P��
�y�A���@���Т��d ��w�B�HԖЉ�Y���\�  �� ���#	B��?*	���҄����#W�v��>���Qh����pp� �'8[P2Kt����� ��//��7.� ��A]/���ݱѕ/3 ��|�Z��/�/??+6����F7�/�)�r7^	�>��?l��	�N�5>L���?�1N��"U�<#�
q��p�?92�886a"��	�� ��5QB���5@���4 ��}Ol4���F�M��e�B��5:� _!_�3__W_i_|���=�uB�4!??�_�#�It$ �_$B>%��2
�_gA�$o�_-o�_�VR0+��=�ye.����eQ1�$敕�e(4$�ܡeYokk;��.��e>��H�e�a5����e8M�Y�eY-=�0uQ2>"�7I[m��w
 ?o������� >�P�b�5o��}�����������	ӏ(�� L�7��ow������� ԟ�O���Y�k�}ߏ� �߳�E_����{��� 1ﯯU��y���� ��������=�O� �s�}�;�M�n�ͯ߯ �_��g�9�K�]�o� �ϓ��������-ߣ� �?_��߃��������� ��K�%7I�� �O��ɿW��b� t�������EW���� (:L^p� ����A/S/e/w/�/ �/�/�ˏQcu� =?O?a?s?�?/�?�? �?�?�?/O�/9OKO ]OoO�/�O�O?�O�O �O��y?�?�?�?�?�? }_�_�?�!Og��_�_ o/O%O�OIO�oyo�o �o�O�o�o�o�o	 -�_�_�_�_�_o/� 4ooXojoQo�ouo�o �o�o�O�o�o' Tfx;����[� �[O��,�>�P�O? ����տ���'�/� �?��?�ߥ���s� ��������+�)�O� a�3�������ˏݏ� ����ɯ7�I�[�m�ۯ ��㟵�ǟٟ�1�� !�3��ߓߩ�����'� d����#�5�c�Y�k� }������N����� ���1�ӿU������ �&�����\�n��� ������������ ������; �����������/��� ��/��%/7/=�[/ m/��/�/�/�/�/ t?!?3?E?W?i?� �/(//L/^/�?O �/�/�O�eOwO�O�/ �/6?�/�O�O__S? =_O_a_s_�_�_�_2O DOVOhOzO�o/?�O�O �O�O�O
_�O._@_R_ %?v_m__�_�_�_�_ ��_oo<o�]o� �o�o�o�o�og�y��o �c�u�C��;/q� ���;�M�_� q���������ݿ�� #5GYku�3� y���ˏE����� 1�C�U�g�U�����_� ��ω�3�E�W�a�{� �ϟϱ���1������ �/�A�ʿi�w߉ߛ� ��O���Z�l�~ϐ�+� ��O�������� �2� D�V�h�z��'�9�K� ]��߁��������7� I�v�m�#5#�Yk �������� 1CUg��� ��ͯ��_q� -/���u/�/y� A?C�/#?�� E_?q?�?�?/�?�? �?�?OO%O�/�/�/ �/�/_?,??P?7? t?�?m?�?�?�?��? �?�?OOLO^O!o�O mOO�OSo�Owo __ $_6_H_�o�o������ ����w�_�_ oo� ����o��ɟ۟ퟣ_ �go5�/�Y�{_Mo�_ �_�_�_�o��./o AoG�wo�o�o�o�o E�'��og�y��� �����J����	�� -�?���c�u�W����� ��܏U�j��Ϲ�;� ��֯�����Ϲ�+� T�f�x���������ҿ ����ߣߵ������� ���7O-O������ �ϟ��7�����p�� �/�A�S�e�w����� ������k�}�+ m�O�������2� D�V�����Ϟ���O ]���
��=� ��/G5/G/Y/k/ }/*<N`r �?�}�����  /&/8/J/S/�/w/ �/�/�/�/�O�/�/"? ?�U?�O|?�?�?�?��=�$CCSCH�_GRP12 3�����1&� x�� o_5�Yk^O�!� �O�O�O����O1� ��U�g�y���_���� ӏO�OZ_LObOpOz_ 8oJoko�O�O�O\o_ $_6_H_�_�o�o�_�_ �_��:�)�;�� xoq�����SϹ�H�ݟ ��%�7���[�� ��T��_�q����� ��!�3�ɟ���%� 7�I�[�m�����o� /�֯\�e�{ω�0�ҏ �/i�`�r����+�6� O�a�υߗߩ߻��� ���߀��'�9�K�� 䏁������H�v� ���ߌ�����Y�k��� ��9�7a?������>� ��F���Ugy�� �����	���� ������/1A gN�r����� ��$Qcu ?����.��/ /)/;/M/��?_/�_ �_�_oo,o��?? ��o�o�o(?�o �o (~?LF�p�/ d?�/�/�O�/�?�O�O �OF?X?j?�O�?�?�? �?�?�?._OO0O~ p/�_oJ��ao��  �2�`�V��oz����� ��Xo
�����BO �_R�����#��� ПY�k�}�������ŏ ׏���:_��̯ޯ ����&�8��Dʟ ܟ����ȿڿ��� ��"�4�F�X�jϋ��� ���������q�0�� ��B�T�f�,o��%� �I�[����h���� �b�t��Ϟ�3��� 4�����L�:�L�^� p�������/�A�S�e� w����������� ���+�=�O�"�s�j� |������������  9�Z�ρ�� ��ȿv/�NO`OrO ���O�O:π>�po� ��J_\_n_�_�_ �_��_�_� 2 DVhr/0?B?�� ��T?
/\/./@/R/ d/�?�/�/�/�_o"O 0oBo�O�Oxo�o�o�o �o�o�o�o,> �_bt�_��LO� Woio{o�o�o:�L��o �o�o/ASe w�$�6�H�Z�p�~� ���/��=�4�F�s�j� �2��V�h�z�o�� ���Oԯ�o�
���.� @�R�d�퟈������� п⿘On�������ů ׯrτ���>�l�� ���l����>�\�n� �ߒ�̿���������� �"�Ͻ�������� ��)��M�4�]߃�j� �߹��ߞ�������%� �I�[�F<��|�� P��t���!�3�E� ��P��?�/�/��? ������{�l?~?�� �?�?�?�?�?�t2O ,oVO+���������� �����,>D� /������� �vO�O?�O�O ���O__*_X_�? `_r_�_�_�_�_CO�_ �_oo&o�/Jo�O�O �O	_�o_�oQ_c_u_ �_�_�_�_�_�_�_� ����\o��~ 0��_�o�o�o�o���� �oҏ���,�>� P�b�t���������Ο ��i���(�F?L�^� ؏���� �A�S��  ��o������Z���~� ������ؿ���� ��2�D�V�h�zϐϞ� '�9�K�]�o��ߓ��� ��ɿ������#�5� G��P�i�tφϘ��� �Ϛ�������1���R� ��yߋߝ߯���\�n� 4/x/j<���f� x����/��0/B/ T/f/�/��/�O�/ �����*�<�N�h� (�������:��� �&�8���n����� �/�/~(?:?�V p?�?�?�?�?&/�?�? �O$O6OU�/�/~O �O2�O?O?a?s?�?  _2_�?�?�?�?OO 'O9OKO]OoO
oo.o DoRodozo�o_�Ϧ� G_>_P_i_*�_N `�_������ ���&�8�J��_�_ �������oȏ�T* �j���j�x_n_ �6�`�֟_�����z� $���T�f�x������� ��ү���|������� ǟٟ�
�����E� ,�i�P�y�����ï�� ̯����/�A�S�� w�b������οl������+�<��$CC�SCH_GRP1�3 3����^�&� xn�߮������ �����4�bt �%ߪ���� {�("?L��a����� �����߱�����C�U� g���ߝ߯���g�Y� +�	��-�Zl�� ��^����/�O 2/�V/h/�/�/�/ .�/~�/���.?� ��/ /�?�?B/h/ z/�/�/�/�/�/�/�/ 
?��O�OO?��O�O _�?K ��?�?�?O �_�_�?�_�_�O�_o "o4oFoXojo�O�o�o �o�o_]�o0 B�_�_O"ooFoXo ��O	O�o��ڿP� �ot��o�oQΏ�� ���(�:�L�^�p� ��,�>�P�b�t����� ��������Ǐ��(� :�L�;%�g������� ʟܟ����6�!� �i�~�������Ư}_ s�دK�]�o���� 7o}���m���#��� G���k�}��������� ����ݿ/�A��e� o�-�?�`߿�ѿ�Q� �Y�+�=�O�aϧ߅� �ϩ�������OQ ��u�����=� �);��_q �����I��Tfx ��7/I/��� ,>Pbt��}� 3?E?W?i?{?/�?�? ���C/U/g/�//OAO SOeOwO ?�O�O�O�O �O?_�?+_=_O_a_ �?�_�_�?�_�_�_�� kO�O�O�O�O�Ooo�o �O�/_Y��o�o�o!_ _�_;_�k}��_ ��������o �o�o�o�o!�& J\C�g��� �_�����F�X� j�-���y���M�ӏM_ ����0�B�AO�x� ������/�!߳O�� �O�����e����� �������A�S�%� ��������ϟ�믩� ��)�;�M�_�Ϳ��կ ����˯ݯ#���%� s��ϩ���V��� ��'�U�K�]�o��� ������@�����v� #��G�������� ��N�`�r������� ������������ ���	/w�-/�� ����?�/��/�/ �/��?)?/�M?_?� �?�?�?�?�?f/O O%O7OIO[O��/? ?�/>?P?�O�O�?}? �_�W_i_{_�?�?(O �?�_�_�_oEO/oAo Soeowo�o�o$_6_H_ Z_l_�!O�_�_�_�_ �_�_�_ o2oDoOho _oqo�o�o�o�o���o 
�o.ɏO�v� ���Y�k���U� g�5��-?c�u��� �����-�?�Q�c�u� �폫ϥ��Ϥ��� '�9�K�]�g�%�k��� ����7������#�5� G�Y�G�}���Q���� {�%�7�I�S�m�ߑ� ����#��������!� 3��[�i�{���A� ��L�^�p߂����A� ������ ��$�6�H� Z�l�+=O�� s����w�)�;�h� _�'�K]��� �������/ #/5/G/Y/�}/�/�/ ���/�/Qc�?y ��g?y?k��3O5/ �?/�?�//�/7/QO cOuO�O?�O�O�O�O �O	__�?�?�?�?�? oOOOBO)OfOxO _O�O�O�O�/�O�O�O �O_>_P_t___q_ �_E�_i�_oo(o :o������㟵� �i�o�oa�s��� ����ͯ߯�o�Y '�!�K�mo?�o�o�o �o����� �!39� ��i{���7�� ���Y�k������� ��<�Ϗ�����1� ��U�g�I��ϝϯ�Ο G�\���	߫�-߄�ȿ ڿ����߫��F�X� j�|ώϠϲ������� ������������ ��)__�߷����ߑ� ��)�����b���! 3EWi{��� �]�o��_�A ����� ��$6H ����ߐ�/�_O/� s/���/�/�/�/ ?9'?9?K?]?o?� 
//./@/R/d/�O�/ o/�/�/�/�/�/�/? *?<?E?r?i?{?�? �?�?�_�?�?O�?��GO�_nO�O�O�O�M��$CCSCH_G�RP14 3�����A&� x�ao'� ��K�]�P_��z_�_ �_ۏ����_#�u�G� Y�k�}��_����ş_ �_Lo>_T_b_lo*< ]�_�_�_Noo(o :o�o���o�o�oӟ �,����-�׏jc� u���E߫�:�ϯᯋ� ��)���M���q�� F���Q�c�u������ %ϻ�����)�;� M�_�q���z�!�ȿ N�W�m�{�"�ğ�?[� R�dϑ���(�A�S� ��w��������� r���+�=���֟s� ��������:�h�ϛ� ~����K]�ς�+� )SO�s��0���8� ��GYk}��� �������� ���/#
3Y@ }d������� ///C/U/g/	O�/ v/�/�/ �/�/	?? -???���OQ?�o�o�o �o���?O�x ��O����� �pO>�8�b��?VO�? �?|_�?�O�_�_�_8O JO\O�_�O�O�O�O�O �O o�O_"_p�b?�o <�ʏS� ��$� R�H��l�~������� J���s��4_�oD� ͏ߏ�����¯K� ]�o���������ɟ۟ �,/�_����п��� z��*���6/��ί� ��Ϻ�������y�� &�8�J�\�}���	Ϥ� ������c�"��v�4� F�X�������;� M�����Z������/T� f�x��ߐ�%��&�� ��>�,>Pbt ��!�3�E�W�i�{� ��������������� /A�e\n� �����/�+ �/L��s���� ��h?�@_R_d_���_ �_,�r/0�b�
/�/ �/<oNo`oro�o�o�/ �o�o�/ //$/6/H/ Z/d?"O4O�/�/�/�/ FO�/N? ?2?D?V?�O z?�?�?�o�o_"4 �_�_j|���� �����0��oT� f��o����>_��I[ m�,�>���� ��!�3�E�W�i�� �(�:�L�b�p����? ��/�&�8�e�\��$� �H�Z�l������_ ƿؿa����� �2�D� V�߯zόϞϰ����� �_`�����v���ɿd� v�����0�^������ ^�ϡ�0�N�`�r�� �Ϩ���������� �߯���������� �?�&�O�u�\��� �����������;� M�8.���n���B�� f��%7�� B|O�?�?��O��� �m^OpO� �O�O �O�O�O�f$_H_ /|������ �/�06/�/
?x ������/�/ �/h_z_�?�_�_�/�/ �_�_
ooJo�ORodo vo�o�o�o5_�o�o�o �?<�_�_�_�_ �o�CoUogoyo�o �o�o�o�o�o������ ��ȏN���p/"��o ���������ğ ֟�����0�B�T� f�x���������ү[� ����8O>�P�ʟܟ �����3�E���� r��Ϯ�Lώ�p����� ��������� ߆�$� 6�H�Z�l߂ߐ��+� =�O�aπ�ϗ�~ϻ� ���������'�9�� B�[�f�xߊ߷��ߌ� ������#��D���k� }����N`&/�/ j?\/.��/�X�j��� �/�/�/|�"?4?F?X? �|?���?�_�?��� 
��.�@�Z� �����,���� *��`r��?�? 
/p/O,O�/HbOtO �O�O�O?�O�O�/_ _(_G/�?�?p_�_$/ �_�?AOSOeOwOo$o �O�O�O�O�O__+_ =_O_a_�o 6D Vlz o�ߘ�9o0o Bo[o
���o@�R��o v���������Џ�� ��*�<��o�or��� ������/F��y�\� ������\�jo`o	�(� R�ȯQ��u�l���� F�X�j�|�������Ŀ ֿ�n���������˯ ݯ������7��[� B�k������������ ���!�3�E��i�T� ��x�����^��������.��$CCSC�H_GRP15 �3���P��&� x `/��r����� �����&�Tfx� ������m�/ O>/��S�������� �������5�G�Y��� }����Y�K�� ��L/^/��/�/ P���/�/ ?�_$?� H?Z?/~?�?�? ��? p/�?{/� O�/�/�/  ??�O�O4?Z?l?~? �?�?�?�?�?�?�?�� �_�_AO��_�_�_�O =/��O�O�O
_�o�o �O�o�ov_�o& 8J\�_���� oO/���"�4��o �o_�o8Jď֏ _�O�����B��f� ���C���ҟ��� ��,�>�P�b�t�� 0�B�T�f�x�v����� ��ҟ����ݟ�,�>� -��Y���}�����ί ூ���(����[� p���������ooe�ʿ =�O�a�s�����)o� ��_����9� ]o���Ϸ�/� ����!�3���W�a�� 1�R������C���K� �/�A�Sߙ�w߉ߛ� �ۿ����_C��g y����/�� 	//-/��uoc/��/ ��;��/FXj|� )?;?����// 0/B/T/f/��o�%O7O IO[OmO�/�O�Ox/�� 5?G?Y?�?!_3_E_W_ i_�?�_�_�_�_�_�? �_�Oo/oAoSo�O�o �o�O�o�o�o��]_~_ �_s_�_�_as�_w? oK����o	o�o -o��]�o����o���� ɏۏ������� ������<�N� 5�r�Y��������oޏ Տ� ��8�J�\�� ��k���?�ş?o��� �"�4�3_�j����� ��?��_믩_�� �/����W��������� ����3�E��y��� ������ӯݿ�ϭ�� -�?�Q���u�ǿ���� ��Ͽ����e�w� �ߛ����H����� G=Oas�� �2���h��� 9��������
�� @Rdv���� ��}/�/�/�/�/�/ �/�/i�?���� ��O�?��?�?�?�� 	OO!�?OQO�/uO/ �O�O�O�OX?�O__ )_;_M_��?�?O�? 0OBO�_�_xOoO�oן Io[omo�O�O_�O�o �o�o�o7_!3EW i{�o(o:oLo^o }�_�o{o�o�o�o�o �o$6	_ZQc ���������  ���A�ߟh�z����� ��K�]�����G�Y�'/ }�OU�g�������� y��1�C�U�g���ߟ �ߗ��ߖ�����+� =�O�Y��]������� )������'�9�K� 9�o���C�����m�� )�;�E�_�q����� ���������%��� M�[�m����3ϵ�>� P�b�t���3���� ������(�:�L�^� �/A��ew 鯛i�-ZQ/ /=/O/ws/�/�/ �/�/�/�/�/??'? 9?K?�o?�?�?�Ϸ? �?C/U/v/Ok/�/�/ YOkO]�/%_'?�O? �Or??{?)?C_U_g_ y_�?�_�_�_�_�_�_ 	o�O�O�O�O�O�o�O _�O4__X_j_Q_�_ �_�_�?�_�_�_�_o 0oBo�foQoco�o7� �o[��o�o,Ǐ ُ��q��կ���[/ ���S�e�w���� ����ѿ���K��� =�_1�����ӏ ������%�+���[� m������)��ُ� ��K�]σ�鯓ϥ�.� ���������#ߑ�G� Y�;�}ߏߡ���9�N� ���ߝ��vϺ����� �ϋ���8�J�\�n� �ߒߤ߶�����u��� ������������y�o o�������� ��T��%7 I[m���O� a���/Q3/��� ���(:�/�� ���?�oA?�e?� ��!/�?�?�?�?+/ O+O=OOOaO�/�/?  ?2?D?V?u_z?a?s? �?�?�?�?�?
OO.O /7OdO[OmO�O�O�O �o�O�O_�Os/9_�o�`_r_�_�_�]�$C�CSCH_GRP�16 3�����Q&� xٯS��=� O�Bos�lo~o�o͟ ߟ�o�g�9�K�]� o��o���Ϸ��_�o> 0oFoTo^�.�O��o �o�o@��o,� ď��t��ůׯ� ����ɟ\�U�g�y� 7,���ӿ}���	� ϙ?��c���8��� C�U�g�y����߭� ӿ���	��-�?�Q� c�u�l����@�I� _�m�߶��OM�D�V� ������3�E���i� {�����������d��� /��ȯew� ��,�Z��ߍ�p��� ��=O~�t�/E_ �e�"�*�9/ K/]/o/�/�/�/�/�/ �/�/������ �?/�%/K/2/o/V/ �/�/�/��/�/�/�/ ?5?G?Y?�O}?h?�? �?�?�?�?OO1O ���_CO����� ����O�O؟j�|��� _���֏����b_ 0�*�T�vOH_�O�Ono �O�_�o�o�o*_<_N_ �or_�_�_�_�_�_ �_oob�TO� �.� ��E������D�:� ��^�p�������<��� ܯe� �&o�6���џ ��������=�O�a� s���������ͯ߯? �o�ϰ�������l�
� ��(?����ҿ���� �߾�����k���*� <�N�o�r��ϖ��� ��U���h�&�8�J� �����	���-�?��� ��L��~��?FXj ��������� 0�0BTfx� %7I[m�/� x�����! 3�WN`y�� ���?��/�?>/ ��e/w/�/�/�/��ZO �/2oDoVo��zo�o� d?"�T���/v?�?. @Rdv��?�� �?�/??(?:?L?VO _&_�?�?�?�?8_�? @OO$O6OHO�_lO~O �O��o�&��o�o \�n���������ȏڏ ����"��F�X�� |���0o��;�M�_�q� ���0���ˏݏ�� �%�7�I�[����� ,�>�T�b�t��O��!� �*�W�N� �� �:� L�^� ��ϔϚo���� S���|��$�6�H�ѿ l�~ߐߢߴ���|oR� sυ�hϩϻ�V�h��� ��"�P/������P��� ��"�@�R�d�v��ߚ� ������������� ������������1� �A�g�N��������� ������	 -?*/  u`�4/�X/� �)�/�/4n_ �O�O���O����_ P_b_x��_�_�_�_ �_v/X/o�:o?n ������/�?�/ /"/(?�?�?j/|/�/ �/�/�/�?�/�/�?Zo lo�O�o�o�?�?�o�o �o<�_DVhz ��'o����
� �O.��o�o�o�o���o ��5GYk}�� ���r��������� @�ޟ�b?������ ӏʏ��������ȯ�� ����"�4�F�X�j� |�������ĿM���� �*_0�Bϼ�ί﯊� �%�7�����֏d��� ��>߀�b��z����� ��������x��(�:� L�^�t����/�A� S�r�w߉�p߭ߔ��� ������+���4�M� X�j�|���~���� ����6��]�o��� ����@R?�?\ON?  �r?ԯJ\}�?�? �?nO&O8OJO nO ��O�o�O�����  2L�/��� �/���
�/ �/Rdv�O�O�/b? __�?:/T_f_x_�_ �_
O�_�_�?�_oo 9?�O�Oboto?�o�O 3_E_W_i_�_�_ �_�_�_�_oo/oAo So� ��(�6�H�^� l��o���+"4M ����2�D��h�z� ������ԟ���
� �.���d�v���ʏ ��r?8��k�N����� ��N�\R���D��� C�޿g�^����8�J� \�nϤ��Ϥ϶����� `�u���������Ͽ�� �ڿ�)��M�4�]� �ϕϧ�z��������� �%�7���[�F��j� 쯲�P�������� ���$CCSCH_�GRP17 3����B�?&� xR?�� �d/�����~��� ���F/X/j/	��/�/ �/�/�/�/_�?_0? s�E����������� ��'�9�K��o��� ����K=���� >?P?���?�?B/� �?�?�?�oO�/:OLO �/pO�O�O��Ob?�O m?�_�?�?�?�?O ~_�_&OLO^OpO�O�O �O�O�O�O�O�zo�o 3_�/�o�o�o�_/?� �_�_�_�_v��_� �ho����*�<� N��or��������oA? ޏ����&����_ ��*�<���ȟ�_�_ ������4�ޏX����� ��5���į֯���� �0�B�T�f��"�4� F�X�j�hώ�u���į ���ϯ��0��	� K�x�o�������ҿt� ����ϋ�M�b�t� �ϘϪ�aW��/A Sew��a�s�Q/ ����+}Oa s��ߩ�?����� �%���I�S��#�D� �ߵ���5���=��!� 3�E��i�{����� y�o5/�Y/k/}/ �/�/�/!�/�/�/? ?�gU?�y?��- �?8/J/\/n/�/O-O �/�/�/�/�/?"?4? F?X?��a�_)_;_M_ __�?�_�_j?��'O9O KOxOo%o7oIo[o�O o�o�o�o�o�O�ot_ !3E�_�{�_ ����Oopo�oeo �o�oS�e��oiO�o=� ��я��o��� O�a�s��������͟ ߟ��������ԏ ��
��.�@�'�d� K�������Пǟٟ ���*�<�N��r�]� ��1Ϸ�1ޯ��� &�%o��\�������? ����oݿ�o�{?u� �Iϧ��������� ��%7	�k�}����� ��ſ�ύߟ���1� Cϱ�gϹϋϝϯ��� �����	�Wi� ���:����9 /ASew��$ ��Z�/��+/� �����/�/2D Vhz����� o?�?�?�?�?�?�?�? [�O�/�/�/�/�/y_ �Oy/�O�O�Oy�O_ �1_C_�?g_�/�_�_ �_�_JO�_�_	oo-o ?o���O�O�O�O"_4_ �o�oj_a_�ɯ;M _�_w_o�_��� �)o�%�7�I�[�m� �,>Po�o �m������ �(��_L�C�U���y� ���������ُ��� 3�ѯZ�l�~�����=� O�����9�K�?o�_ G�Y�؟�����k�� #�5�G�Y��ѯ�� ������/�A� K�	�O��������u� �����+�=�+�a� s�5�����_�	��-� 7�Q�c�u������� ��������?M _q�%ߧ0�B�T� f�v�%�������� ��,>P�� /!/3/�W/i/ۿ�/ [LC�/?� /?A?ie?w?�?�?�? �?�?�?�?OO+O=O �/aOsO�O�ߩO�O5? G?h?_]?�?�?K_]_ O�?oO�_�?�_dO �?mOO5oGoYoko�O �o�o�o�o�o�o�o�_ �_�_�_�_��_o�_ &ooJo\oCo�o�o�o wO�o�o�o�o�o"4 ��XCU�)��M� �������˟�� c���ǿ��M?ÏՏ ��E�W�i�珍ϟϱ� ��y���=���/�Q� #�u�������şs��� ������M�_�q� �������˟ݟ�=� O�u�ۿ�ߗ� ϳ��� �������9�K�-� o��ﲿ+�@����� ���h߬߾�����}� ���*�<�N�`�r�� ������gy�� ����k��� ������u��� F��//)/;/M/ _/q/�/�/�/AS�/ �/?C%?뿱�� �//,/�?����t/ �O�3O�/WO�/�/�/ ?�O�O�O�O?__ /_A_S_�?�? OO$O 6OHOgolOSOeO�O�O �O�O�O�O_ _�/)_ V_M___�_�_�_s�_ �_�_�_e?+o�Rodo�vo�o�m�$CCS�CH_GRP18 3����a�&� x˿E��ݯ/�A�4 e��^p���ѯ� ��Y�+�=�O�a�� ��ߩ��o�0�"8 FP�� �A���� 2�����ď���� f�x�����ɿ�v��� ϻ�N�G�Y�k�)��� �����o�����ߋ 1�ۿU��*���5�G� Y�k�}���	������ ������1�C�U�g� ^������2�;�Q�_� 憎}_?�6�H�u��� �%7��[m ����V��� !v���Wi{�� Lr�b��// A/p�f�?7o�/W �/r�+?=?O? a?s?�?�?�?�?�?�? �/�/�/�/�/�/�O? �/?=?$?a?H?�?�? �?��?�?�?�?�?'O 9OKO�_oOZO�O~O/ �O�O�O�O_#_���o 5_����̏ޏ���� �_�_ʯ\�n����_�� ��ȟڟ���To"�� F�h_:o�_�_`�_�o ���o.o@o�do �o�o�o�o�o��o�o T�F_|�� ���7� ү����6�,���P� b�t�����.���οW� ���(ϱ�ïկ� ���Ϧ�/�A�S�e�w� ��������ѿO��� �ߴ�����^����� O�ϲ����ό��� ����]���
��.�@� a�d��߈�������G� ��Z�*<��� �������1���>� ��p��O8J\~�t� 	��
/���"/ "/4/F/X/j/|/ );M_~?�j� ����//%/�� I/@/R/k/v/�/�/�/ �O�/�/?�O0?��W? i?{?�?�?��L_�?$ 6Hv�l~�VO� F����?hO�O �2�D� V�h�z�xO�����O�? �?OO,O>OH_oo �O�O�O�O*o�O2__ _(_:_�o^_p_�_Џ ��o��v�N�`� r���������̟ޟ� ����8�J�ӏn��� "��-�?�Q�c�u�� "�����ϟ���� )�;�M������0� F�T�f��_���
�� I�@�����,�>�P� �t߆ߌ�߼�E��� n���(�:���^�p� �����nD�e�w� Zߛ߭�H�Z����� B?������B��߅�� 2DVh���� ������������ ���~�����#
3 Y@}��t��� ���1?g R�&?�J?��� 	//�?�?&/`o�_�_ ���_���/�/Q/BoTo j/�/�o�o�o�o�oh? J?�,O`/r/�/ �/�/�/�?�O�??? O�O�O\?n?�?�?�? �?�O�?�?�OL^�_ ���O�O��� � .��o6�H�Z�l�~��� ��Ə؏����_ � ����z����'� 9�K�]�o��������� ɏd�v�������2�Я �TO�ԏ����ş�� r���r������޿� ��&�8�J�\�nπ� �Ϥ϶�?�������o "�4߮����|�ֿ� )�����ȟVϐ��0� r�T���l��ϔϮ��� ����j���,�>�P� f�t����!�3�E�d i�{�b�������� ������&�?�J�\� n�����p������ �(�Oas�� 2/D/
O�ON_@O�dO ƿ<No�O�O�O` __*_<_�`_��_ ~�_��� $ >/�/�/}/~��/? ����/�?v?D/ V/h/�_�_�?TO�_o �O,?FoXojo|o�o�O �o�o�O�o�o+O�_ �_TfO��_%o7o Io[o��zo�o�o�o �o�o�o!3E�� ���(�:�P�^�� ��|���&�?�� � ��$�6���Z�l�~��� ����Ưد���� � ��̏V�h�z�����dO *� �]�@�������@� N�D���6��5��� Y�P�����*�<�N�`� ���ߖߨߺ���R�g� yϋϝϯ��������� ����?�&�O�u߇� ��l����������� )���M�8�q�\�޿���B���������$�CCSCH_GR�P19 3����4�&� xDO��/V? �/�/���/p�����
 8?J?\?���?�?�?�? �?�?Q�?�_"Oe�7 ����������� +=�as�� =///��0OBO �/�/xO�O4?��O�O �O�_�?,_>_�?b_ t_�_��_TO�__O�/ o�O�O�O�O�Opo�o _>_P_b_t_�_�_�_ �_�_�_�l~%o�? ���o!O�߸o�o �o�oh�z��o����Z ԏ���
��.�@�� d�v������3OП� ������ŏ�o��ۏ �.������o�o���� ��&�ПJ���럕�'� ����ȿڿ����"� 4�F�X���&�8�J� \�Z߀�g�������ڿ �����"����=�j� a�sϠϲ���f����� ���}�?�T�f�xߊ� ��S�I���!3EW i{�S�e�C?�� �w�/o/A/S/e/w/ ��/�O�/�߳��� ��;�E�6��� ��'��/���%�7� }[�m���/���k �'?�K?]?o?�?�? �?/�?�?�?�?O� Y�GO�/kO���O*? <?N?`?r?__�?�? �?�?�?OO&O8OJO ��S	oo-o?oQo�O uo�o\O��_+_=_j_ );M�_q� ����_�fo�� %�7��o�m��o���� ��{AbtW�� E�W��[_�/߱�ß ՟�������A�S� e�����������ѯ� ��~�������Ɵ؟�� ��� �2��V�=�z� ����q�¯��˯�� �.�@��d�O���#� ��#�п����� ��Nϝ������O���� ��ύ�mOg���;� �������� )��]�oρϓϥϷ� �������#�5ߣ� Y߫�}ߏߡ߳����� ����I[q���� ,����+/!/3/ E/W/i/{/�/�/�/ L�/�/��?��� ���?�?$/6/H/Z/ l/~/�/�/�/�/aOsO �O�O�O�O�O�OM�_ �?�?�?�?�?ko�_k? �_�_�_k�_�_#o 5o�OYo�?}o�o�o�o <_�o�o�o1�� �_�_�_�_o&o�� \oSo����-�?�Q��o io�o�o����Ϗ� ��)�;�M�_�q�� ��0�B�a��ox�_� ������ҏ������ �o>�5�G�t�k����� ������˟���%�ÿ L�^�p�����/�Aϟ� ��+�=�Oa�o9�K� ʯ�����]���'� 9�K��ÿ��{��z� ٯ����!�3�=��� A�{������g�տ� ����/��S�e�'� ����Q����)�C Ugy����� ��	��1?Qc u�"4FX� h/������ 0B�/�/?? %?�I?[?��?M� />/5/�?�?�!O3O [/WOiO{O�O�O�O�O �O�O�O__/_�?S_ e_w_��_�_'O9OZO �_OO�O�O=oOoA/�O 	_�o�O�oV_�O__ _'9K]�_�� �����vo�o�o �o�oݏ�o�o�o�o <N5r��i_� �����&��J� 5�G������?�ȏڏ ����������U��� �ϋ/��?O��ǟ�7� I�[�ٟߑߣߵ�k� ��/�����!�C��g� y�������e�w����� 	����?�Q�c�u��� ���ϯ�/�A�g� ��w��ߥ������� ���u�+�=��a�s� �����2������� Z�������o��� �.�@�R�d�v����� ����Yk}��� ��]����� �g/y/��/�/8�/ �/�/	??-???Q?c? u?�?�?3E�?�?�? 5/O�ϣ/y/�/�/�/ ??�O��f?�_�� %_�?I_�?�?s?O�_ �_�_�_O�_o!o3o Eo�O�O�O__(_:_ Y^_E_W_�_{_�_�_ �_�_ oo�?oHo?o Qo~o�o�oe��o�o�o �oWO��DVhz��}�$CCSCH�_GRP1A 3�����q&� x�� 7���Ͽ!�3�&�W��/ P�b�����ÿտt��� K��/�A�S�ʏw�q� �����"��*�8�B�  ��3�������$�ڏ ��������z�X�j� |��ϻ��h���߭� @�9�K�]���ϥ� ��a�������}/#��� G����}�'�9�K�]� o�����߷������� ���#�5�G�Y�P��� ����$�-CQ��� oo1�(�:�g����� )��M_q�� ��H��//h ��I/[/m//�/> d�qT��!?3?b� X�/�?)�?I/�?/ d//�/O/OAOSOeO wO�O�O�O�O�O{?�? �?�?�?�?�_�?�?	O /OOSO:OwO�O�O�/ tO�O�O�O�O_+_=_ �oa_L_�_p_�/�_�_ �_�_oo��'o�� ����П�����o�o ��N�`�r��o��诺� ̯ޯ�F��8�Zo ,~o�oR��o�|��� �� 2��V�z ��������F� 8on����)�Ŀֿ ���(�ό�B�T�f� xϊ� ����I���
� ��ߣ���ǿٿ뿆� ��!�3�E�W�i�{ύ� �ϱ���_̏���� ����P��� ���_�� �߶���~��������� O����� 2S�V ��z���9��� L�
.�������� ��#��0��b �_*/</N/pf�� �/�/�/�/??&? 8?J?\?n?�	//-/ ?/Q/pOu/\/�/�/�/ �/�/�/??�;?2? D?]?h?�?�?�?|_�? �?O�_"O�IO[OmO O�O��>o�O�(�:� h�^�p�H_8��� �OZ_�_�$�6�H�Z� l�j_����t_�O�O�O __0_:o�o
x_�_ �_�_�_$o�_oo ,orPobotoԟ� ��
�h���@�R�d�v� ��������Я���� ��*�<�ş`�r���� �1�C�U�g��ϝ� ����ӯ���	��-� ?��������"�8�F� X��o|�����;�2� ������0�B��f� x�~����7���`��� ��,���P�b�t��� ����`�6�W�i�L�� ��:L����4O� ��4���w��$6 HZ��~���� ��s�����/ p����%K2 o��f����� �/#/O/Y/D/}/ O�/<O�/�/�/�/? �O�O?R�o�o���o |�?�?C?4F\?�? |����ZO<O� ����OR?d?v?�?�? �?�Ot_�O�?O_�_ �_NO`OrO�O�O�O�_ �O�O�_>�P��ot��� �_�_��Ώ��� �r (�:�L�^�p������ ��ʟܟo����� ��яl�Ꮠ��+�=� O�a�s���������V� h�z�����$�¿ԿF_ ��Ɵx�������d�v� d��Ϭ�ԯ������� �*�<�N�`�r߄ߖ� ��1��������&� �ϲ���n���	�߶� �ﺯH߂���"�d�F� ��^��߆ߠ������� \���0BXf ����%�7�V[�m� T���x����������� ��1<N`� �b/�����/ �/ASew�$?6? �O�_@o2_�V_��./ @/a/�_�_�_R/�_
o o.o�Ro�/vop��o ��/��//0?�? �?o?p/�/�?O�/�/ �/�/ ?�OhO6?H?Z? �o�o�OF_�o�_O 8J\n��_�� �_���_�o�oF� X��O|��o);M ���l����� ���%�7�ҟ��� ��,�B�P�֏xn ���1���x�� (���L�^�p������� ��ʿܿ� �Ϭ��� H�Z�lϮ���V_�� O�2�s�����2�@�6� ߿��(��'���K�B� �~��.�@�R��v� �����D�Y�k�}� �ߡ߳����߾���� ��1��A�g�y��^� ���������	��� ?�*�c�N��ϖ�4����������$CC�SCH_GRP1�B 3����&&� x6_�v?HO�?�? ��?b����*O<O NO�rO�O�O�O�O�O C�O�o_W)�� ���y/�/�/ /�/Sew�//!? �/���"_4_{?�? j_|_&O�/�_�_�_�� �_�Oo0o�OTofoxo ���oF_�oQ_�?�o�_ �_�_�_�_bt
o0o BoTofoxo�o�o�o�o �o�/^�p��O���� ʏq_����� Z�l�w����L�Ɵ؟ ���� �2���V�h� z����%_¯ԯ��� 
�������͟� � ������z�xϢ�� ¯<��ݯ����Ϩ� ����������&�8� J�����*�<�N�L� r�YςϨϏ��ϳ��� �����/�\�S�e� �ߤ߶�X��������� o�1�F�X�j�|��C#5G/�/Q? C/�g/ɟ`�r����/ �/�/��	??-???� c?���?�_�?����� $�6�H�b"��� ���4���� 2 ��hz��?�?/ x/OO�/PIO[OmO O�O ?�O�O�/�O�O _O/�?�?W_i_,/�_ OIO[OmOO�_o�O �O�O�O�O_!_3_E_ W_i_�o�o+= Sao���Ao8oJo co���o'�9��o]� o���������ɏۏ� ���#��o�oY�k�}� ����/N�$���d��� ��ɏC�roho��9� ��Y�ӯ}�t����-� ?�Q�c����������� Ͽv���������ӯ� ��	���?�&�c�J� s���������ƿ�� ��)�;�M���q�\ϕ� �����E�����%����D������x ���o b����,� Zl~���� ���s� /OD/��Y� �߽����������:� ;�M�S�������� ��Q3��%�R/d/ ��/�/V���/�/ ??*?�N?`?c�? �?�?�a/v/�?O� &O�/�/�/??�O�O 7?`?r?�?�?�?�?�? �?�?O|_�_�_�_�_ �_�_�_�O"���O�O �O�O�o�oC_�o�o|_ �o,>Pbt ����w_�_�� �yo:�!�o�o�o >Pb܏__��� ��H��l����I� Ɵ؟���S� �2�D� V�h��$�6�H�Z�l� ~�|�������؟���� ��2�D�V�)�_��� ����¯ԯ毈�
��� .����a��ψ�������8�J�EU�g�y�?� �u�G_���o�Ϥ� ������;M_ qHϕ߹�/� � ��D�V�h�zϔ�B�T� ��������f��.�@� R�d�����߬߾�� �D���3E����{ ����R���� ///A/����/�/ ^��/7{���+? =?��////A/S/ e/w/�/�/O'O9OOO ]OoO�O�O:?����s? j?|?�?#_5_�?Y_k_ O�_�_�_�_�_�_�_ oo1oCoUoO"O�o �o�o_�o���_V_�_ �_�_�_�_u�?�?Co A�k���o��o�oPo �o_�q������o��ˏ ݏ������� ���;�"�4�q�X� ��|���ˏݏ��o�� %��.�[�m��!��� ��ǟ��4��w�!�3�E�W�ѿ�F� �� �ߪ����?2�_+� =�^�����O����� ��
��.���R�Lv� ����ݯ���-��� ��l�m�����ϵ�ǿ ٿ�����e�3�E�W� ������C�������� &8J\��� ��������" 4��X��&8J ��i����� ��"4�/�/�/ �/�/??,?�T�J� ///./�?�?u/�? O�/(O:OLO^OpO�O �O�O�O�O�O�O�/�/ $_6_H_�?l_S�O�? LO/OpO�O�Oo=/3/ �O�o�zo$_�oH_?_ �O{_�o
.�_R dv��AoVohozo �o�o�o���o�o�o
 �o.>dv�[_ ��������� <�'�`�K��_����� ̏ޏ��j�|�G���� ��q�Cߵߧ�y/��-O ğ֟��%�7�I��m� ߑߣ�z���>����� �R�$�v�������Ư t���������N� `�r��������̯ޯ ��/�v���e�w�!� ������������� +�.�O�a�s���,�A� ��������i����� ��]o�+�=�O�a� s�����������GY k�����l� �����U/g/ �/�/G�/�/�/�/	? ?-???Q?c?u?�?B T�?�?�?D/O�ϲ/ �/�/�/	??-?�O� �u?s_��_�?7_�? �?�?O�_�_�_�_O �_�_o!o3o�O�O_ _%_7_I_Gm_T_f_ �_�_�_�_�_�_o!o �?*oWoNo`o�o�o�o S��o�o�o�ofO,��@Sew���H � 2�D�
�ܿN�@�d� �/]�o�����п⿁� ��*�<��`�׏�� ~������!�3�E� _�����������1� �����/�����e� w��������u���� ��M�F�X�j�|ߎ�� ����ǿ�����L��� ��T�f�)����F�X� j�|������������ ����0�B�T�f��� ��(:P^� �o|o>�5�G�`��  ��$6��Zl~� ������/ / ����V/h/z/��/�� K!~a���@? o�e�/O6�?V/�? z/q//�/*O<ONO`O �/�O�O�O�O�Os?�? �?�?�?�?�?�_O�? �?<O#O`OGOpO�O�O �O�/�O�O�O�O&_8_ J_�on_Y_�_}_�/�_�B�_�_o"o��wI �����u��ٟ�� ��_�o)W�i�{� ����ïկ�o��p ��A��oV�o�o�o �o�����7�8JP� ʏ�����N�0� ��"�O�a������ ��S��߿���'� ��K�]�`��ϓϥ�� ^�s�����#ߛ�߿ ��Ϗߡ�4�]�o� �ϓϥϷ��������� y������������ ��__�������߇� ��@����y��� );M_q��� �t���v�7 �������;M_ ���ߧ�/�_E/� i/
�F�/�/�/ �/P?/?A?S?e?/ !/3/E/W/i/{/yO�/ �/�/�/�/�/�/	?/? A?S?&\?�?�?�?�? �?�?�_O�?+OO� ^O�_�O�O�O�O5oGgJRodovo<����r� D���_�_�_��� ��_8�J�\�n�E_�� 	o����ڟ_�_A_S_ e_w_�o?Q�o�_�_ �oco+o=oOoao� ��o�o�o���A��� 0�B��x������� ��O�������,�>� ~��������[���4� x�������(�:�ͯ�� ��,�>�P�b�t��� ���$�6�L�Z�l߂� ��7ϸ?�?p�g�yϒ�  �2���V�h�ߌ�� ����������
��.� @�R��߈������ ����}�S������� ��r�ϗ�@�>hO� ������M���\n ��������� �����? 81nU�y� ������"//+/ X/j/|/O�/�/�/�/ 1�/tO?0?B?T?�O�GK�O�O_�o�� ��/��(O:O[O� ��LO�����? +��OO�I�s��?�O�? �?�?O*_�_�_i_jO |O�_�_�O�O�O�O�O �obo0_B_T_�����o @ɏۏ�o�#�5� G�Y��}������ş ן�����1��oU� ͏�#�5�G���ӯf� ������şן���� �1�����Ͽ��� �)�ЯQ/G/	� �� +�����r���߫�%� 7�I�[�m�ߑߣߵ� �����ߦ���!�3�E� ��i�P���I�,�m� ߑ��:�0�����? w�!��E�<���x��� +��Oas� �>�S�e�w������� ���������+ ;as�X��� ���/9$] H��?���� �