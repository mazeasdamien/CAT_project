��   g�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����BIN_CF�G_TX 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG���DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST�  �DwNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !�� FT� @�� LOG_8	,C�MO>$DNL�D_FILTER��SUBDIRCAPC� �8 .� 4� H{A�DDRTYP�H NGTH����z +LSq� D $ROB�OTIG �PEEyR�� MASK��MRU~OMGD�EV�gPINF�O.   �$$$TI ���RCM+?T A$( /�QSIZ�!S~� TATUS_%�$MAILSER�V $PLAN~� <$LIN�<$CLU��<�$TO�P$CC�&FR�&YJEC�|!Z%ENB ^� ALAR:!B��TP,�#,V8 S���$VAR�)M��ON�&���&APPL�&PA� �%�N�'POR�Y#_�!>�"ALERT�&i2URL }Z3�ATTAC��0ERR_THROU3�US�9H!�8� CH�- c%�4MAX?W�S_|1��1MOD��1I�  �1�o (�1PWD � � LA��0�N�D�1TRYFDE�LA-C�0G'AERcSI��1Q'ROBICLK_HM 0Q'� �XML+ 3SGF�RMU3T� !OU�U3 G_�-COP 1�F33�AQ'C[2�%�B_AU�� 9 R��!UPDb&PC�OU{!�CFO ?3 
$V*W��@c%ACC_HYQS�NA�UMMY1�oW2"$DM*  $DIS��gSM	 l5�o!�"%Q7�IZP"�%� �VR�0�U�P� _DLVSP�AR��QN,�
3 �_�R!_W�I�CTZ_IND9E�3^`OFF� ~URmiD�&f�   t Z!N`MON��cD�.�bHOUU#E%A�f��a�f�a�fLOCAܗ #$NS0H_[HE���@I��/  d8`ARP�H&�_IPF�W�_* O�F``QF�AsD90�VHO_�� 5R42PSWq?�wTEL� P����90WORjAXQE� LVt�[R2�ICE���p�$cs  O����q��
���
�p�PS�A�w[# XK	�Iz0�AL��' �
���F����!�p��i��$� 2Q��P���������� Q���!�q�����$� _FLTR � �\� ��
��������$Q��2��7rSH`D +1Q� P㏙�f���ş��韬�� П1���=��f���N� ��r�ӯ�������ޯ �Q��u�8���\��� ����󿶿�ڿ;��� _�"�XϕτϹ�|��� ��������6�[�� �Bߣ�f��ߊ��߮� ��!���E��i�,�� P�b���������� /���(�e�T���L���l��z _LUA1�_x!1.��0���p���1��p�25c5.0��r��n���2����d %7I[3e��� ����[4���T'9[5U��� {���[6���@D �//)/s��Q�ȁMA��M?A�P����� Q� ��u.<�/?&?�/J?\? n?A?�?�?m�P�?�? �?�?�?O.O@OROOvO�O�Ou.kOl�q���O�L
ZDT ?StatusZO�O�5_G_Y_n�}iR�Connect:� irc{T//alert^�_�_�_ �_mW#_oo,o>oPo�bot�^�P~2g���go�o�o�o�o�o�o 	-?Qcul��$$c962b3�7a-1ac0-�eb2a-f1c�7-8c6eb5�6401a8  (�_�_���"�Rp�1!W��(��" S��JE�� X��C� ��,$���W���ˏ ���֏��%��I�0� m��f�����ǟ��������!��u�R������ DM_�!�����SMTP_CTRL 	����%����DF��� ۯt�ʯ��'��Lz�N�� 
j��y��q�u���������#L�USTOM' j������ � ���$TCPIPd�j��H�%�"��EL�����!���H!T�b<�n��rj3_tp�d7� ��i�!KCLG�L�i���5�!CRT�ϔ�����"u�!CON�S��M�[�ib_Osmon����