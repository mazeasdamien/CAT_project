��   �c�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����DCSS_C�PC_T 4 �$COMMEN�T $EN�ABLE  �$MODJGRP�_NUMKL\�  $UFR�M\] _VTX �M �   $�Y�Z1K $Z�2�STOP_T�YPKDSBIO�IDXKENBL_CALMD��USE_PRED�IC? �ELAY�_TIMJSPEED_CTRLKOVR_LIM? *p D� �L�0�UT�OOi��O���&S. ǰ 8J\TC �u
!���\�� jY0 � � �CHG�_SIZ�$A�P!�E�DIS"�]$!�C_+{#�s%O#J�p 	]$J d#� �&s"�"{#�)�$��'�_SEEX�PAN#N�iG�STAT/ D�FP_BASE_ $0K$4�!� .6_V7>H�73hJ- � q}�\AXS\3UP�LW�7����a7r � < w?�?�?��?�?�x//	7ELEM/ T �&B.2�NO�G]@%CNHA��DF#� $DAT�A)he0  �PJ�@ 2� 
&P5 �� 1U*n   �_VSiSZbRj0jR(��VyT(�R%S{TR/OBOT�X�SAR�o�U�V$CUR�_��RjSETU~4"	 $d �P_MGN�INP_ASSe#�P B!� `CiH�77`e��.fXc1�CONF�IG_CHK`E_�PO* }dSHRS�T�gM^#/eOTH�ERRBT�j_G]�R�dTv �ku�dVALD_7h�e�4hT1r
0R HLH8t� 0  lt<NerRFYhH~t�5"�1� ��W�_Ag$R��UPH/ (G%Q�Qt�Q3?wBOX/ 8�@F!�F!��G �r��s tUI}Ri@  ,��F�pER%@2 {$�p l��_Sf�uUIZ}N/ 0 IbF(@�p��Z_�0 _�0?wu0  �@�QWyv	*��~  ��$$CL`  ����!���Q���Q�VERSI�ON� � XK2�IRT�UAL�0�' 2� ?�Q  Q(�����&@^�
��ʐ����ϟ�(������d<�9�Cz  P�8���a� ��������ׯ��� ��.�@�R�d�f��� ���������Կ	�� *�<�N�`�r����ϫ� ��̿����߮�8� J�\�n�)ߒϧ߶��� �������%�4�F�X� ~�|ߎߣ�.������� ���!�0�B�T�f�x� �������������� />�P�b���v�� ��������+ :L^p���� ��� /'/9/H Zl/�/��/�� ��//#?5?D/V/h/ z/�/�?�/�?�/�/�? 
?O1OCOR?d?v?�? �O�?�O�?�?O	_�O -_?_NO`OrO�O�O�O �_�_�O�Oo_)o;o �_\_n_�_�_Mo�_�o �_�_�oo7IXo jo|o�o�o�o�R�o �o�3�E�Tfx �����Տ��ݏ ��A�S�b�t����� ����џ�����(� =�O�^�p��������� ʟ߯� ��$�9�K� ]�l�~���6���Ưۿ ����#�2�G�Y�h� z���������Կ���� 
��.�C�U�g�vψ� �ϬϮ��������<� -��Q�c�r߄ߖߨ� ����������)�8� M�_�������q� ���������4�&[ m|������������ v3BWix ������� />?/e/w/�� ���/��///(/ =?L/a?s?�/�/�/�/ �/�?�/O?$?9OH? ]OoO�O�?�?�?ZO�O �?�OO O2OG_VOk_ }_�O�O�O�O�O�_�O o_._CoR_goyo�o �_�_�_�_�o�_	o *o`oQ@u��o�o �o�o�o�o��&8 M�\q������� �����"�4��X� J��������ď������$DCSS_CSC 25���Q  P�;���Z���~� A�����w�د������  ��D�V��z�=��� a�¿��濩����߿ @��d�'ψ�KϬϾ� ���ϥ����*���N� �r߄�Gߨ�k��ߏ� �߳��&���J��n� 1��U��y��������GRP 2N� ����	� s�^������������� ��'��7]H� l������ �5 2kV�z ������/
/ //U/@/y/d/�/�/�/ �/�/�/	?�/-??*? c?N?�?r?�?�?�?�? �?�?OO'OMO8OqO \O�O�O�O�O�O�O_ �O%__"_[_F__�_ �_n_�_�_�_�_o�_�oEo0oio�_GS?TAT 2�E���< 6���`u�����<��#���?�`A=sǜ��=s�=.93��~{C���B� .C�����X`<�e?G��?� 47��R�84��s�?��`�`��`4��Z����e��l�Ͼ=�M�?t�C�>���ɾ��	�y�$�����D)�� y=�� �=�	�?}�`<� 5�`����vɿE������>=��P�c>�=%��?|ఀp���p��p�?���H�+�~Q�C|��CJ�+�D?Q y?H���?�׼#��G��p?�p=~��==t$�.9��?�a��AB�?c�D�� y�o �o�m��\�n��P� ������Џ����jp ������z!�O�5�G� i�k�}���͟��՟� �����ŏ{����� ��ï��������O� 5�c�-�k�Q�c����� �����Ͽ���� 9�g�i����ۯ���� �����'��/�]�� Eߓߥ�?����ߵ��� �����G�Y�3�}�� i�{���������� 1�C��/�y�o߁߯� ��[���������-? cuO���� ���)5_ 9K������w �/%/�I/[/5/c/ �/k/}/�/�/�/�/? �/?E??1?{?�?g? �?�?�?�?�?��?/O AO�?eOwOQOcO�O�O �O�O�O�O_+___ a_;_M_�_�_�_�_�_ �_�_oOOKo]o�_ io�omoo�o�o�o�o �oG!3}� i������� 1�C�9oG�y��e��� �������я��-�� �c�u�O��������� ៻�͟�)��M�_� 9�g���O�}�˯ݯw� �����I�#�5�� ��k���ǿ������׿ �3�E��i�{�U�g� �ϧ������ϓ��/� 	��e�w�Qߛ߭߇� ���߽����+��O� a�;�m��q������ ��������K�]�7� ����m����������� ��5G!O}W i������ 1��gy�� �����/-// Q/c/=/O/�/s/�/�/ �/�/??�/?M?C U�?�?/?�?�?�?�? OO�?7OIO#OUOO YOkO�O�O�O�O�O�O 	_3___i_{_q?_ �_K_�_�_�_�_o/o 	o7oeo?oQo�o�o�o �o�o�o�o�oO a;��q���_ ����9�K�%�7� ��[�m���ɏ����� ُ�5��!�k�}�W� ������������ 1�˟=�g�A�S����� ��ӯ寿������ Q�c�=�����s���Ͽ ��������M�� 9σϕ�oϹ��ϥ��� �����7�I�#�m�� Y߇ߵߏߡ������� !�3��;�i�#�Q�� ��K������������ 	�S�e�?�����u��� ��������=O );�{���g ���9K%o �[������ �#/5//A/k/E/W/ �/�/��/�/�/�/? 1??U?g?A?o?�?w? �?�?�?�?	OO�?#O QO+O=O�O�OsO�O�O �O�O_�/�O;_M_�O q_�_]_o_�_�_�_�_ o�_%o7oo#omoGo Yo�o�o�o�o�o�o�o !_)_Wiu� y������� )�S�-�?�����u��� я��ݏ���=�O� ES����q���͟�� ��ݟ�9��%�o� ��[����������ǯ�ٯ#�5��Y�k�a���$DCSS_JP�C 2`�Q ( DQ�����ʴԿذ���� ʿܿ1� ��$�y�H� ��l��ϐ��ϴ�	��� ��,�Q� �2߇�V�h� z��ߞ��������;� 
�_�.�@��d�v�� �������%���I�� m�<�N����������� ������3W&{ J�n����� ��AO4�X �|����/� �O//0/B/�/f/�/ �/�/�/?�/'?�/? ]?,?>?P?�?t?�?�? �?�?O�?5OOOXO }OLO^O�O�O�O�O�O �O_�OC__g_6_�_ Z_l_�_�_�_�_	o�_�o4c��S����L ouo&o�o�`ddo�o �o�o�o	�o-�oQ u<�`r�� ����;��_�&� ��J���n�ˏ��ُ�� �ڏ����m�4��� X���|�ٟ����ğ!� �E���0�y���f� ï��篮��ү/��� S��w�>���b����� ��������=��a� (υ�Lϩ�p��ϔ��� ������%�K��o�6� ��Z߷�~��ߢ����� #���1��k�2�D�V� h����������1� ��U��y�@���d�v� ����������? c*�N�r�� ����q 8�\����/��%/�FdMODE�L 2Skx\�o(
 <o$c (_  o&�( �/�/�/�/�/�/�/�/ ??d?;?M?�?q?�? �?�?�?�?O�?ONO %O7OIO[OmOO�_�O y/�O�O&_�O_\_3_ E_W_�_{_�_�_�_�_ o�_�_oXo/oAo�o eowo�o�o�o�o�o �o�O�O�O/� �������� P�'�9�K�]�o���Ώ �����ۏ����#� 5���Y�k���Se�� ���������1�C� ��g�y�Ư������ӯ ���D��-�z�Q�c� u���������Ͽ�.� ɟ۟	�ψ��qσ� �ϧϹ������<�� %�7߄�[�mߺߑߣ� ��������8��!�n� E�W��?�Q�cϑ�� y�����F��/�|�S� e�w������������� 0+=Oa� ��������> ���]o�� ������/#/ p/G/Y/�/}/�/�/�/ �/�/$?�/?Z?1?C? U?+�?O}?�?�?�? �?2O	OOhO?OQOcO �O�O�O�O�O�O_�O __d_;_M_�_q_�_ �_�_�_�_�?*o�?�_ oroIo[o�oo�o�o �o�o�o&�o\3 EWi{���� �����/�A�o ��;oi�{�菿�я� ����+�=�O���s� ��ҟ����͟ߟ�� P�'�9���]�o����� ���������߯�^� 5�G���k�}���ܿ�� ſ����H��1�C� ��g�y��ϝϯ����� ����D��-���'� U�g���O߽������� �R�)�;��_�q�� ���������<�� %�7�I�[�m������� ���ߝ�����J��3 EWi{���� ���/|S e������� 0///f/A/S/ �/;/�/�/?�/�/>? ?'?t?K?]?o?�?�? �?�?�?�?(O�?O#O pOGOYO�O}O�O�Ow/ �/�/�O�O�O_1_~_ U_g_�_�_�_�_�_�_ �_2o	ooho?oQoco uo�o�o�o�o�o�o �Ov_?Q' �����*��� %�7�I�[������ޏ ��Ǐُ����\�3��E���i�{���Җ�$�DCSS_PST�AT �����Q  �  �� � (&�K�2�o���� ������$�˟į֯���� ����'��SETU�P 	�B�����X�r����������ۿ�g��T?1SC 2
K����Cz�#�5�G; �CP R�D$�Dl�Ϥ�^�� ���ϻ��"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t����� ����������( :L^p���� ~������-� Qcu����� ��//)/;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?m?? �?�?�?�?�?�?�?O !O3OEOWOiO{O�O�O �O�O�O�O�__/_ BS_e_w_F_�_�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o �������� �#�5�G�Y�k�}��� ����ŏ׏����� 1� _U�g�y��_���� �������	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{�J��� ��ğ���������/� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������� #5GYk}� ��������/ 1/C//g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_� !o3oEoX/io{o�o\o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟��� �#�5�G�ok�}��o ^���ů������� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹������� ��%�7�I�[�m������$DCSS_�TCPMAP  ������Q @ �������������������	���
����������W�  ���������*������⡋�U��������U���� ��!��U"��#��$��%��U&��'��(��)��U*��+��,��-��U.��/��0��1��U2��3��4��5��U6��7��8��9��U:��;��<��=���>��?��@��UI�RO 2����������� 0BTfx��� ����,1��U��y��� ����	//-/?/ Q/c/u/�/�/�/6�/ Z�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7O�/[O�/O �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_�_�_NO�_��UIZ�N 2��	 �����(o:oLoR�%o zo�o�oao�o�o�o�o 
.�oRdvE �������� *�<�N�`�#�����e� ��̏ޏ�����&�8� �\�n���C�����ȟ ������ӟ4�F�X� '�|�����c�u�֯������0��_��UF�RM R��� ����w���������ѿ �����+�=�O�a� sυϗϩϻ������π��'�9�K�\�r��\߄ߖ�qߺ��ߧ� �����&�8��\�n� I����������� ���4�F�]�o�|��� -������������� 0TfA��w �����> Pg�t�%��� ���/(//L/^/ 9/o/�/�/�/�/�/�/  ??�/6?H?_l?~? ?�?�?�?�?�?�?�?  O2OOVOhOCO�O�O yO�O�O�O�O
_�O._ @_W?d_v__�_�_�_ �_�_�_�_o*ooNo `o;o�o�oqo�o�o�o �o�o&8O_!n ������� �"��F�X�3�|��� i���ď�����Տ� 0�B�Yf�x������ ��ҟ䟿�����>� P�+�t���a�����ί ����߯(�:�@�