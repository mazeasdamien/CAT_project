��  
�,�A��*SYST�EM*��V9.4�0107 7/�23/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����ADV_I�N� 0   � O�PEN� CRO �%$CLOS�� $�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�o#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO>""ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� _"��!_I�F� � $_ENABL@t#T� P dt#UE5K%1CMA�s �"�
� �OG�f J0CUR�R_u1P $�3LI�N@�1z4$t$AU�SOK4� OD2$�SEV_AND_�NOA 3PPIN�FOEQ/  ��L �0p1�5�1� H �749E�QUIP 3n@NAM0�,B�_OVR�$V�ERSI� �!P�COUPLE]  o	 $�!PP�1�CES0�2eG  �"P�0�2
 �� $SOFT��T_ID�2TO�TAL_EQ 0Ă1�@N" �@U SP�I
 �0^�EX�3C�RE -DdBSI�GJ@dOvK�@P�K_FI90	�$THKY"WPA�NE�D � DU/MMY1dIT1�TU4QQ���AR�x1R� � /$TIT91� �� � �Td�T0�ThP�TU5�V6�V7�V8�V9�W0�W�WOQ�U�W�gQ�U�W1�W1�W1��W1�W2�R�SBoN_CF�!@$<!J� ; ;2�1�_CMNT�$�FLAGS]�C�HEK"$�b_O�PTJB � ELL�SETUP � `@HO8@9 P�R�1%�c#�aREPR�hu0D+�@���b{uHM9 MN�B;16 UTOB�J U�0 }49DEVIC�STI/@�� �@b3�4pB�d�"VAL��#ISP_UNI�tp_DOcv7�yFR_F�@|%u13���A0s�C_WAx�t,q�zOFF_T@]N�DEL�Lw0pdq�1�Vr?^q��#S?�o`Q"U��t#*�QTB��bMyO� �E � �[M�����RE�V�BIL���!X�I� v�R  �!D�`��$NOc`M�|����ɂ/#ǆ� �ԅ��ނ�@Ded �p E RD_E���h�$FSSB�6�`KBD_SEV�uAG� G�2Q"!_��2b�� V!�k5�p`(��C�00q_ED|� � � t2d�$!S�p-D%$� ��#�B�ʀ_�OK1��0] P_C�� ʑ0t��U �`LACI�!�a�Y�� ��qCOMM� # $D
� ��@���J_�\R BIGALL;OW� (Ku2:-B�@VAR���!|�AB   �BL�@� � ,K�q��r�`S�p�@M_O]�˥��CCFS'_UT��0 "�A�Cp'��+pXG��b�0� 4� IMCM ��#S�p�9���i �_�"t\b���M�1 h$�IMPEE_F�s���s��� t����D_(�����D��F��� �_����0 aT@L��L�DI�xs@G�� �P�$I�'�����CFed XF@GRU@��Mb��NFLI�\Ì@U�IRE�i42� SgWITn$`0_N�`�S 2CF�0M�' �#u�D��!���v`����`J�tV��[ E��.p�`��>�ELBOF� � շ�p`0���3����� F�2T��A`��rq1J1��z _To!��p��g����G� �r0WARNM�p#tC�v`�ø�` � COR-�UrFLTR��TR�AT9 T%p� $ACCVq��� ��r$ORI�_&��RT��S<��HG*�0I���TW��A��I'�T���H9K�� �2028�a1��HDR�2��2�2J; S���3���4��5��6��7
��8��9��׀
 �2� @� TRQB�$vf��'�1�<�c_U<�G� COec  <� P�b�t�x53>B_�LLEC��}!~�MULTI�4��"u�Q;2�CHI�LD��;1ذO�@T�� "'�STY 92	r��=��)2��������ec# |@r056$J ђ��`����uTO���E^	EXTt����2��22"����$`@D	�`&��p������(p�"��`% �ak�����s�����A&'�E�Au��Mw��9 �% ��TR>�� ' L@�U#9 ���At�$J�OB����P��}IG��( dp��� ���^'#j�~�L��pOR�) tf$�FL�
RNG%Q@�TBAΰ �v&r� *`1t(��0 �x!�0«+P�p�%4��*��͐U��q�!�;2MJ�_R��>�C<QJ�8&<J D`5CF9���x"�@J���P_p�7p+ \�@RO"pF�0��I9T�s�0NOM��>Ҡ�4s�2�� @U<PPTgў�P8,|Pn�ć0�P�9�͗ RA����l�?C�� �
$�TͰtMD3�0TD��pU�`�΀+AYHlr>�T1�JE�1 \�J���PQ��\Q��hQ�CYNT�P��PD'BGD̰�0-���PU6$$Po�|�u��AX����TAI�sBUF,�O!�A�1�. ����F�`PIV|�-@PvWMuX�M�Y�@�VFvWSI�MQSTO�q$7KEE�SPA��  @?B�B>C�B�2��/�`=��MARG�u2��FACq�>�SLEW*1!0����
�4ذs�CW$0'����pJB�Ї�qDE�Cj�e��s�V%w1 Ħ�CHNR�;MPs�$G_@�g�D�_�@s��1_FP�5�@TC�fFӓC@�Й���qC��+�VK��*��"*�JRx���SoEGFR$`IOh!v�0STN�LIN>�csPVZ�z�Ц@�D2����r 2��hr�r��1��3` + ^?���եq�`��q|`������t��|aSI!Z#�!� �T�_@%�I��qRS�*s���2y{�Ip{�pTpLpF�@�`��CRC����CCTѲ�Ipڈ�a8���bL�MIN��aP1순���D<iC �C/���!uc�OP4�n �j�EVj���F��_
!uF��N����|a�֔=h?KNLA�C=2�AVSCA�@�A�WQ�a�4�  cSF�$�;�Ir�Kঠ'��05��	 D-Oo%g��,,m�����ޟ��RC�6� n���sυ��U��R�0HANC���$LG��ɑDQ�$t�NDɖ��AR۰N��aqg��ѫ�X��ME��^�Y�[PS�RAg�X�AZ�П���:rEOB�FCT��A���`�2t!Sh`0ADI��O��y�s"y�n!@�������~#C�G3�t!��BMPmt@�Y8�3�afAES$���v��W_;�BAS#?XYZWPR��*��m!��	y�U�87/  ƀI@d��2�8\�p_C:T����#��_L
 � 9K ���C�/�(z�J�LB�$�3�xD��5�FORC��b�_AV;�MOM$*�q�SaԫBP`Ր� y�HBP�ɀE�F�����AYLOAD&$�ER�t&3�2�X�rp�!ҁ�QR_FD��� : T`IH�Y3��E�&��Ct���MS�PU
$0(kpD��9 �b��;�B�	EVId�y
�!_IDXY�$���B@X�X�<&�SY5� � �HOPe�<��AL�ARM��2W�r}rR9_�0= hb P�nq�`M\qJ@$PiL`A&�M#�$�` ��� 8�	���V�]�0�U�qU�PM{�U���>�TITu�b
%�![q�BZ_;�.��? �B pQk���6NO_HEADE^az��}ѯ��`� �����dF�ق�tc`����@�@��uCIGRTR�`��ڈL���D�CB@4�RJ�� 1�[Q���A�2>�&��OR�r��O����T`UN_OO�Ҁ�$����T������I�VaCnp�DBP�XWOY���B��$SKADR��DB]T�TRL��C���րfpbDs��~�DIJj4 _�DQ}���PL�qwbWA���WcD�A��A�=�2�UMMY�9��10�VIȾ ����D;[QPR�� 
M�Z���gE O�Y1$�a{$8��L)�F!/��
����0G�G/��9�PC�1H�f/3#PENEA@T�f�I�/���RE�COR`"JH y@ �E$L�#F$#PR���+jp���nq�_D$�qPROSS]�
���R�r�` >u�$TRIG96�PAUS73ltETgURN72�MR:�eU 0Ł0EW$�~�SIGNALA��QR$LA�З5�1�G$PD�H$PDİ�AI�0�A�C�4�C��DO�D�2�!��6GO_AWA�Y2MOZq�Z��,CS��CSCB�g�K Իa#���E+RI�0Nn�T�`$�����FCBPL�@QBGAGE���P��ED`|BD�wA[CD�OF�q�[F0�FoC��MPM�AB0XoC�$FRCIN��2Dk��@��O$NE�@�FD�L8�� L� �����=��Rw�_��P>� OVR10����lҠ�$ESC_|�`uDSBIO��p��pTe�E�VIB�� `s��Z��V��p�SSW��$�VLY�:�Lk��X���ѣ�0bQ����USC�P��qA=�	Q��MP1%e@&S*`�(bt`'c5۳ESUd��-cWg&S Wg?cWd����Wd��Wd<.���AUTO$�Ya҃�ac�SB����-d���&SwB[��GB�f_$VOLT�g ���  �GAOD!��q���@:�ORQ�ҀKra�$DH_THE&0�Rgp� <qtnwALPHnt��o��w0 Vp]�$�.�Ra�[��s�5�`r�CQ�#BUD�S� F1M���sV
��;��L�b�tk���BRTHR��L��T`�Z���Vɖ��D)E  �1��2�⋅ ��������kѯ�a� �Tt0V�ꆸ������@̈Я�-�"�N~���sS2����INHB��ILTG0ɡ�T?� �3$�w��E��PqQxQ��TqPe��0Y�AF}�O�ນ��ڗ ��qPڳē����bPܙ���PL?���3���TMOU��ēS��� � ��s�/�S18���O��Aܙ��I����CDqIƑ˩o�STI��գ�O:ҋ�,0���AN��Qg�S��+r�#x$�����w�1_����PRA�P`�vC����MCN�eQe�����VER�S��r�oPIw�F�PåǲШ۷G.�DEN��G>�����F�2H�Ƿ�M�7�F��_�MN�D̠,���@�d�{ƭa����OB����U˱z���DI ���#���3�����A��w�Fx���3�O�N�5��Q��VAL��CR[�_SIZp��b�;Qn�REQ�R�b��]2b���CH q�΂�ڃ�Ռ�����:�n�S_U��X��wW�FLG���wU$CV�iMGP�QδFLXP�923R�u�L��EAL�P-�C	�F+rT��W��� �R��c���NDMS�7� ��K>S�P_M'0h�STWv������AL�P���Q����U���U�IAG@,�o��d�U�-�T"	A-`� ���A��� ��H`��Q`��6��Pq_D&��1s��.�P��F�"2�T�� ?7 1A>���#�#L��?`_=i @@>LD�pc�F�0�FRI�0 `Ѐ��1}Ѳ�IV\1�*�^1�U�P`��a��C�L!W��
`L=S&-c&&S�C.w��  L���!����d�Q$w!�҇��$w��p��
�P�5RSM��P���V0h � r�l�d^2AW�a_TRp�}�8@NS_PE�A����< ��$�SAVG�8�6G]%���CAR �`�!�$���"CRa���$ d�#qE�@��"STD���!Fpo��'QOF0��%��"RC���&RC۠�(F�2A�R#7����%, gMA�Q_�a��
QQ��al2��%u4Ib�r7I�R�9�wQ�7�8M/��!C:pR�  �p�2F<�SDN�a0 � W2QM P $Mi��s$cA �$C�cm�9���4���AT�0CY_ �N LS!IG1@x'yB��y@@H2Y��NO����SDE�VI�@ O@�$�RBT:VSP0�3�CuT�DBY|�A�	W`3CHNDGD�AP H@GRP�HE iXL�U��VSЌFx2� DL1p aQ6ROp��FB�\]�FEN�@��S���ChAR d�@DyOd�PMCSb���P薇P�R��HOT�SWz42�DMpEL�E�1/ex\8`�RS T�@���r� hf��`OL�GHA�Fk�Fs�����C�A@�T � $MD�LUb 2S@�E ���q�6�q	0�i�c�e
�cJ��	uݢ�#~X5t+w�PTO��� x�byU DSLAVS�� U  ��INAP �	V�ЊyA_;�wENUAV $R��PC_�q�2 1bLp�wpp B�pSHO+� W ���A�a�qB�2�r�v�u�v�b�_CF� X�` ,f��r�OG� gE��%D�h��p2C�Iߣi�MA��D��x AY?�W� p�N3TV	�D�VE�0@�SKI��T�`g?Ň2�� JZs�! �Cꆻ��f�_SV</ �`XCLU��H����ONL��'�Y��T��OT:eHI_�V,11 APPLY���HI4`;�U�_M�L�� $VR�FY8�	�U�M{IGOC_I���J 1/d��߃O�@X�LSw"�`@$DUMMY�4���ڑ�Cd L_TP���kC��^1CNFf���E��@HT�y� D_#UQ_��ݥ�YPCP��=�� ������uJ �ҟ Y +�
0R�T_;P��uNO�CCb Z�r�TAE���=�פ�DG��@[ D�P_B�Ae`kc�!I��_��H�t~T��E \�pyAb=cARGI�!�$���`[��SGNA] ��`U���IGN�Տ��� ���V������ANNUN��&�˳�EU�<J'�ATCH���J��B��u^ <`@g�����:c$Va������ᑴaE�F] I�� _ �@@FͲITb�	$TOTi �C�O��c� @EM�@NIF�a`tB��c��ùA>���DAY@CLOAD�D\�n���� �EF7�X�I�Ra��K���O�%��a�ADJ_)R�!@b��>�H2��"[�
 c�%��`a�͠MPI�J��D��qA��?�Ac 0� �х�� ��Z�ϡ��Ui ��CTRLܖ Yp d��TR�A8 ?3IDLE_�PW  �Ѡ��Q��V��GV_���`c ��o�;Q@e� �1$��6`<cTAC�-3��P�LQ�Z�Rdz\ A-u:ɰSW;�A\���/Jղ�`b�K�OH�(OsPP; �#IRO� ��"BRK��#AB  �������� _ ���F���`d͠, j@�S�RQDW��MS��P6X�'z��IF�ECAL�� 10^tN��V��豊�V�(0}f�CP
��Nr� Yb�0FLA_#f�OVL ��HE��>�"SUPPO��ޑ�\�L�p��&2XT�$Y-
Z-
W-
���/��0GR�XZl�q�$Y2�CO�PJ�SA�X2R��*r�!���:��"�rI�0)��f `�@CACH�E��c��0�s0L}AZ SUFFI, C��q\��哹6��QMSW�g� 8�KEYIM[AG#TM�@S���n
2j�r���ROC�VIE��~�h ��aBGL����`�?G� 	Q���i��m!`STπ!� �����n����/EMAI�`N��`A��`Z�FAU� �jH�"�qa��U�3�qq� }�k< �$I#�US�� �IT'�BUF`�r�DNB���SUBu$��DC_���J"��"SAV�%�"k�������';��P�$�UOR	D��UP_u �%��8OTT��_B`��8@�LMl�F4��C7AX�@Cv���Xu 	��#_uG��
 @YN_��R�l6���D�E��UM����T��F���caC�DI`BED%T)@C��~�m�rI��G�!c�&��l`���-�P��FZP n (�pSV� )d\��ρ���2ΰ��o�� ����>"$3C_R�IK��kB���hD{pRfgE.(AD�SP~KBP�`�II�M�#�C�Aa�A��UЂG���iCM! IP`��KC��� �DTH� ȷS�B*�T��CHS�3�CBSC��� ���V�dYVSP�#[T_D^rcCONV�Grc�[T� �Fu F�ቐd0�C�0j1��SC5�e�]CMER;dAFBgCMP;c@ETBc� p\FU D�Ui ��+�~�CAD�I%P702#@O��B�qWӏ�SQ��QǀSU��MSS�1ju�4`��TB�Aa��A�1r�� "�Й��4�$ZO@s���l�U�6�&��eP���eCN�c�l��l�l�iGRO�U�W)��S c�MN�kNu�eNu�eNpR|b|�i�cH�pi��z
 �0CYC���s�w�c���zDEL�_D��RO�a���qVf���v{�O�2���1���t��:R�ua�.#�� ���AL� �1s@ˢI1¡�J0�PB��,렒�ER^�T�Gbt ,!@��5��aGzI1LcR1s 
�0&ԠNO��1u����H�����P����Cڠ	�����!���J0��0vH *	�L U�1#J�Q��V
�[�7A z���z��z�n�z�Ѩz�Fz�7w�8w�9Pw���y���1��1��U1��1��1Ě1њU1ޚ1�2��2�����2��2��2��2�Ě2њ2ޚ2�3J��3��3����3��U3��3Ě3њ3ޚ�3�4���EXTF��1w6�.(�0�f�0��U�0ŷ�e.�FD�R5�xTU V�E��?1���SR��R�E�F���OVM�~C)�A2�TROVf2�DT� R�MXa��IN2���Q�2�IN	Dp�r�
���0�0�0�Gu1��[�G`��{�D_�[�RIV�P��oGEAR~AIOr�	K"N�0�y�p��5`@�a�Z_MC�M� ���F��U�R�Ryǀ��!?3 ��p?nЋ�?n�ER�v�Gme��!�P��zIj:�PXqB�RI0%�>`�#ETUP2_� { ���#TDPR�%TBp�������K�"BAC�2| QT��"�4)�:%	`t^B��p�IFI���� Mc���.�PT|��I �FLUI��} � ��K UR�c!���B�1SPx NE�EMP�p�2$��]S^�?x��Jق�0
3VRT���0x/$SHO��Lq�6 ASScP=1��PӴBG_�������FORC�3" �i�d~)"F%UY�1�2\�2
A�h� p� |��N�AV�a��������S!"��$VI�SI��#�SCM4S�E����:0E�V�O���$���M����$��I��@��FMR2��� �5`�r�@ �� �2�I�9 F�"��_���LIMI�T_1�dC_LM�������DGCLFl����DY�LD����5������F  ���D u	 T�sFS0Ed� P���QC�0$EX_QhQ1i0�P�aQ53�5��GoQ��g� ����RSW�%�ON�PX�EBUG���'�GRBp�@U��SBK)qO1L� ��POY 
)�(�P��M��OXta`KSM��E�"�0�����`_E � x
@F���TERMZ%9�c%�aORI�1_ Y�c%d�SMepO��B_ �|&.�`�(�c%��e:�UP>� ?�� -���b����q#� ���G<�*� ELTO��p�0�PFIrc�1Y���P�$�$�$UFR�$��1L0e&� OTY7�PT4q��k3NST�pPATz�q4PTHJ�a�`EG`*C�p1AR�T� !5� y2$2R�EL�:)ASHFTPR1�1�8_��R�P�c�& � $�'@�@� ��s�1 @I�0�U�R G�PAY�LO�@�qDYN_�k���.b�1|��'PERV��RA��H��g7��p�2�J�E-�J�R�C���ASYMFgLTR�1WJ*7����E�ӱ1�I��aUT�pbA�5�F�5aP�PlC�Q1FOR�p�M��GRI!����W��/&�0F0�a H��Ed� �m2N���5`OC1!?�$OP����c��c���bRE�P�R.3�1a�F��3e���R�5e�X�1(�e$PWR��_���@�R_�S�4��et$3U�D��.�Q72 ����$H'�!�`AWDDR�fHL!G�2(�a�a�aT��R��U�w� H��SSC����e-��e���e��S�EE��HSCD���� $���P_"�_ B!rP����}T!HTTP_���HU�� (�OB�J��b(�$�fL�Ex3pWq�� �� ���ะ_��T�?#�rS�P��z�KRN�LgHIT܇5��P ���P�r������PL���PSS<�ҴJQUERY_FLA 1��qB_WEBSOC���HW�1U����`6PINCP	U���Oh��q�����d���d���� �I�HMI_ED� T� �RH�?$��FAV� d�Ł��wOLN
� 8��yR�@$SLiR�$INPUT_�($
`��P�� �؁SLA� ����5�1��C���B��IO6pF_AuS7��$L%�}w%�A��\b.1��0���T@HYķ������Qh�UOP4� `y�ґ�f�¤�������`PCC
`���#���aIP_M�E�񵁗 Xy�I�P�`�U�_NET�9���Rĳs�)��DSP(�Op=��BG�����M��A��� lp:CTiAjB�pAF TI�`-U��Y ޥ�0PSݦBUY IDI�rF ���P�q�� �y0��,����Ҥ�N�Q�Y R��IRCA|�i� � ěym0�CY�`EA������񘼀�CC����R�0�A�7QDAY_<���NTVA�����$��5 ���SCA�d@��CL���� ���𵁛8�Y��2,e�o�N_�PCP�q��ⱶ��,�N�����
�xr���:p�N� �2��Ы�(ᵁ�p���xr۠LABy1���Y ��UNIR��Ë ITY듭��e�ւR#�5���R�_URL���$AL0 EN��ҭ� �;�T��T_U��A�BKY_z��2DI�SԐ�kSJg�����P�$���E��g�R���З A�/���J����FLs��7 Ȁ|���
�UJR� ���F{0G��E7��J7 O^ R$J8I�7�H�R�d�7��E�8{��H�APHIQ�S��DeJ7J8�B��L_KE*� � �K��LM�[� � <X�X�Rl�u���WATCH_VA��o@D�tvOFIELc��cy��L��4� � o1Vx@��-�CT[�9�m�� ��LGH���� $��LG_SIZ�t�z�2y�p�y�FD��Ix���+!�� w�\ ����v��S��� 2��p�������\ ��h�A�0_gCM]3NzU
RFQ\v�v�d(u�"B ��2�p����I��+ �\ ��fv�RS���0  ��ZIPDUƣp�L)N=��ސ�p��z6���f�>sD�PL�MCDAUiEA`Fp���TuGH�R�.OGBOO�a��� C��I�IaT+���`��RE����SCR� �s��D�I��SF0�`RGIO"$D�����T("$�t|�S�s{�W$|��X��JGM^'MN3CH;�|�FN��a&1K�'uЅ)UF�(1@n�(FWD�(HL�)STP�*V�(%Г(,��(RS9HIP�+��C[T�# R��&p:'^9U=q�$9'�H%C�d���"Gw)�0PO�7��*��#W}$���)E]X��TUI�%I�� �Ï���rCO#C� N*�$S��	)���B@�NOFAN1A|��Q
�AI|�t:��EDCS��c�CT�c�BO�HO�GS����B�HS�H(IGN������!O���DDEV<7LL�ѩ�|��­Ц(�;�T��$��2�p������#A
���(�`�{�Y���POS1�U2�U3��Q	��2�@�Ш ��{�PtD�����&q)��0�d��VST�ӐR�Y��B@ ` _�$E.fC.k��p<p=fPf���4�ѩ LRТ� ��x�c �p��<�Fp�d��?"�/_ �����Kqx&���c �MC7�� ���CLD�PӐ��TRQLI0#ѽ�ytFL��,r��5s8�D�5wS�LqD5ut5uORG���91HrCRESERAV���t���t���c~�� � 	u095t5u��PTp���	xq�t�vRCLMC�������q�q�M��k�������$DEBUGMA�S��ް��?U8$T�@��Ee�g���MF�RQՔ� � �j�HRS_RU�7��a��A��k5FgREQ� �$/@x�OVER��n�t�V#�P�!EFI�%�a��g��d���tǯ \R�ԁd�$9U�P��?A��SPS�P��	߃C���͢a��U\�l��?( 	�MI;SC� d@�QkRQ��	��TB �� Ȗ0A՘AX����ؗ�EXCE�SjҔЪ�M��\���W����ԝ���SC>�P � H��̔�_��Ƙǰ]���
�MKHԳK�J� �m�B_K�FLIC��dB�QUIREG3MO��O˫3���ML�`MGմ @�`��T���a#NDU�]��>���k�G�Df��INAsUT���RSM>�a��@N�r]3-��p�5�PSTL\�� �4X�LOC�VRI�%��UEXɶANG�uBu�R�ODA��ŷ�������MF O����Y�b@�e4Ŝ2k�SUP�e��F�X��IGG� � �A��c���c Q6�dD�%�b|�!`�Ȁ!`��|��3w�ZWa�T!I��p�a M��[��� t��MD��I��)֟@���H8ݰM��DIA��ӂ��W,!�wQ�1�D��)��O���]��[ 0�CU��VPА�p���!_V��ѻ� ��P�S�X�5�	�����P��0N��ЍP��KES2���-�$B� ����ND2x����2_TX�d�XTRA�C?�/��qM�|q�`�Pv�`�XҰ�Pt SBq`^�USWCS��T��<	���PULS��A��NSޔ��R��JOIN��H��~`j�=��b��b�����P�=��$��b$���TA����S���S�HS�ME��SCF�aPJ���R��PLQ� 
M��LO��н.�L��^����8��Ҹ����0�RR2���O 1��eA�q/ d$��Iΐ+��G�A2+/� ;�PRIN�w<$R SW0"��a/�ABC�D_�J%�¡u��_J3:�
�1SPܠe�u�P��3��р`
u��J/���r�q�O8QIF��CSKAP"z{�{�J���QL2LBҰ�_AZ�r�~ELxQ��OCMP���T���RT�����c1�+���P1��t>@�Z�SMG0���=�JG�`SCL<�͵SPH_�@���%V�u� RT�ER`  �< A_�@G1"�A�@c���\$DI�
"23U�DF�}!LWn�(VELqIN�b)@� _BL�@u��$ G�q�$�'�'�%`<��� ECHZR/�TS�A_`����E�}`<����5�Bu�Ht1}`_�� �)5 D2d%��A4I��N9t&FR�DH�A���ÀP�$V `�#>Aa$��Ͳ�$Q���R}ӆ��H? �$BELvᵆ><!_ACCE�!c�x�7/��0IRC_] ���pNTT��S'$PS�rL�d� /Es��F{�@F
��9gGCgG36B���_�Q�2�@�A���17_MGăDD�A]"ͲFW�`���3�EC��2�HDE�KPPA�BN>G��SPEE �B�Q%_pB�QY�Y�|�11$USE_��,`Pk�CTReTYhP�0�q P�YN��AAe�V)хQM����ѷ��@O� YA�TINCo�ڱ�B�DՒ�WG֑ENC����u��.A�2Ӕ+@INPO�Q�I6Be��$NT|�#�%NT23_�"ͲIcLO� Ͳ_`��I�_�if� _�k�? ȼ` ej�C400fMOSI�A���ОA䃔�PERCH  �c��B" �g��c��lb =�����oUu@�@		A6B(uLeT	~��1eT�ljgv�fTRK@%�AY��"sY��q 6B�u�s۰�]��RU��MOMq�ՒY�MP�^��C�s�CJR���DUF �BS_BCKLSH_C6B )����f���St�H��R�R��QDCLALM�-d���pm0��CHK����GLRTY ���d��Y��)Üd'_UM]�ԉC��A�!�=PLMT� _AL�0��9��E� .� ��#E)�#H� =�0�Q3po�xPC�ax�HW�頿EׅCMC�E��@�GCN_,N�D�Ζ�SF�1�iV oR��g<!��0r���7CATގSH)�, �DfY��f��7A����܀PAބ�R_P݅�s_ �v��X�s����JG�T]��Y�����TORQ�UaP��c�yPOU`��b��P%�_W�u �t��1D��3C��3C�UIK�IY�I�3F�`6�����@VC�00RQ�t��1���@ӿ��ȳJRK������UpDB M��UpM�C� DL�1BrGR�VJ�Cĭ3Cĳ3$�H�_��"�j@q�COS~˱~�LN���µ �ĭ0�����u�����ē��Z���f$�MY���؊���>�TH�ET0reNK23��3hҧ3��CBm�C5B�3C! AS� ��`u��ѭ3��m�SB�3���x�GTS$=QC������������$DU��Kw�B�%(��%Qq_��a��x�{�K���b(��\сA`Չ��p�{�{�LCPH~�g�Aeg�Sµ ��������g������֚�V��V��0��UV��V��V��V��UV	�V�V%�H��@������G�����H��UH��H	�H�H%��O��O��OV	��O���O��O��O��O*	�O�O�Fg����	�����SPBA?LANCE_-��LE��H_`�SP�!1��A��A��PFULCElTl���.:1��UTO_<����T1T2��22N���29`�!�q�nL�=B�3�qTXpO�v 
A4�INSEG�2�aREV��`agDIF�uS91�8'6t"1�`OB.!t��M��w2�9`��,�L�CHWARRCBA	B�� ��#�`-ФQ 5�X�qPR��&���2�� 
�""��1neROB͠CR0r|5�����C�1�_��T � x� $WEIGH��P`$��?3àI̡Qg`IFYQ�@LA�G�Rq�S�R �RBILx5OD�p�`V2ST�0V2P!t�W0P�11�&1/0�30
�Px�2�QA  2řd^[6DEBUg3L_@z�2�MMY9&E� Nz�D`$D�_A�a$�0��O� � �DO_:@A.1� <B0�6��m�Q�B�2�0N�-cdH_p`�P��2O��� �� %"��T`"a��T/!�4�)@TICKh3| TE11@%�C ��@N͠�XC͠R?��Q�"�E��"�E8@PROMP��SE~� $I�R��Q��R;pZRMCAI)��Q�R4U_r0C2S; �q�PR8�7COD�3FU�Pd6ID_[�vU R!�G_SUFFu� �l3�Q;Q�BD�O�G �E�0�FGR r3�"�T�C�T�"�U�"��Uׁ�T8D�0�B0Hnb _FI�19*c7ORD�1 50�2�36V�+b�Q1@$�ZDT}U 1�0;E��4 *:!L_N�AmA�@�b�EDEF_I�h�b�F�d�E�2��F�4�F�c�E�e�FISP��PAKp�Ds�C�d��44בi��2�D�"�It�3D�O|#OBLOCKEz���S�O�O�Gq�R�PUM�U�b�T�c�T�e�T !r�R�s�U�c�T�d�R �6�q�S� ���U�b��U�c�S�Z��X�@P@` t�@qe�)@W�x4���s 1TE�<D��( l1LO�MB_��ɇ0V2V�IS;�ITYV2A���O�3A_FRI��a SIq�Q!R�@��@�3�3V2�W��W�4����_e��QEAS^3�Rϡ���_�[p:R�4�5��6_3ORMUL�A_Iz���TH]R^2 �Gtg�30�f��<8�5COEFF_O�A	 ��A���GR�^3Sg0BCAnO/C$��]30�1�GRP� � �G $�p�YBX�@TM~w���u�B�s��bCER, Tttsd$`7�  �LL�TSpS~�_SVNt�ߐĸ�$`�@��$`� ���SETUsMEA*P�P��W0�1+b>/0� � h��  @ڐo�l�o�cqDz��b�@cqq`t�P�G��R�� Q\p�*q[p��>�c NPR�EC>at��ASKy_$|�� PB1?1_USER�e"��{ ���VEL@���{ 0�$Ō!I]`���MT�ACFG>���  �@@ =O�"NORE-0l@,o�V�SI.1�d��6��"UXK�fP!��D�E�� $KE�Y_�3�$J3OG��0SV���0���!��}�SW�"�ah\aS�ՐT|�GI����| ^�� 4 �h��'d2�!XYZ�c���31�_ERR#�� 8Ԡ�A�fPV�d��1����/$BUF��X�����MOR|�� HB0CUd�lA�!��GQ�\aB�,"!a$� ���a��u��?��G~�� � $cSIՐ���VO��<T�0OBJE_���ADJU)B��EL�AY���%�DR�O�U.`=ղВQ0b=��T���0���;BDIR���; I�"�0DYNW�2��T���"R���@�0�"��OPWORK����,%@SYSBUy�SOP��ޑ�U�; P�pN�<��PA�t�>�"��OP�PUd!0�`!�Ľl�IMAGw��B0y�2IM�Õ�I�Ne�d��RGOVCRD��-��o�Pq����0��J�Os���"L�pBa���o�PMC�_Ee`���1Ny M� A�21�2T���S�L_��� � $OVSL�ǫ�?qD�`��2�" -�_�� k�P��k�Pu���2�C� �`�Ź�^��_ZER�D��$G�� 82=���� @*����%Oh`RI��� 
 JP8+��=!/��L��ح�T� �0A�TUS��TRC_T���sB��}f�s�9s�1Re`��� !DFAm����L���"`��0a� ޱ��XEw {�����C0�vUP��+p	qPX�P�j�43 � ��PG\���$SUBe�%�qe9JMPWAIT ,z}%LO��F�A�RCVFBQ�@x"�!qR�� �x"ACC� �R&�B�'IGNR�_PL9DBTB2�0Pqy!BWbP�$2w�Uy@�%IGT�P=I��TNLN�&2�R��rL�NP��P�EED \HADCOW�06�w��E[pq4jO!�`SPDV!� LbAz�`�07�3UNIr��02"!R��LYZ`� �o/PH_PK���e�RETRIE9{�q���0'P;FI"�� �G`�0�D 2�g�DB�GLV�#LOGS�IZ��EqKT�!Ud��VDD�#$0_T�
G�MՐCݱ��|@eM�RvC}�3�CHECAK0���0O�V!�kЙI��LE(!��P�ArpT�2K�W��0I�P2V!� h $ARIBiR� c�a�/�O�P8�ӐATT ��2�IF|@z�Aq4S��3UX����PL9I2V!� $g���OITCHx"[�W ��AS9�wSLL�BV!�� $�BA�DYs��BA�M!���Y9�PJ�5��Q��R6�V�Q_�KNOW�Cb��UF��AD�XV��0D�~+iPAYLOAt���Ic_��Rg�RgZ�OcL�q��PLCL=_�� !7��bP�QB��d���fF�iAC֠�js��d�I�h!Rؠ�g�ҢdB���љJ��q_J�a#���AND��Ĳ.t�bؤaL!q�PL0AL_ �P�0���QTրC��DNcE����J3CpWv� TPPDCK������>P�_ALPHgs�s�BE��gy|��K�1�� � �\��HoD_1Oj2ydDP�AR�*��;��&���TIA4U�5:U�6��MOM��a����n���{�Y�B� A�Da���n���{�PUB��R��҅n�҅{��/2�Wp��W � � PMsbT� �BxQ���� e$PI��81���TgJ��niJ�IV�Id�Ir��[��3!��>!��r�Ӫ�U3HIG�SU3�%�4� �4�%� ���"����!x
��!�%SAMP����^��_��%�P4s ю���[ 	ӝ� 3 ���0���&�C��� ��^��Sp��H&0	�IN�SpB�������"��6��6�V�GA�MM�SyI�� E�Tْ��;�D�tA�
�$ZpIBR!62I.T�$HIِ_���$C�˶E��ظAҾ���LWͽ�
���7Ơ��rЖ,0�qC�%C�HK��" �~I_A�����Rr� Rqܥ�Ǚ��ԥ���Ws� �$�x �1���I7RCHk_D�!� RN{��#�LE��ǒ!,���x���90MSWF�L�$�SCR((1#00��R@��3]B�րç��a����َ0��P�I3A9�METHaO����%��AXH��XX0԰62ER)I��^�3��R�0$u�	��pF{�_���$?ⲣ1�L�L�_�a�OOP����wᲡN��APP:���F��`�@{���أRT�V�OBp�0T����;��� 1�I��� ��lr���RA�@MGA1o���SSV-�w�P_@CURg��;�GRO[0S_�SA�Q��Y�#NO�pC!"�tY�� Zolox�������!b��,��&�DO�1A���A ����Х��A���A"�0WS�c L"h�*�� � ��YQLH�qܧ��SrZ�]B�o�=�q�Ô�q_�C1��M_W���g���c�M� �`Vq�$Ap�x1o�3"�PMJ�,�� �'A� 9�!YWi:�$�LWQ |ai�tg�tg�tg{t� �N`���S��JSpX�0O�sRqZ���P� *�� ���M��������������PX��� ��5L�q_~R� |�q#(Y����& n��&{�Y�Z��'�&t���Q��D�#0��@�}`�$PQ�PMO�N_QUc� �{ 8�@QCOU��n%PQTH��HO�n^0HYS:PES�RF^0UEI0O��0O|T�  �0PGõz�RUN_TO�r@Oْ.�� PE`�5C��A<�IND}E�ROGRA�nP� 2g�NE_NO�4�5IT��0�0�INFO�1� p�Q�:A��$PA�B� (��SLE�QݖFAѕF@�6� OySy�T� 4�@�ENAB��0PT�ION.S%0ERV�E���G���1{BGC]F�A� @R0J$�Rq�2���R�H�O�G "�EDITN�1� �v�K�jޓʱE�NU0W�*XAUTu�-UCO�PY�ِN\����M�ѱNXP\[q�PRU�T9� _RN�@OUC�$G�2�T����$$CL`?0[��&������Г �P�S�@�X��PXK�QIGRTU��_�PA� _WRK 2 e��@ 0 � �5�QMoYh\Jo|m |l	�`�m�o��`��o�o�f�e�l}�aI�[ct'`BS�*� �1�Y� <7����� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P��b�t���������srC�C��LMT?0����s  dѴIN�ڿ�дPRE_EXE��)�Ƅ0jP���za'`DV��S��@e)�%s�elect_macro����kϤ�qt�IOCNVVB�� 5��P��USňw����0V 14kP $$p��a�|�`?���߰>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ ���$�ѰLARMRE?COV ^������LMDG ��Ь�LM_�IF ��d�  YST-04�0 Operat�ion mode AUTO S���ed TELEOP)�������9��K�]�o��, 
� ���#�8� ~ǘLINE 0Ǒ�قABORTED�ǖS/WORLD? 100 %������$��1��8�A��ATAǒؑ3��גؒ��i���į�֯��NGTOL � @� 	 A� |���ѰPPI�NFO ��� f�L�^�p����  ������k���ۿ ſ�����5��Y�C�iϏ�%���ٯ���� ������'�9�K�]��o߁ߓߙ�PPLI�CATION ?}t��|��HandlingToolǖ� 
V9.40�P/17���
�883ǀ����F0�	�549������>��7DF5�О��ǓNone���FRA�� 6�9��_ACTIV�E1�  �� �  ���ڀMOD���������CHGAP�ONL�� �O�UPL[�1	���� >�B�T�f���CUREQ 1
��W  Tp�p�p�	��������l����� ��������i3l��p����^H��A�t
?HTTHKY�F Xv|��* <N`����� ���//&/8/J/ \/�/�/�/�/�/�/�/ �/�/?"?4?F?X?�? |?�?�?�?�?�?�?�? OO0OBOTO�OxO�O �O�O�O�O�O�O__ ,_>_P_�_t_�_�_�_ �_�_�_�_oo(o:o Lo�opo�o�o�o�o�o �o�o $6H� l~������ �� �2�D���h�z� ������ԏ���
� �.�@���d�v�����������TO������DO_CLEAN����E�NM  �� p��������ɯۯv�DSPDR3YRL���HI��o�@��G�Y�k�}����� ��ſ׿����ϻ�MAX��,�呿���=�X,�<�9�<���PLUGG,�-�9���WPRC��Bm�q�6�(ϗ�O����/SEGF�K����  �m��G�Y�k�}ߏ�����LAP$�7ޡ ������+�=�O�a��s����� �TO�TAL_ƈ� �USWENU$�1� �������RGDIS�PMMC�d�CL�O�@@�1�O"��D��-�_STR�ING 1��
_�M��S���
��_ITEM1��  n����� ���� $6HZ l~��������I/O �SIGNAL���Tryout �Mode��In�pNSimula�ted��Out�`OVERR~!� = 100���In cycl�T��Prog OAborj��J�Status��	�Heartbea�t��MH Fa�ul��Aler �!/!/3/E/W/i/p{/�/�/�/ (� ��(����/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFO�/WORИ�~A�/XO �O�O�O�O�O __$_ 6_H_Z_l_~_�_�_�_p�_�_�_�^PO�� �"`�KoEoWoio{o �o�o�o�o�o�o�o /ASew��bDEV%n�p9o� ���#�5�G�Y�k� }�������ŏ׏������1�C�PALT�-j��OD������� ȟڟ����"�4�F� X�j�|�������į֯X�GRIB������ �6�H�Z�l�~����� ��ƿؿ���� �2�@D�V�h�z�����R�- ��&����������"� 4�F�X�j�|ߎߠ߲߀�����������PREGn�W���0�~� �������������  �2�D�V�h�z����������$�$ARG�_~@D ?	�����  	$$W	[]�$�:	��SBN_CO�NFIG�X�WqRCII_SAVE  $�zm��TCELL�SETUP �
%  OME_�IO$$%MO�V_H� ��RE�P��#��UTOB7ACK� 	tFRA:\D�� .D�z '`r�D�w� ��s  25�/11/29 20:26:16D�;D���#//h��C/j/|/�/�/�/�/D�X/�/??(? :?L?�/p?�?�?�?�? �?�?g? OO$O6OHO ZO�?~O�O�O�O�O�O\�O���  c_F�_\ATBCKCTL.TM�)_;_pM___q_8INIm���j~CMESSAG� �Qz �[ODE_D� �j��XO�p�_@PA�US6` !� , 	�; x:oHg,		2o loVo�ozo�o�o�o�o �o�o 
D.Pz}�d`TSK  �mw}_CUPDT��P�Wd�p�VXW?ZD_ENB�Tf
�vSTA�U�u���XISX UNT �2�vwy � 	� ������F��I����E��mD�R�������������p���D��R��F� ��� ��� '��W�� �I���������,�/�M[ET��2@��y �PQ�@���@�&K@���@��MU@zK�@��H��R�>caU=����=�ӌ<����>�f>�iz5�SCRD�CFG 1�Y ��w ����%�7�I�pD�Q�	ܟ������ϯ ��Z��~�;�M�_��q�������6���FG�R9��p�_ԳPNA�� 	FѶ_�ED�P1��� �
 �%-PEDT-¿ R�vυ��Es� -FE�D��;9/�>���  ����2�����B�  ����{�����j�����3��#� �G�Y���@G�ߠ�6�����4� �����Yި��Z�l������5K������ Y�t���&�8���\���6��d��Y�@� ���(��7�S 0wY�w��f����8�W��{�I Z��C/��2/���!9{/��//LZݤ/�?V/h/�/�/��CR ���?�?Tn?�? ?�2?�?V?԰!�NO_�DEL�ҲGE_�UNUSE޿дI�GALLOW 1��   (�*SYSTEM�*
�	$SER�V_GR[�@`REG�E$�C
��@�NUM�J�C�MP�MU?@
�LA�YK�
�PM�PAL�PUCYC10 N3^P!^YSULSU_�M5Ra�CLo_�TBOX�ORI�ECUR_��P�MPMCNV6V�P10I^�PT4DLI�p�_�I�	*PROGRA��DPG_MI!^Ko]`AL+ejoTe�]`B�o�N$F�LUI_RESU`9W�o�O�o�dMR�N�@�<�?�;M_ q������� ��%�7�I�[�m�� ������Ǐُ�����!�3�E�W�2BLAL_OUT �K����WD_ABO�R:PcO��ITR_�RTN  �$��빸�NONSTO��� lHCCF�S_UTIL ��̷CC_AU�XAXIS 3$� h}�j�|������ƽCE_RIA3_I`@�נ���FCFG �$�/�#��_L�IM�B2+� ��� � 	��B\T���$� 
Ԡ��)[�Z�%�/���b��[����� ��H�!�����L��(
5������PA�`GP7 1H������A�S�e�w�6�CCV� C7��J��]���p������� CU������������U���é�̩�ձ�Uߩ�������ę;���PCk������������������R��ɱ���������� D� DU!�!�!�!�� ��&?��HE@ONFIpCѷG_P�P1H� +EH��ߟ߱�����������C�KPA�US�Q1H�ף IR�S�H�A��e� ������������� �E�+�i�{�a����A?Iץ�MؐN�FO 1��� �3��$4��B�]���l��^��e���¤��C*p���*��� B�� Cة�0�T������GwhPb�O� �� ��LLECT_��!�����EN�+`�ʒ���NDEַ#�/��1234567890�"�A��/ҵHw��#)j��< i{��;��/� �/`/+/=/O/�/s/ �/�/�/�/�/�/8?? ?'?�?K?]?o?�?�?@�?�?O�?��$�� ��IO #&��"S▒O��O�O�O`GTR�2'DM(��^�?�NN��(oM Z��_M[OR)q3)H��7� �U3��Y�_�_�_�_�_P�[bR�kQ*H�,S�I?<�<Ѡ<cz�KFd����P,�� ;ϒo�o�o˿�o�oœh�UY@E�oS� �sja.�PDB.���4�cpmidbg03��Рs:��>uq�pz��v  E��>x��}.���}�`��|�<�m!gP���t��~f��������@ud1:��?��XqDEF �-��zC)*�c�O�buf.txt�J��|K�[`�/DM��>���R�A���MCiR20_{RCdX���hS21�����G���CzA�d4�A���A��A����Bj��B�a:C&8/�Cp
B�DW�C6��D
�r�D"�D��E��8D�)��E}�F5���F^F��aA���Ufg23DL�D�	>z�!� 2���}��yc
�@�x9��Ĵ  �D4G������ � E%q�F�֟ E�p�u�F��P E��fF�3H ��G�M��Ъ5�>�G33��?�xn9�:q@�Q5����R�pA?a��=L��<#�QU�@,�C�ϒ���RSMOFST +i������P_T1Ɠ4DM�A =ք�MODEg 5dm�@��	Q,�M;��%���?���<�M�>��Ͷ�TES�Tc�2i�`�R�6(�O�K�CN�AB����n� 8��\�n�C6dB���Cpp�s����p:d�QS ��� ����T��4�I7>����>B8m5$�RT�_c�PROG �%j%��d�1�h@N�USER��x�KE�Y_TBL  �e�����	
��� !"#$�%&'()*+,�-./(:;<=�>?@ABCc�G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~����������������������������������������������������������������������������>��͓���������������������������������耇����������������������4A8�LC�K��F�y��STA�T��2�X�_AL�M�����_AUT/O_DO�E��FDR 3:i�2hi�US�x��i�$g��A�� ����T* g�2� bf��/ �/9/;�*pm�P/z/ �~/h/�/�/�/�/�/ ?"=�G?Y?k?/|? �?L/�?�?�/�?�?O O�?*O@OvO�O6?�O �O�O~?�O	_�?*_$_ BOD_6_p_~_T_�_�_ �_�_�Oo)o;o�OLo qo_�o�o�_�o�o�o �o�o�oFXo ��No���o�� ��@�N�$�b�x� ����n������ A��b�\�z�|�n��� ����ʟ���(�֏O� a�s������T�ʯį ��֯����2�H� ~���>���ɿۿ��� ϼ�2�,�J�L�>�x� ��\Ϛϰ����Ϧ�� 1�C��T�y�$Ϛߔ� �ϴߦ��������� N�`�߇���V߼� ���������H� V�,�j�������v��� ��$I��jd ���v����� 0��Wi{&� �\�����/ &/�:/P/�/�/F�/ �/�/��/?�:?4? R/T?F?�?�?d?�?�? �? O�/'O9OKO�/\O �O,?�O�O�?�O�O�O �O�O
_ _V_h_O�_ �_�_^O�_�_�O
oo "_$ooPo^o4oro�o �o�o~_�o	�_, Q�_rl�o�~� ����&�8��o_� q���.����dڏԏ ��� �.��B�X� ����N�ǟٟ럖��� !�̏B�<�Z�\�N��� ��l����������/� A�S���d���4����� ¯Ŀ�����Կ�(� ^�p���ϩϻ�f��� �Ϝ���*�,��X� f�<�zߐ����߆��� �#���4�Y��z�t� �ߔ����������� .�@���g�y���6�� ��l�����������( 6J`��V�� ����)��JD bdV��t�� �/�7/I/[/l/ �/<�/�/��/�/�/ ?�/?0?f?x?&/�? �?�?n/�?�?�/OO 2?4O&O`OnODO�O�O �O�O�?__+_�?<_ a_O�_|_�O�_�_�_ �_�_�_ o6oHo�Ooo �o�o>_�o�ot_�o�o o�o0>Rh ��^o����o� 1��oR�L�jl�^��� ��|���Џ���?� Q�c��t���D����� ҏԟƟ ���"�8� n���.�����˯v�ܯ ���"��:�<�.�h� v�L�����ֿ迖�� !�3�ޯD�i���τ� ���ϖ����ϴ���� >�P���w߉ߛ�FϬ� ��|�����
����8� F��Z�p���f��� ������9���Z�T� r�t�f�����������  ��GYk�| �L������� �*@v�6� ��~�	/�*/$/ BD/6/p/~/T/�/�/ �/�/�?)?;?�L? q?/�?�?�/�?�?�? �?�?�?OFOXO?O �O�ON?�O�O�?�O�O O__@_N_$_b_x_ �_�_nO�_�_o�Oo Ao�Obo\oz_|ono�o �o�o�o�o(�_O aso��To�� �o�����2�H� ~���>��ɏۏ�� ��2�,�J�L�>�x� ��\����������� 1�C��T�y�$����� ��������į�� N�`��������V��� ῌ�������H� V�,�jπ϶���v��� �߾�$�I���j�d� �τ�v߰߾ߔ����� �0���W�i�{�&ߌ� ��\������������ &���:�P�����F�� ����������:4 R�TF��d�� � ��'9K��\ �,������ ��
/ /V/h/�/ �/�/^�/�/�
?? "/$??P?^?4?r?�? �?�?~/�?	OO�/,O QO�/rOlO�?�O~O�O �O�O�O�O&_8_�?__ q_�_.O�_�_dO�_�_ �O�_�_ o.ooBoXo��otc�$CR_F�DR_CFG };re�Q?
UD1:�W�TJ�d  �`�\�bHIST 3<rf�  �`  �?�R@tA�tBtC�PpD�tEtItg�P�potw�_��bI�NDT_EN6p~�T�q��bT1_DO  1�U�u�sT2��w�VAR 2=�g�p hq  �{P�{P4�R��4�{��m[�:�RZ�`STO+����`TRL_DEL�ETNp�t ��_�SCREEN �re�rkcs�c�rUw�MMEN�U 1>��  <�\%�_��T ��R��S/�U���e� w�ğ������џ�	� B��+�x�O�a����� ������ͯ߯,��� b�9�K�q�������� ��ɿ����%�^�5� Gϔ�k�}��ϡϳ��� �����H��1�~�U� gߍ��ߝ߯������� 2�	��A�z�Q�c�� ����������.�� �d�;�M���q�������������YӃ_M�ANUAL{��rZCD�a?�y�rG� ���R�fx"
�"
?|(��P�dTGRP 2@:�y�B� � �s��� �$DwBCO�pRIG����v�G_ERRL�OG A��Q��I[m �N_UMLIM�s���u
�PXWOR/K 1B�8����//�}DBT;B_�� C%����S"� �aDB__AWAY��Q�GCP �r=���m"_AL�F�_�Y+����p�vk � 1D� , 
��/"�/%?/(c_M�pqw,@�=5�ONTIM���f�t�_6�)
�0~�'MOTNENFp�F�;RECORDw 2J� �-?�SG�O��1�?" x"!O3OEOWO�8_O�O �?�OO�O�O�O�O�O (_�OL_�Op_�_�_�_ A_�_9_�_]_o$o6o Ho�_lo�_�o�_�o�o �o�oYo}o2�oV hz��o��C �
��.��R��K� �������Џ?��ߏ �*�����+�b�t�� ������Ο=�O��� ��:�%���p�ߟ񟦯 ��O�ǯ�]������ H�Z���������#��5����ϩ�i"TO�LERENCv$B�ȿ"� L��� C�SS_CCSCB� 2K�\0" ?"{ϰϟ���7�� 
����@�R�d�3߈���"�x�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C�Ugy��� �������R�LL]�La�m1T#2� C�C�p�F�^ A�C�%pC���#�0�? 	 A����B���?�  ��$����\0����0��B��`#sߠK/]/o/�ϓ/��/�/s/�/�/�K����K�D���� �:U>:�?�Ȧ��/�Q�/`?;�@���O?�?�?�?Ȏ0A0F��?{F�A OO��7�1���9M	AB 
AZOdBAE�9$O�O�O��Oi:P��`�@0��DJCA� @5��
X-.
[N#_   M?�>O� ڴ�q_�_�_�_:W�A<o:[<ǲ/o�/�_+oPobotoL�eACHC�V�W-B$�Dz�cD�`�a =/�o�oo�oW�a.+�!��2=t,yD�"ŻYqC�z) I?�-t�s�js�w�y j�������Q���@`��$��� ��A����Bމ�o� �'�9��_]�o�N��� r���ɟ۟_�B�ʄ���YZ>`3�m$���0B�!�@�1�<%�R��Z�l�~����`_м¯� ��
���̯9�,�]�o� �� �H�����ٿ뿊� �ƿ3�E�W�iϬ��� $ϱ����� Ϟ���� /�A�S߶�w�V�h߭�`���S���ߐ�_ �f	��H�?�Q�~�u� ����������� �D��-�g�q����� ��������
@ 7Icm��߾�  �����) M@qdv�� �����//I/ P�m/�v/�/�/�/�/ �/�/�/?3?*?<?i? `?r?�?^/�?�?�?�? �?O/O&O8OJO\O�O��O�O�O�O�O�O�g	o  Q�PՄs �PC4p*p�p6U6P�\C9p/p��� ]V^PM]�6P�b:P�>P�VJ_�^P��bP�fP�Vr]v�	�Tp Q
k���_o�o�id1Q&oNo �;o_co�oˏUUA �  �o�k1Q@� � �o�k�b�����Up �� 1��>6��1C���C��cPfL��?#�c>_�{���`�cP��@@�d��r�`Be�cP>�s�qC��p癙��b�t<��o?�PH�)S�B�tq�q�p�r��`B���eIC��&�Q�4( �oz�UU�� �>��B��@�2�<���S}LQ��-R���?G����F�Bn����b��`ځ` � ?�p���U�[?����}t��$����$DCSS_CL�LB2 2M���p�P�^?�NSTCY 2N����  �������ʟ؟� ��� �2�D�Z�h�z� ������¯ԯ��SA��DEVICE 2%O��!�$��4& V�h�������˿¿Կ ���
�7�.�[�R�π�ϣϵ�����4(A�HNDGD P���*�Cz�A�LS 2Q��_�Q�c�u���ߙ߽߫���?�PA?RAM RP���1�`�&�RBT 2}T�� 8�P9<C�'p �qi�2l��s@"�R��(q�I�X��0�pB C7W  ��B\x�N�0�`Z����%��)���X�j��p����zq������B �(s,� F�p�V��q���b�,��B ��4&c �S� e�l�4+����H1�~����D�C�$Z��b����A,� 4�u@��X@��^@w����]B���B��cP%��C4��C3:^C4Ս�nЬ ��p8��-B{B���A���� l���C�C3��JC4jC3���yn+�3 D�ff 2�A PB W4+@:�]o� W�����/� /P/'/9/K/]/o/�/ �/�/�/?�/�/�/? #?5?�?Y?k?�?�?�o �?�?O�?6O!OZOlO WO�O�Es�?�?�?�O �O_�O�OL_#_5_G_ Y_k_}_�_�_�_ o�_ �_�_oo1o~oUogo �o�o�o�o�owO  D/Aze��� �O�o�o
��o��R� )�;���_�q������� ���ݏ�<��%�r� I�[�m��������ǟ ٟ&�8��\�G���k� ������گů���� �F��/�A�S�e�w� Ŀ������ѿ���� �+�x�O�aϮυϗ� �ϻ�����,���b� t�ﯘ߃߼ߧ����� ����:��C�U߂� Y�k��������� ��6���l�C�U�g� y����������� �� 	-?Q��� ����@+ dvQ����� ���*///%/r/ I/[/�//�/�/�/�/ �/&?�/?\?3?E?�? i?{?�?�?U�?�?"O 4OOXOCO|OgO�O{ ��?�O�?�O�O0__ _f_=_O_a_s_�_�_ �_�_�_o�_oo'o 9oKo�ooo�o�o�o�o �o�O:%^I�������H�$�DCSS_SLA�VE U��}�	���z?_4D  	���AR_MENU V	� �j�|�������ď�BY�� ���~?�SHOW 2}W	� � �b �aG�Q�X�v�������@��П֏���� @� :�d�a�s��������� �߯��*�$�N�K� ]�o�������̯ɿۿ ���8�5�G�Y�k� }Ϗ϶����������� "��1�C�U�g�yߠ� �߯��������	�� -�?�Q�c��s��� ����������)�;� M�t������������ ����%7Ip� m��������� �!3ZWi� ��J����/ /DA/S/e/��/� �/�/�/�/�/?./+? =?O?v/p?�/�?�?�? �?�?�??O'O9O`? ZO�?�O�O�O�O�O�O O�O_#_JOD_nOk_ }_�_�_�_�_�O�_�_ o4_.oX_Uogoyo�o �o�o�_�o�o�oo Bo?Qcu���o�:���CFG �X)�3�3q�5p�FRA:�\!�L+�%04d�.CSV|	p}�� �qA g�CHo�zv�	����
3q�����́܏�� ���4��JP�(���qp1� ��RC_OUT -Y��C���_C_FSI ?�i�  .�������͟���� �>�9�K�]������� ��ίɯۯ���#� 5�^�Y�k�}������� ſ�����6�1�C� U�~�yϋϝ������� ���	��-�V�Q�c� uߞߙ߽߫������� �.�)�;�M�v�q�� ����������� %�N�I�[�m������� ����������&!3 Eni{���� ���FAS e������� �//+/=/f/a/s/ �/�/�/�/�/�/�/? ?>?9?K?]?�?�?�? �?�?�?�?�?OO#O 5O^OYOkO}O�O�O�O �O�O�O�O_6_1_C_ U_~_y_�_�_�_�_�_ �_o	oo-oVoQoco uo�o�o�o�o�o�o�o .);Mvq� �������� %�N�I�[�m������� ��ޏُ���&�!�3� E�n�i�{�������ß ՟������F�A�S� e���������֯ѯ� ����+�=�f�a�s� ��������Ϳ���� �>�9�K�]φρϓ� ������������#� 5�^�Y�k�}ߦߡ߳� ���������6�1�C� U�~�y��������� ���	��-�V�Q�c� u��������������� .);Mvq� ����� %NI[m��� �����&/!/3/ E/n/i/{/�/�/�/�/��/�/�/3�$DC�S_C_FSO �?���71� P  ??T?}?x?�?�?�? �?�?�?OOO,OUO PObOtO�O�O�O�O�O �O�O_-_(_:_L_u_ p_�_�_�_�_�_�_o  oo$oMoHoZolo�o �o�o�o�o�o�o�o%  2Dmhz�� �����
��E� @�R�d���������Տ Џ����*�<�e� `�r���������̟�� ���=�8�J�\��������?C_RPI4>F?��������3?�&�o����� >SLү@d������ %�7�`�[�m�Ϩϣ� �����������8�3� E�W߀�{ߍߟ����� �������/�X�S� e�w��������� ���0�+�=�O�x�s� ������������ 'PK]o�� ������(# 5Gpk}��� ��Q���/6/1/C/ U/~/y/�/�/�/�/�/ �/?	??-?V?Q?c? u?�?�?�?�?�?�?�? O.O)O;OMOvOqO�O �O�O�O�O�O___ %_N_I_[_m_�_�_�_ �_�_�_�_�_&o!o3o Eonoio{o�o�o�o�o �o�o�oFAS e������>��NOCODE }ZU��?��PRE_CHK �\U��pA �p�< ��p�U�]�o�U� 	 < Q��������ۏ�Ǐ �#����Y�k�E��� ��{�şן��ß�� ��C�U�/�y�����s� ��ӯm���	���?� �+�u���a������� ɿ�Ϳ߿)�;��_� q�K�}ϧϝ������� ����%����[�m�G� �ߣ�}߯��߳���� !���E�W�1�c��g� y������������� A�S�-�w���c����� ��������+= asM_���� ��'�]o 	������ /#/�G/Y/3/e/�/ i/{/�/�/�/�/?�/ ?C?9Ky?�?%?�? �?�?�?�?	O�?-O?O OKOuOOOaO�O�O�O �O�O�O�O)_____ q_K_�_�_a?�_�_�_ �_o%o�_Io[o5oGo �o�o}o�o�o�o�o �o�oEW1{�g ���_����/� A��M�w�Q�c����� �����Ϗ�+��� a�s�M���������ߟ ���'���3�]�7� I������ɯۯ��� ����G�Y�3�}��� i���ſ�������� 1�C���+�yϋ�eϯ� �ϛ���������-�?� �c�u�Oߙ߫߅ߗ� �������)��M�_� U�G���A������ �������I�[�5�� ��k����������� ��3EQ{q�� ��]����/ AewQ��� ����/+//7/ a/;/M/�/�/�/�/�/ ��/?'??K?]?7? �?�?m??�?�?�?�? O�?5OGO!O3O}O�O iO�O�O�O�O�O�/�O 1_C_�Og_y_S_�_�_ �_�_�_�_�_o-oo 9oco=oOo�o�o�o�o �o�o�o__M_ �ok�o���� ����I�#�5�� ��k���Ǐ��ӏ��׏ �3�E��i�{�5c� ��ß�����ӟ�/� 	��e�w�Q������� ѯ㯽�ϯ�+��O� a�;��������Ϳ߿ y����!�K�%�7� �ϓ�mϷ��ϣ����� ����5�G�!�k�}�W� �߳ߩ������ߕ�� 1���g�y�S��� ���������-�� Q�c�=�o���s����� ��������M_ 9��o���� �7I#m Yk������ !/3/)/i/{//�/ �/�/�/�/�/�/?/? 	?S?e???q?�?u?�? �?�?�?OO�?%OOO E/W/�O�O1O�O�O�O �O__�O9_K_%_W_ �_[_m_�_�_�_�_�_ �_o5oo!oko}oWo �o�omO�o�o�o�o 1UgAS�� ����	���� Q�c�=�����s���Ϗ �o������;�M�'� Y���]�o���˟��� �۟�7��#�m�� Y������������ !�3�ͯ?�i�C�U��� ����տ������� 	�S�e�?ωϛ�uϧ���ϫϽ�������$DCS_SGN� ]	�E��-����29-�NOV-25 2�2:59 ��N�0�:27_�x�x�� [}�t��q��т�xҚك�JѨ��EƼÞ� �ۈǖ�  1�HO�W ^	�� x�/�VE�RSION �=�V4.5.�2��EFLOGI�C 1_���  	�����C���R�%�PROG_E_NB  ��:��{�s�ULSE  �X��%�_AC�CLIM������d��WRSTgJNT��E��-�EMO|�zя�$���INIT `2�����OPT_S�L ?		�	�
 	R575��V]�74b�6c�7c�50��1���C��|�@�TO  L��� �V�DEXҞ�dE�x�PA�TH A=�A�\k}��HCP�_CLNTID y?�:� D���ռ��IAG_G�RP 2e	�����z�	 �@�  
ff�?aG���BG�  2��/�8�[I@c�ς!��7@�z�@^��@
�!���mp2m15 �89012345�67���� � ?��?��=q?��
?���R?�Q�?ѯ�?�����?(�?�z����x�@�  A_�A�p !7A�8�8_�B4�� ��L�x�
�@����@��\@~��R@xQ�@q���@j�H@c��
@\��@U�@Mp��//�'$�; �O)H���@Ct >d 9���@4�/\)@)�� #t {@��/�/�/�/�/P'�?���?����_ ?}p�?u?n{?s ;?\�Q�? ?�2?D?V?h8�
=?�����0w5�z��H?p�h��?^�R�?�?�?�?��?h8��t0����@�?��0� ;@&O8OJO\OnOP' �$_�_Y_k_�O?_ �_�_�_�_�_s_�_�_ 1oCo!ogoyoo�o���Bj"� �2{1�@"?���f�t0�d"�5!�
u4V��u"�B3t�A>u��U?@[q��@`,�=q�=b���=�E1>�J��>�n�>��H�"<�o �z�s��q��� �x�C��@<(�Uz� �4�� ����A@x�?*�o��m*� P�b���tn���2����Ώ�����i>J���&�bN2�"�'�G�N��o@�@v�奈0����@f�fr!l ��33����(��"C��� ƒI�CH��)C.dB؃�"8"����' ���"~�A?�&"K���,�pf�B��@�p��������p�Ŀ`u������<�"����?`A�=s��=s��=.9ӿ~|�C� B��CC���xВ������3��N�T�����C0�T������Gw@�"����ǿ����ֿ���$��-=�+[��V���_��<��L����'�!�o��C�T_CONFIG� f��|��egY��ST�BF_TTS��
@����О�}���1��MAU������MS�W_CF��g� � # ��OCVIE�W��h!�-�� �s߅ߗߩ߻��ߟ� a�����,�>�P��� t�������]��� ��(�:�L�^���� ����������k�  $6HZ��~�� ����y 2 DVh�����X��v�RC�i���!�0./S/B/w/�f/�/�/�/��SBL�_FAULT �j*6��!GPMS�K���'��TDIAOG k��-�������UD1�: 6789012345I2��=1���%P\υ?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�Od696�I�r�
t?�O|�TREC	P"?4:
B44_[7M[ s?p_�_�_�_�_�_�_ �_ oo$o6oHoZolo�~o�o�O�O�O�o7�U�MP_OPTIO2=��.�aTR���:�)uPME���Y_TEMP  �È�3BG�rgp�B�QtUNI�����gq�YN_BR�K lL�7�EDITOR�a�a@�r�_
PENT 1m�)  ,&?TELEOP^P �z��pPSNA��:�&MTPG��p+�=��/����� z�����ۏ���� 5��Y�k�R���v��� ş���П����C� *�g�N�v�������������ޯ��?�Q����EMGDI_S�TAzuV�gq�uNC�_INFO 1n<!��b���X����������n�1o!� C��o����
�d�oU�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫���  u����
��*�B�*� P�b�t������� ������(�:�L�^� p���������2����� ��9�CUgy �������	 -?Qcu�� ������//1 ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?��? �?�?O)/OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�?�?�_�_o�_ 3O=oOoaoso�o�o�o �o�o�o�o'9 K]o����_�_ ����+o5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� �������ӟ���	� #�-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ����7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߹��������� �%�/�A�S�e�w�� ������������ +�=�O�a�s������� ���������'9 K]o����� ���#5GY k}�	����� �/1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? ��?�?�?�?/O)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�?�_�_�_ �_O�_!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �_�_����o� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o�������ɟ ۟���#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߝ��߹� ���������%�7�I� [�m��������� �����!�3�E�W�i� {��߇���������� /ASew� ������ +=Oas����� �����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?���?�?�?�?� �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�?�_ �_�_�_�?�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m�_u����_ ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�� ������u������ +�=�O�a�s������� ��ͯ߯���'�9� K�]�w���������ɿ �����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g߁� �ߝ߯���ۿ����	� �-�?�Q�c�u��� �����������)� ;�M�_�y߃������� ������%7I [m����� ��!3EWq� c��������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?i{�?�?�? �?��?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_�? s?}_�_�_�_�?�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qk_u�� ��_�����)� ;�M�_�q��������� ˏݏ���%�7�I� cQ���������ٟ ����!�3�E�W�i� {�������ïկ������/�A�[� �$�ENETMODE� 1p��_�  k�k��f�����j�OAT�CFG q�����Ѵ��C����DATA 1�rw�Ӱ���*	�*��'�9�K�]�"l�dlύ�e��� ����������'ߡ� ��]�o߁ߓߥ߷�1� ��U����#�5�G�Y� ���ߏ��������� ��u��1�C�U�g�y� �����)�������	 -����cu�����j�RPOS/T_LO��t�[�
׶#5Gi�R�ROR_PR� �%w�%L�XTA�BLE  w��ȟ����RSE�V_NUM ��?  ���  ��_AUTO_ENB  ���Xw_NO5! uw����"  *�*x �x �x �x + �+w �/�/�/Q$FLsTR=/O&HIS#�]�J+_ALM �1vw� �[x,e�+�/Q?c?u?��?�?�?�/_"W   w�v!���:j��TCP_VER �!w�!x�?$E{XT� _REQ�&s�H)BCSIZKO�=DSTKhIf%��?BTOL  �]Dz�"�A =D_BWD�0�@�&��A���CDI�A �wķ���]�KST�EP�O�Oj�POP�_DO�Oh�FDR_GRP 1xw��!d 	�?�_��yP�s�Y�Q'��M"���l���T� �����VyS�_�]yPAU���A��A���P�A1)l�BVJ@�[[A�?�P@����_k Ko6oooZoo�o�o�o�i<`�>@p��?�"�o�F@#c�`]?�G@�o(2�o�oZE�~�]p�u@S33�u�]@�q�g���yPq�|yPG� � @�Fg�fC�38RL��]?�pi�ޏ~6�X����8�75t��5��ߛ5`+��~�\�� m,�����[���&��e��e���FE�ATURE y����@��H�andlingT�ool �]�English �Dictiona�ry�4D St���ard��An�alog I/O�>�G�gle Sh�iftZ�uto �Software Update��matic Ba�ckup���gr�ound Edi�t ��Camer�aU�FY�CnrR�ndIm���om�mon caliOb UI��nˑ��Monitor�$�tr�Reli�abn��DHCP� �[�ata Ac�quis3�\�ia�gnos��R�v�i�splayΑLi�censZ�`�oc�ument Vi�ewe?�^�ual� Check S�afety��hanced����s�Frܐ�xt�. DIO /�f�i��@�end�E�rr>�L��\�4�s�[�rP�K� �@
�F�CTN Menu���vZ���TP I�n��facĵ�G�igE־�Đp �Mask Exc��g=�HT԰Pr?oxy Sv��igh-Spe��Ski�� Ť�O�m�munic��onsV�ur����q�V��ײconnect� 2��ncrְsGtru!��ʴ�eۡ���J���KARE�L Cmd. L��ua���Runw-Ti<�Env��^��el +��s��S/W�ƥ���r��Book(Sys�tem)
�MAC�ROs,M�/Of'fseu�p�HO����o�u�MR8�4���MechStop+�t����p�im�q���ax�R�����odo�witch�ӟ�y.��4�OptmF�,�fil䬳�g���p�ulti-T��Γ�PCM fun�Ǽ�o������^��Regie�rq���riݠF���S�Num Sel��|/�:� Adjua��*�W�q�h�tatu���ߪ�RDM �Robot�scgove'���ea���<�Freq An;lyq�Rem��O��n5�����Serv�oO�!��SNPX� b-�v�SN԰C�liܡ?r�Libr&�_�� ��q +�oJ�t��ssag���@ ����	�@�/Iս�MILI�B��P Fir�m���P��Acc<Ő͛TPTXk��eln���������orquo�imGula=��|u(��Pa&��ĐX�B�&�+�ev.���ri���TUSB poort �iPf��aݠ&R EVN�T� nexcept�����%5���VC�rl�c���V@���"�%q�+SR sSCN�/SGE�/��%UI	�Web Pl��>��A43���ۡ��ZDT A�pplj�
�{1EOAT����&0?�7Grid�񾡬=�?iR�".5� F����/גRX-10i�A/L�?Alar�m Cause/���ed(�All ?Smooth5��ОC�scii+�V�L�oad䠌JUpl��@w�toS ��r�ityAvoidM(�s7�t�@�ycn�����_�sCS+���. c��XJo���-T3_H��.RX��U���Xco�llabo����R�A�:�.9���in8���NRTHI
��On��e Hel�����ֿ�����1t�rU�ROS Eth$��A������;,��G �B�,|HUp0V�%�W�t ԰�_�iRS�ݐ�64M?B DRAM�o�c�FRO���L8F CFlD�����2M �A&:�opm�ԕex@V�F
�sh�q��wce�d�u��p��|tyn�sA�
�%�r����J���^�.v� P)Q/s�bS�`���O�N��mai��U���R�mq�T1�^FC+��%̋Fs9�ˌk̋n��Typ߽FC%��hױV�N Sp�FoarްK��Ԭ�lu!�x���cp�PG j��ҡ�RJ�[L`Su�p"}��֐f��c�rFP��lu� ��al�����r��i�
�q�4@а�ues�t,IMPLE  ׀6*|HZ���c0�BTea(�|���$�rtu���V�9HMqI�¤��UIFc�'pono2D�BC� :�L�y�p��������� ʿܿ	� ��?�6�H� u�l�~ϫϢϴ����� ����;�2�D�q�h� zߧߞ߰�������� 
�7�.�@�m�d�v�� �����������3� *�<�i�`�r������� ��������/&8 e\n����� ���+"4aX j������� �'//0/]/T/f/�/ �/�/�/�/�/�/�/#? ?,?Y?P?b?�?�?�? �?�?�?�?�?OO(O UOLO^O�O�O�O�O�O �O�O�O__$_Q_H_ Z_�_~_�_�_�_�_�_ �_oo oMoDoVo�o zo�o�o�o�o�o�o 
I@Rv� �������� E�<�N�{�r������� Տ̏ޏ���A�8� J�w�n�������џȟ ڟ����=�4�F�s� j�|�����ͯį֯� ���9�0�B�o�f�x� ����ɿ��ҿ����� 5�,�>�k�b�tφϘ� �ϼ��������1�(� :�g�^�p߂ߔ��߸� ������ �-�$�6�c� Z�l�~�������� ����)� �2�_�V�h� z��������������� %.[Rdv� ������! *WN`r��� ����//&/S/ J/\/n/�/�/�/�/�/ �/�/??"?O?F?X? j?|?�?�?�?�?�?�? OOOKOBOTOfOxO �O�O�O�O�O�O__ _G_>_P_b_t_�_�_ �_�_�_�_oooCo :oLo^opo�o�o�o�o �o�o	 ?6H Zl������ ���;�2�D�V�h� ������ˏԏ��� 
�7�.�@�R�d����� ��ǟ��П�����3� *�<�N�`�������ï ��̯����/�&�8� J�\�����������ȿ �����+�"�4�F�X� ��|ώϻϲ������� ��'��0�B�T߁�x� �߷߮���������#� �,�>�P�}�t��� �����������(� :�L�y�p��������� ������$6H ul~������  H5�52��21R�7850J6{14ATUP'�545'6VC�AMCRIbU�IF'28cNR�E52VR63�SCHLICޒDOCV�CS]U869'02�EIOC�4R{69VESET?vUJ7UR68�MASKPRXuY{7OCO#(�3?+ &3j&J�6%53�H�(L{CHR&OPLG?�0�&MHCRS&S��'MCS>0.'5=52MDSW+7u';OPu'MPRv&���(0&PCMzR�0q7+ 2� �'51�J51�80JPR�S"'69j&FRD�bFREQMC�N93&SNByA��'SHLBF�M1G�82&HT=C>TMIL��TPA�TPTXFcFELF� �8�J95�TU�Tv'95j&UEV�"&UECR&UFR�bVCC
XO�&V�IPnFCSC�FC�SG��IWE�B>HTT>R6���H;RVCGiWI�GQWIPGS�VRmCnFDGu'H7�7�R66J5'R��8R51
(6�(2��(5V�J8�86B�L=I% �84g�662R64N�VD"&R6�'R8�4�g79�(4�S�5i'J76j&D0��gF xRTSFC�R�gCRXv&CL9IZ8ICMS�Sp�>STYnG6)7C�TO>��7�NNj&ORS�&C &wFCB�FCF�7�CH>FCR"&F[CI�VFC�'J�PjO7GBfM�8OLax�ENDS&LU�&C�PR�7LWS�xC��STxTE�gS6�0FVR�IN�7IHaF�я��� ��+�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ��ɯۯ����#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E Wi{����� ��/ASe w������� //+/=/O/a/s/�/ �/�/�/�/�/�/?? '?9?K?]?o?�?�?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_�_�_�_�_ �_	oo-o?oQocouo �o�o�o�o�o�o�o );M_q�� �������%� 7�I�[�m���������Ǐُ�  �H552��2�1�R78�50��J614�AT�UP7�5457�6��VCAM�CR�I��UIF7�28n��NRE�52v�wR63�SCH��LICƚDOCV��CSU�869z7�0F�EIOCǛ�4�R69v�ES�ETW�u�J7u�R{68�MASK��PRXY��7�OCO��3W����6�m3�J65�536��H$�LCHƪOP�LGW�0�MHCuRǪS��MCSV��0��55F�MDS�W���OP��MP�R���6�06�PCM��R0E˓�F����6�51f�51��0nf�PRS��69��FRD��FREQn�MCN�936��SNBAכ%�SH�LB�ME��ּ2�6�HTCV�TMI�L�6�TPAV�T7PTX��ELړ��6�8%�#��J95n��TUT��95�wUEV��UECƪwUFR��VCCf��O��VIP��CS�C��CSGƚ$�I��WEBV�HTT�V�R6՜��S���C�G��IG��IPGmS'�RC��DG���H7��R66f�5t�u�R��R51f��6�2�5v�#�J׼��6��LU�5�s��v�4��66F�R6�4�NVD��R6n��R84�79��4��S5�J76��D0uFRT�S&�CR�CRX���CLI&�e�CMqSV�sV�STY��6�CTOV�#�V��75�NN�ORS�����6�FCBV�F�CF��CHV�FC�R��FCIF�FCR��J#��G
M�̻OL�ENDǪL]U��CPR��Lu��S�C$�StTE�S60�FVR6V�IN��IH��� m??�?�?�?�?�?�? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�_ �_�_�_�_�_oo+o =oOoaoso�o�o�o�o �o�o�o'9K ]o������ ���#�5�G�Y�k� }�������ŏ׏��� ��1�C�U�g�y��� ������ӟ���	�� -�?�Q�c�u������� ��ϯ����)�;� M�_�q���������˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���!�3�E�W�i�{� �ߟ߱���������� �/�A�S�e�w��� �����������+� =�O�a�s��������� ������'9K ]o������ ��#5GYk }������� //1/C/U/g/y/�/ �/�/�/�/�/�/	?? -???Q?c?u?�?�?�? �?�?�?�?OO)O;O MO_OqO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_�_�_ �_o!o3oEoWoio{o �o�o�o�o�o�o�o /ASew�� �������+� =�O�a�s����������͏ߏ�ST�D�LANG ���0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h��zߌߞ߰���RBT
�OPTN����� �'�9�K�]�o������������DPN 	���)�;�M�_�q� �������������� %7I[m� ������� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo 1oCoUogoyo�o�o�o �o�o�o�o	-? Qcu����� ����)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� ������ǟٟ���� !�3�E�W�i�{����� ��ïկ�����/� A�S�e�w��������� ѿ�����+�=�O� a�sυϗϩϻ����� ����'�9�K�]�o� �ߓߥ߷��������� �#�5�G�Y�k�}�� ������������� 1�C�U�g�y������� ��������	-?Qc�f�������99��$�FEAT_ADD ?	����  	 �#5GYk}� ������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ���������DEMO� y   �L�B�T߁�x� �߷߮���������� �G�>�P�}�t��� �����������C� :�L�y�p��������� ������?6H ul~����� �;2Dqh z������ / 
/7/./@/m/d/v/�/ �/�/�/�/�/�/?3? *?<?i?`?r?�?�?�? �?�?�?�?O/O&O8O eO\OnO�O�O�O�O�O �O�O�O+_"_4_a_X_ j_�_�_�_�_�_�_�_ �_'oo0o]oTofo�o �o�o�o�o�o�o�o# ,YPb��� �������(� U�L�^����������� ʏ����$�Q�H� Z���~�������Ɵ�� ��� �M�D�V��� z�������¯ܯ�� 
��I�@�R��v��� ������ؿ���� E�<�N�{�rτϱϨ� ���������A�8� J�w�n߀߭ߤ߶��� ������=�4�F�s� j�|��������� ���9�0�B�o�f�x� �������������� 5,>kbt�� �����1( :g^p���� ��� /-/$/6/c/ Z/l/�/�/�/�/�/�/ �/�/)? ?2?_?V?h? �?�?�?�?�?�?�?�? %OO.O[OROdO�O�O �O�O�O�O�O�O!__ *_W_N_`_�_�_�_�_ �_�_�_�_oo&oSo Jo\o�o�o�o�o�o�o �o�o"OFX �|������ ���K�B�T���x� ������ۏҏ��� �G�>�P�}�t����� ��ןΟ�����C� :�L�y�p�������ӯ ʯܯ	� ��?�6�H� u�l�~�����Ͽƿؿ ����;�2�D�q�h� zϔϞ���������� 
�7�.�@�m�d�vߐ� ���߾��������3� *�<�i�`�r����� ���������/�&�8� e�\�n����������� ������+"4aX j������� �'0]Tf� �������#/ /,/Y/P/b/|/�/�/ �/�/�/�/�/??(? U?L?^?x?�?�?�?�? �?�?�?OO$OQOHO ZOtO~O�O�O�O�O�O �O__ _M_D_V_p_ z_�_�_�_�_�_�_o 
ooIo@oRolovo�o �o�o�o�o�o E<Nhr��� ������A�8� J�d�n�������яȏ ڏ����=�4�F�`� j�������͟ğ֟� ���9�0�B�\�f��� ����ɯ��ү����� 5�,�>�X�b������� ſ��ο����1�(� :�T�^ϋςϔ��ϸ� ������ �-�$�6�P� Z߇�~ߐ߽ߴ����� ����)� �2�L�V�� z������������ %��.�H�R��v��� ������������! *DN{r��� ����&@ Jwn����� ��//"/</F/s/ j/|/�/�/�/�/�/�/ ???8?B?o?f?x? �?�?�?�?�?�?OO O4O>OkObOtO�O�O��O�O�O�O__0]  'XF_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |������� ��0�B�T�f�x��� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
�|�.�  /� )�J�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x��������������� ,>Pbt� ������ (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�?�? �?
OO.O@OROdOvO �O�O�O�O�O�O�O_ _*_<_N_`_r_�_�_ �_�_�_�_�_oo&o 8oJo\ono�o�o�o�o �o�o�o�o"4F Xj|����� ����0�B�T�f� x���������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ ؿ���� �2�D�V� h�zόϞϰ������� ��
��.�@�R�d�v� �ߚ߬߾�������� �*�<�N�`�r��� �����������&� 8�J�\�n��������� ��������"4F Xj|����� ��0BTf x������� //,/>/P/b/t/�/ �/�/�/�/�/�/?? (?:?L?^?p?�?�?�? �?�?�?�? OO$O6O HOZOlO~O�O�O�O�O �O�O�O_ _2_D_V_ h_z_�_�_�_�_�_�_ �_
oo.o@oRodovo �o�o�o�o�o�o�o *<N`r�� �������&� 8�J�\�n��������� ȏڏ����"�4�F� X�j�|�������ğ֟ �����0�B�T�f� x���������ү��� ��,�>�P�b�t��� ������ο���� (�:�L�^�pςϔϦ� �������� ��$�4�8�+�N�`�r߄� �ߨߺ��������� &�8�J�\�n���� �����������"�4� F�X�j�|��������� ������0BT fx������ �,>Pbt �������/ /(/:/L/^/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n��� ������"�4� F�X�j�|�������ď ֏�����0�B�T� f�x���������ҟ� ����,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D� V�h�zߌߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N�`�r��� ������������ &8J\n��� �����"4 FXj|���� ���//0/B/T/ f/x/�/�/�/�/�/�/ �/??,?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O �O�O�O�O�O __$_�6Y�$FEAT_�DEMOIN  �;T�fP�<P�NTINDEX[[�jQ�NPILECO�MP z����QiRIU�P�SETUP2 �{�U�R� � N �Q�S_AP2BCK 1|�Y?  �)7Xo"k%�_8o<P�P&o co9U�_�oo�oBo�o �oxo�o1C�og �o��,�P�� ���?��L�u�� ��(���Ϗ^�󏂏� )���M�܏q������ 6�˟Z�؟���%��� I�[��������D� ٯh������3�¯W� �d������@�տ� v�Ϛ�/�A�пe��� �ϛ�*Ͽ�N���r��� ߨ�=���a�s�ߗ� &߻���\��߀��'� ��K���o���|��4� ��X������#���G� Y���}������B����f�����1�Y�PP��_ 2�P*.cVR8���*��������l PC����FR6:D�2�V�TzP z�w�]PG���*.Fo/��	�:,�^/�STMi/�/ /"�-M/�/�H�/?��'?�/�/g?�GIFq?�?�%�?D?V?�?�JPG�?O�%O0�?�?oO�
JSyO�O���5C�OMO%
J�avaScript�O�?CS�O&_�&�_�O %Cas�cading S�tyle She�etsR_��
AR�GNAME.DT�_��� \�_S_�A��T�_�_�PDISP*�_���To�_��QLaZooCLL�B.ZIwo2o$ :�\�a\�o�i�AC?ollabo�o�o�
TPEINS.gXML�_:\!�[o�QCustom� Toolbar�biPASSWO�RDQo��FRS�:\�dB`Pas�sword Config���/�� (�e��������N� �r�����=�̏a� �����&���J���� �����9�K�ڟo��� ����4�ɯX��|��� #���G�֯@�}���� 0�ſ׿f������1� ��U��y��ϯ�>� ��b���	ߘ�-߼�Q� c��χ�߽߫�L��� p��ߦ�;���_��� X��$��H�����~� ���7�I���m����  �2���V���z���! ��E��i{
�. ��d���� S�wp�<� `�/�+/�O/a/ ��//�/8/J/�/n/ ?�/�/9?�/]?�/�? �?"?�?F?�?�?|?O �?5O�?�?kO�?�OO �O�OTO�OxO__�O C_�Og_y__�_,_�_ P_b_�_�_o�_oQo �_uoo�o�o:o�o^o �o�o)�oM�o�o ��6��l� �%�7��[�����  ���D�ُh�z���� 3�,�i���������ßR��v�������$FILE_DG�BCK 1|������� < �)
S�UMMARY.DyG!�͜MD:U����ِDiag� Summary�����
CONSLOG��n���ٯ����Console� log���	T�PACCN�t�%�\�����TP A�ccountin�;���FR6:I�PKDMP.ZI	PͿј
�ϥ����Exceptio�n"�ӻ��MEMCHECK���������-�Memory� Data�����Bn )��RIP�E�~ϐ�%ߴ�%��� Packe�t L:���L�$y�c���STAT���߭� %~A�Status��^�	FTP�����	��/�mmen�t TBD2�^� �>I)ETHERNEw�
�d�u�����Ethern�J�1�figura�Aϩ��DCSVRAF&���7������ verify �all:����4=��DIFF/���'���;�Q�diff��r�d���CHG01������A����it�2���270 ���fx3���I �p��VTRNDIAG.LSu&8�z��� Ope���L� ��nosti�c��`�)VwDEV�DAT������Vis~�Device�+IMG��,/>/��/:�i$Imag�u/+UP ES�/�/FRS:\�?Z=��Upda�tes List�Z?��� FLEXEVEN��/�/�?����1 UIF �EvM�M���-v�Z)CRSEN�SPK�/˞�\�!O���CR_TAO?R_PEAKbOͩ�PSRBWLD.CM�O͜E2�O\?�.�PS_ROBO�WELS���:GI�G��@_�?d_��G�igE�(O��N��@�)UQHAD�OW__D_V_�_���Shadow C�hange����.�dt�RRCMERAR�_�_�_oo��4`�CFG Erro�ro tailo �MA�k�CMSGLIBgoNo`o�o0|R�e��z0ic�o�ao�)�`ZD0_pO�os��ZD�P�ad�l �RNOTI�Rd����Notificx����,�AG�� P�ӟt���������Ώ ]�����(���L�^� 폂������G�ܟk�  ����6�şZ��~� �����C�د�y�� ��2�D�ӯh������ ��¿Q��u�
�ϫ� @�Ͽd�v�Ϛ�)Ͼ� ��_��σ�ߧ�%�N� ��r�ߖߨ�7���[� ����&��J�\��� ����3����i��� ��"�4���X���|��� ���A�����w��� 0��=f���� �O�s�> �bt�'�K ���/�:/L/� p/��/�/5/�/Y/�/  ?�/$?�/H?�/U?~? ?�?1?�?�?g?�?�?  O2O�?VO�?zO�OO �O?O�OcO�O
_�O._ �OR_d_�O�__�_�_ M_�_q_oo�_<o�_ `o�_mo�o%o�oIo�o �oo�o8J�on �o��3�W�{ �"��F��j�|�� ��/�ď֏e�������0��$FILE_�FRSPRT  ��������?�MDO?NLY 1|S��� 
 �)�MD:_VDAEXTP.ZZZ1��⏹�ț6%�NO Back �file ���S�6P�����>�� K�t�����'���ί]� 򯁯�(���L�ۯp� �����5�ʿY�׿ � ��$ϳ�H�Z��~�� �ϴ�C���g���ߝ� 2���V���cߌ�߰� ?�����u�
��.�@����d��߈��C�VI�SBCKq�[����*.VD����S��FR:\��ION?\DATA\��v��S�Vision VD���Y� k����y��B����� x���1C��g�� �,�P��� �?�Pu� (��^��/� �M/�q/�/>/�/6/ �/Z/�/?�/%?�/I? [?�/??�?2?D?�?�9�LUI_CON�FIG }S�����; $ �3v�{S�;OMO_OqO0�O�O�I#@|x�?�O �O�O__%\�OH_Z_ l_~_�_'_�_�_�_�_ �_o�_2oDoVohozo �o#o�o�o�o�o�o
 �o.@Rdv� �������*� <�N�`�r�������� ̏ޏ�����&�8�J� \�n��������ȟڟ 쟃���"�4�F�X�j� �������į֯�� ��0�B�T�f����� ������ҿ�{��� ,�>�P�b����ϘϪ� ������w���(�:� L�^��ςߔߦ߸��� ��s� ��$�6�H��� Y�~������]��� ��� �2�D���h�z� ��������Y�����
 .@��dv�� ��U��* <�`r���� Q��//&/8/� \/n/�/�/�/;/�/�/ �/�/?"?�/F?X?j? |?�?�?7?�?�?�?�? OO�?BOTOfOxO�O �O3O�O�O�O�O__ �O>_P_b_t_�_�_/_ �_�_�_�_oo�_:o�Lo^opo�o�o$h � x�o�c�$F�LUI_DATA ~����a�(a�dR�ESULT 3��ep �T��/wizar�d/guided�/steps/Expert�o=O as���������z�Cont�inue wit�h Gpance �:�L�^�p�������`��ʏ܏� � �b�-�a�e�0 ��0`��c�a?��ps��������� ҟ�����,�>�P� �0ow���������ѯ �����+�=�O�a��?�1�C�U�e�cllbs�ֿ����� 0�B�T�f�xϊϜ�[� ����������,�>� P�b�t߆ߘߪ�i�{���ߟ�]�e�rip (pſ-�?�Q�c�u�� ������������ )�;�M�_�q������� ���������������`�e�#pTimeUS/DST	 ��������!3E�Enabl(�y���� ���	//-/?/Q/�b�)�/M_q24|�/�/?? )?;?M?_?q?�?�?T f�?�?�?OO%O7O IO[OmOO�O�Ob/t/��/�/Z�"qRegion�O5_G_Y_k_ }_�_�_�_�_�_�_��America !�#o5oGoYoko}o�o��o�o�o�o�o��Ay��O�O3�O_qEditor�o��� ������+�=�� � Touch �Panel rs �(recommenp�)K�������Ə ؏���� �2�D�|��%��I[qaccesoܟ� � �$�6�H�Z�l�~������Connec�t to Network��֯��� ��0�B�T�f�x�����x��@��}����,!��s Introduct!_4�F� X�j�|ώϠϲ����� �����0�B�T�f� xߊߜ߮��������� ɿ��"� i�{���������� ����/�A� �e�w� ��������������+=�H�3��+�O���� � 2DVhz �K������
/ /./@/R/d/v/�/�/ Yk}�/�??*? <?N?`?r?�?�?�?�? �?�?��?O&O8OJO \OnO�O�O�O�O�O�O �O�/_�/1_�/X_j_ |_�_�_�_�_�_�_�_ oo0oBoS_foxo�o �o�o�o�o�o�o ,>�O_!_�E_� ������(�:� L�^�p�����So��ʏ ܏� ��$�6�H�Z� l�~���O��s՟� ��� �2�D�V�h�z� ������¯ԯ毥�
� �.�@�R�d�v����� ����п⿡��ş'� 9���`�rτϖϨϺ� ��������&�8��� \�n߀ߒߤ߶����� �����"�4��=�� a��Mϲ��������� ��0�B�T�f�x��� I߮��������� ,>Pbt�E�� i����(: L^p����� ��� //$/6/H/Z/ l/~/�/�/�/�/�/� ���/?�V?h?z? �?�?�?�?�?�?�?
O O.O�ROdOvO�O�O �O�O�O�O�O__*_ <_�/??�_C?�_�_ �_�_�_oo&o8oJo \ono�o?O�o�o�o�o �o�o"4FXj |�M___q_��_� ��0�B�T�f�x��� ������ҏ�o��� ,�>�P�b�t������� ��Ο�����%�� L�^�p���������ʯ ܯ� ��$�6�G�Z� l�~�������ƿؿ� ��� �2��S��w� 9��ϰ���������
� �.�@�R�d�v߈�G� �߾���������*� <�N�`�r��Cϥ�g� ��ύ���&�8�J� \�n������������� ����"4FXj |�������� ��-��Tfx� ������// ,/��P/b/t/�/�/�/ �/�/�/�/??(?� 1U??A�?�?�? �?�? OO$O6OHOZO lO~O=/�O�O�O�O�O �O_ _2_D_V_h_z_ 9?�?]?�_�_�?�_
o o.o@oRodovo�o�o �o�o�o�O�o* <N`r���� ��_�_�_�_#��_J� \�n���������ȏڏ ����"��oF�X�j� |�������ğ֟��� ��0����u�7� ������ү����� ,�>�P�b�t�3����� ��ο����(�:� L�^�pς�A�S�e��� ���� ��$�6�H�Z� l�~ߐߢߴ��߅��� ��� �2�D�V�h�z� ������������ ���@�R�d�v����� ����������* ;�N`r���� ���&��G 	�k-������ ��/"/4/F/X/j/ |/;�/�/�/�/�/�/ ??0?B?T?f?x?7 �?[�?�?�?OO ,O>OPObOtO�O�O�O �O�O�/�O__(_:_ L_^_p_�_�_�_�_�_ �?�_�?o!o�OHoZo lo~o�o�o�o�o�o�o �o �ODVhz �������
� ��_%o�_I�s�5o�� ����Џ����*� <�N�`�r�1������ ̟ޟ���&�8�J� \�n�-�w�Q���ů�� ����"�4�F�X�j� |�������Ŀ����� ��0�B�T�f�xϊ� �Ϯ����������� ٯ>�P�b�t߆ߘߪ� ����������տ:� L�^�p������� ���� ��$������ i�+ߐ����������� �� 2DVh'� �������
 .@Rdv5�G� Y��}���//*/ </N/`/r/�/�/�/�/ y�/�/??&?8?J? \?n?�?�?�?�?�?� �?�O�4OFOXOjO |O�O�O�O�O�O�O�O __/OB_T_f_x_�_ �_�_�_�_�_�_oo �?;o�?_o!O�o�o�o �o�o�o�o(: L^p/_���� �� ��$�6�H�Z� l�+o��Oo��sou�� ��� �2�D�V�h�z� ����������
� �.�@�R�d�v����� ����}�߯����ٟ <�N�`�r��������� ̿޿���ӟ8�J� \�nπϒϤ϶����� �����ϯ��=�g� )��ߠ߲��������� ��0�B�T�f�%ϊ� ������������� ,�>�P�b�!�k�Eߏ� ��{�����(: L^p����w� �� $6HZ l~���s����� ��/��2/D/V/h/z/ �/�/�/�/�/�/�/
? �.?@?R?d?v?�?�? �?�?�?�?�?OO� ��]O/�O�O�O�O �O�O�O__&_8_J_ \_?�_�_�_�_�_�_ �_�_o"o4oFoXojo )O;OMO�oqO�o�o�o 0BTfx� ��m_����� ,�>�P�b�t������� ��{oݏ�o��o(�:� L�^�p���������ʟ ܟ� ��#�6�H�Z� l�~�������Ưد� ���͏/��S��z� ������¿Կ���
� �.�@�R�d�#��Ϛ� �Ͼ���������*� <�N�`����C���g� i�������&�8�J� \�n�����u��� �����"�4�F�X�j� |�������q������� 	��0BTfx� �������� ,>Pbt��� ����/���� 1/[/�/�/�/�/�/ �/�/ ??$?6?H?Z? ~?�?�?�?�?�?�? �?O O2ODOVO/_/ 9/�O�Oo/�O�O�O
_ _._@_R_d_v_�_�_ �_k?�_�_�_oo*o <oNo`oro�o�o�ogO yO�O�O�o�O&8J \n������ ���_"�4�F�X�j� |�������ď֏��� ��o�o�oQ�x��� ������ҟ����� ,�>�P��t������� ��ί����(�:� L�^��/�A���e�ʿ ܿ� ��$�6�H�Z� l�~ϐϢ�a������� ��� �2�D�V�h�z� �ߞ߰�o��ߓ��߷� �.�@�R�d�v��� �����������*� <�N�`�r��������� ��������#��G 	�n������ ��"4FX� |������� //0/B/T/u/7 �/[]/�/�/�/?? ,?>?P?b?t?�?�?�? i�?�?�?OO(O:O LO^OpO�O�O�Oe/�O �/�O�O�?$_6_H_Z_ l_~_�_�_�_�_�_�_ �_�? o2oDoVohozo �o�o�o�o�o�o�o�O _�O%O_v�� �������*� <�N�or��������� ̏ޏ����&�8�J� 	S-w���cȟڟ ����"�4�F�X�j� |�����_�į֯��� ��0�B�T�f�x��� ��[�m����󿵟� ,�>�P�b�tφϘϪ� �������ϱ��(�:� L�^�p߂ߔߦ߸��� ���� ￿ѿ�E�� l�~���������� ��� �2�D��h�z� ��������������
 .@R�#�5� Y����* <N`r��U�� ���//&/8/J/ \/n/�/�/�/c�/� �/�?"?4?F?X?j? |?�?�?�?�?�?�?�? ?O0OBOTOfOxO�O �O�O�O�O�O�O�/_ �/;_�/b_t_�_�_�_ �_�_�_�_oo(o:o LoOpo�o�o�o�o�o �o�o $6H_ i+_�O_Q��� �� �2�D�V�h�z� ����]oԏ���
� �.�@�R�d�v����� Y��}ߟ񟵏�*� <�N�`�r��������� ̯ޯ𯯏�&�8�J� \�n���������ȿڿ 쿫���ϟ�C��j� |ώϠϲ��������� ��0�B��f�xߊ� �߮����������� ,�>���G�!�k��W� ����������(�:� L�^�p�����S߸��� ���� $6HZ l~�O�a�s��� �� 2DVhz ��������
/ /./@/R/d/v/�/�/ �/�/�/�/�/��� 9?�`?r?�?�?�?�? �?�?�?OO&O8O� \OnO�O�O�O�O�O�O �O�O_"_4_F_?? )?�_M?�_�_�_�_�_ oo0oBoTofoxo�o IO�o�o�o�o�o ,>Pbt��W_ �{_��_��(�:� L�^�p���������ʏ ܏���$�6�H�Z� l�~�������Ɵ؟� ���/��V�h�z� ������¯ԯ���
� �.�@���d�v����� ����п�����*� <���]����C�EϺ� ��������&�8�J� \�n߀ߒ�Q������� �����"�4�F�X�j� |��Mϯ�q������ ��0�B�T�f�x��� ������������ ,>Pbt��� ���������7 ��^p����� �� //$/6/��Z/ l/~/�/�/�/�/�/�/ �/? ?2?�;_? �?K�?�?�?�?�?
O O.O@OROdOvO�OG/ �O�O�O�O�O__*_ <_N_`_r_�_C?U?g? y?�_�?oo&o8oJo \ono�o�o�o�o�o�o �O�o"4FXj |�������_ �_�_-��_T�f�x��� ������ҏ����� ,��oP�b�t������� ��Ο�����(�:� ����A�����ʯ ܯ� ��$�6�H�Z� l�~�=�����ƿؿ� ��� �2�D�V�h�z� ��K���o��ϓ���
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ���������#���J� \�n������������� ����"4��Xj |������� 0��Q�u7� 9�����// ,/>/P/b/t/�/E�/ �/�/�/�/??(?:? L?^?p?�?A�?e�? �?�/ OO$O6OHOZO lO~O�O�O�O�O�O�/ �O_ _2_D_V_h_z_ �_�_�_�_�_�?�?�? o+o�?Rodovo�o�o �o�o�o�o�o* �ON`r���� �����&��_/o 	oS�}�?o����ȏڏ ����"�4�F�X�j� |�;����ğ֟��� ��0�B�T�f�x�7� I�[�m�ϯ������ ,�>�P�b�t������� ��ο�����(�:� L�^�pςϔϦϸ��� �ϛ�����!��H�Z� l�~ߐߢߴ������� ��� �߿D�V�h�z� ������������
� �.������s�5ߚ� ����������* <N`r1��� ���&8J \n�?��c���� ��/"/4/F/X/j/ |/�/�/�/�/�/��/ ??0?B?T?f?x?�? �?�?�?�?��?�O �>OPObOtO�O�O�O �O�O�O�O__(_�/ L_^_p_�_�_�_�_�_ �_�_ oo$o�?EoO io+O-o�o�o�o�o�o �o 2DVhz 9_������
� �.�@�R�d�v�5o�� Yo��͏����*� <�N�`�r��������� ̟����&�8�J� \�n���������ȯ�� я������F�X�j� |�������Ŀֿ��� ��ݟB�T�f�xϊ� �Ϯ����������� ٯ#���G�q�3��ߪ� ����������(�:� L�^�p�/ϔ����� ���� ��$�6�H�Z� l�+�=�O�a������� �� 2DVhz ��������
 .@Rdv�� ���������/�� </N/`/r/�/�/�/�/ �/�/�/??�8?J? \?n?�?�?�?�?�?�? �?�?O"O��/gO )/�O�O�O�O�O�O�O __0_B_T_f_%?w_ �_�_�_�_�_�_oo ,o>oPoboto3O�oWO �o{O�o�o(: L^p����� �o� ��$�6�H�Z� l�~�������Ə�o� �o��o2�D�V�h�z� ������ԟ���
� ��@�R�d�v����� ����Я�����׏ 9���]��!������� ̿޿���&�8�J� \�n�-��Ϥ϶����� �����"�4�F�X�j� )���M����߅����� ��0�B�T�f�x�� ������������ ,�>�P�b�t������� ��{��ߟ�����: L^p����� �� ��6HZ l~������ �/����;/e/' �/�/�/�/�/�/�/
? ?.?@?R?d?#�?�? �?�?�?�?�?OO*O <ONO`O/1/C/U/�O y/�O�O__&_8_J_ \_n_�_�_�_�_u?�_ �_�_o"o4oFoXojo |o�o�o�o�o�O�O�O 	�O0BTfx� ��������_ ,�>�P�b�t������� ��Ώ������o�o �o[���������ʟ ܟ� ��$�6�H�Z� �k�������Ưد� ��� �2�D�V�h�'� ��K���o�Կ���
� �.�@�R�d�vψϚ� �Ͼ�Ͽ������*� <�N�`�r߄ߖߨߺ� y��ߝ�����&�8�J� \�n��������� �������4�F�X�j� |��������������� ��-��Q�� ������ ,>Pb!���� ����//(/:/ L/^//A�/�/y �/�/ ??$?6?H?Z? l?~?�?�?�?s�?�? �?O O2ODOVOhOzO �O�O�Oo/�/�/�O_ �/._@_R_d_v_�_�_ �_�_�_�_�_o�?*o <oNo`oro�o�o�o�o �o�o�o�O_�O/ Y_������ ���"�4�F�X�o |�������ď֏��� ��0�B�T�%7 I��mҟ����� ,�>�P�b�t������� i�ί����(�:� L�^�p���������w� ��������$�6�H�Z� l�~ϐϢϴ������� �ϻ� �2�D�V�h�z� �ߞ߰���������
� ɿۿ�O��v��� �����������*� <�N��_��������� ������&8J \�}?�c��� ��"4FXj |������� //0/B/T/f/x/�/ �/�/m�/��/�? ,?>?P?b?t?�?�?�? �?�?�?�?O�(O:O LO^OpO�O�O�O�O�O �O�O _�/!_�/E_? 	_~_�_�_�_�_�_�_ �_o o2oDoVoOzo �o�o�o�o�o�o�o
 .@R_s5_� �mo�����*� <�N�`�r�������go ̏ޏ����&�8�J� \�n�������c�� џ���"�4�F�X�j� |�������į֯��� ���0�B�T�f�x��� ������ҿ������� ٟ#�M��tφϘϪ� ����������(�:� L��p߂ߔߦ߸��� ���� ��$�6�H�� �+�=ϟ�a������� ��� �2�D�V�h�z� ����]���������
 .@Rdv����k�}�����$�FMR2_GRP� 1���� �C4 w B��	 ���9K6F@ �a@�6G�  ��Fg�fC�8yR�y?�  ���66�X����875t��5����5`+�yAg�  /+BH�<w-%@S339%�!5[/l-6@6!�/ xl/�/�/�/�/?�/ &??J?5?G?�?k?�?���_CFG �TK�?�? OO��9NO �
F0FA K@�<R�M_CHKTYP  ��$&� �ROMa@_MI�Ng@�����@��R XSSB�3��� �7�O���C�O�O�5T�P_DEF_OW�  ��$WI�RCOMf@_�$�GENOVRD_�DO�F��E]TH���D dbUdKT_�ENB7_ KPRWAVC��G�@ �Y�O�_�?o�yo&oI* �V�QOU�NAqIRI<�@���oGo�o�o�o��C�p3��O:
��B�+sL�i�O.�PSMT��Y(��@
t�$HOST�C�21��@̹5 MC���R{���  �27.00�1�  e�]�o����� ��K�ď֏���������	anonymous!�O�a�s���"�� �4����� ���D�!�3�E�W�i� ��������ï柀�.� ��/�A�S���课� П����Ŀ���� +�r�O�a�sυϗϺ� ��������'�n� �������ϓ�ڿ���� ������F�#�5�G�Y� k���υ�������� ��B�T�f�C�z�g��� �������������	 -P�����u�� ����(�:�<) p�M_q����� ���/$ZlI/ [/m//�/����/ /�/D!?3?E?W?/ ?�?�?�?�?�/�?./ OO/OAOSO�/�/�/ �/�?�O?�O�O__ +_r?O_a_s_�_�_�O �?O�_�_oo'o�t~�qENT 1�hk� P!�_no  �p\o�o�o�o�o �o�o�o�o:_ "�F�j��� ��%��I��m�0� ��T�f�Ǐ��돮�� ҏ3���,�i�X���P� ��t�՟��៼�
�/� �S��w�:���^��� ���������ܯ=� �QUICC0J��&�!192.168.1.10c��X�1��v�8��\�2��ƿؿ9�!RO�UTER:��!���a��PCJO�G��e�!* �0��U�CAMP3RT�϶�!��߆��RTS���x� �!Softwa�re Opera�tor Pane�lU߇���7kNAM�E !Kj!R�OBO����S_C�FG 1�Ki ��Aut�o-starte�d�DFTP�O a�O�_���O������ ����E_�.�@�R�u� c�	�����������cN :�L�^�;r���R� ������� %H�[m�� �jO|O�O�O4!/h E/W/i/{/�/T�/�/ �/�/�//�//?A?S? e?w?�?����?? �?</O+O=OOO?sO �O�O�O�O�?`O�O_ _'_9_K_�?�?�?�? �O�_�?�_�_�_o#o �OGoYoko}o�o�_4o �o�o�o�of_x_ �_g�o��_��� ��o��-�?�Q�t u��������Ϗ�( :L^`�2��q��� ��������ݟ��� %�H�ʟ[�m������ ����� �ί4�!�h� E�W�i�{���T���ÿ տ�
�Ϟ�/�A�S��e�w����_ERR� ��ڇϗ�PDUSIZ  ��^6����>��W�RD ?(�����  guest���+�=��O�a���SCD_GROUP 3�(�� ,�"�IFT��$PA��OMP�� ��_SHv��ED�� $C���COM��TTP_AUTH 1���� <!iPendanm�x�#�+�!KAREL:q*x���KC��������VISI?ON SET��(� ���?�-�W�R��� v������������������G�CTRL ����a�
�FFF9E3���FRS:DE�FAULT��FANUC We�b Server �
tdG����/�� 2DV��WR�_CONFIG ����������IDL_CP�U_PC� �B����� BH�M�IN����GNR_IO������Ȱ�HMI_EDIT� ���
 ($ /C/��2/k/V/�/z/ �/�/�/�/�/?�/1? ?U?@?y?d?�?�?./ �?�?�?�?OO?OQO <OuO`O�O�O�O�O�O��O�O__;_�NP�T_SIM_DO��*NSTAL�_SCRN� ��\UQTPMODN�TOL�Wl[�RT�YbX�qV�K�EN�B�W�ӭOLN/K 1�����o�%o7oIo[omoo�RM/ASTE��Y%�OSLAVE ���ϮeRAMCA�CHE�o�ROM�O�_CFG�o�S�cU�O'��bCMT_�OP�  "��5sYC�L�ou� _ASG� 1����
  �o������� "�4�F�X�j�|����k�wrNUM����
��bIP�o�gRTR�Y_CN@uQ_�UPD��a��� �bp�b��n��M���аP}T?��k ��._������ɟ ۟퟈S���)�;�M� _�q� �������˯ݯ �~��%�7�I�[�m� �������ǿٿ��� ��!�3�E�W�i�{�
� �ϱ��������ψϚ� /�A�S�e�w߉�߭� ����������+�=� O�a�s���&���� ��������9�K�]� o�����"��������� ������GYk} ��0���� �CUgy�� ,>���	//-/ �Q/c/u/�/�/�/:/ �/�/�/??)?�/�/ _?q?�?�?�?�?H?�? �?OO%O7O�?[OmO O�O�O�ODOVO�O�O _!_3_E_�Oi_{_�_ �_�_�_R_�_�_oo /oAo�_�_wo�o�o�o �o�o`o�o+= O�os����� \n��'�9�K�]� ���������ɏۏi��c�_MEMBER�S 2�:��   $:� ���v���1����RCA_ACC� 2���   [~	�I P�R s�� H� 3�e@l�-l��  �3*�  �������  
l���a�B�UF001 2��n�= �u0�  u0������u0g����u0�l����u0^��u0��-:�D:��p��p�>��=�=��  B�B��^�D=�=U��:��r��r�!���
Z�J_X_�X��fu06�>�Xq����������u0A4 k݊��:�ҤU#Ҥ9ҤPҤgҤ�|:� ���,�C�X��o���������=h=h  �	<sPY�Ȼ	I�	SW�W�0����r��r��r�������*�6�E��Q�`�k�w�ߙ2������x���s�P ��78=�(�q= 0�r��8�J�p\�n�����r���<�±�t� `������u ȯگ�����"�4�F�X�sP V�a��h�j�p��x� }ҁ�}҉�}ґ�� ¡�©�±�¹� ����ɰ�Ѱ�ٰ���ߙ3����� ����!��)�G� 1�>�B�>�J�>�R�>� Z�>�b�l�i�n�r�n� ���n��n�3���� ���⡠��䰣���� �Þ�������l����� ��������������� 
�l�����"�� *��2��:��B�� J��R��Q�l�X�f� a�o�l�p��~򁲏� ~򑲟�⡲��Ⱳ ��������Ѳ�����ݖCFG 2��n� 4��	l�
l�<l�47�a��HIS钜n� ��� 2025�-11-3�l��    #� &��  7 珪�����(7[}�Rq29}	7v���������l�;  ��   % �  � -�RO  *� l��B��aN/`/r/�/�/ �/�/�/�/�/'/9/&? 8?J?\?n?�?�?�?�? �?�/?�?O"O4OFO XOjO|O�O�O�?�?�O �O�O__0_B_T_f_ x_�O�O�O�_�_�_�_ oo,o>oPo�O��([m
8��c���b _o�o�o�o); M;M_���� ����$:�a U2l�d ,l�c 1  \�_�_m� �������Ǐُ��� ��_X�E�W�i�{��� ����ß՟��0��� /�A�S�e�w������� ��������+�=� O�a�s��������� ߿���'�9�K�]πoρ�J�Ѐo�o

 n���������*�<� N�`�r�`r����� ������&�8�&��2��� Z� �־� п����������� �&�8�o��n����� ������������G� Y�FXj|��� ���1�0B Tfx����� 	//,/>/P/b/�t/�/�/�Ϙ�I_C�FG 2��� �H
Cycle� Time�B�usy�Idl��"�min�+�1Up�&��Read�'D�ow8? 2��#Count�	ONum �"����<��b�qaPROmG�"�������)/softp�art/genl�ink?curr�ent=menu�page,1133,1�/OO/OAO�3b5leSDT_ISOLC  ���� �@�.J23�_DSP_ENB�  vK0�@IN�C ��M�ӄ@A�   ?�  =���<#�
�A�I:�o���N_����O<_�GOB�0C�C5�FVQG_GROUP 1�vKw<6�<�P�C�٢_D_?���?�_��Q�_o.o@o�_ dovo�o�o��,_NY�G_IN_AUT�OcT�MPOSRE�^_pVKANJI_�MASK v�HqR�ELMON ��˔?��y_ox������.6r�3��7ĲC���u�o�DKCwL_L�`NUM�@��$KEYLOGOGING�����Q��E�0LANGUA_GE ��~���DEFAUgLT ����LG�!���:2��x��@W�80H  ����'��  � +
��ћ��GOUF� ;��
��(�UT1:\��  �-�?�Q�h�u����������ϟ�����(�g4�8i�N_DISP ��O8�_��_��LOCTOL����Dz`�A�A���GBOOK ����d�1
�
�۠X����#�5�G�Y�`i���3{�W�	��@쉞QQJ¿Կ1���_BUFF 2�NvK ���25�
�ڢVB&�7 C�ollaborativ�=�OΗώ� �ϲ���������'�� 0�]�T�fߓߊߜ��?DCS ��9�B �Ax���Rh�%�-�?�|Q���IO 2���� ���Q� ������������ �*�<�N�b�r����� ����������&�:e�ER_ITMsNd�o����� ��#5GYk }����������hSEV��M.dTYPsN�c/pu/�/
-�aRST5����SCRN_FLW 2�s��0��� �/??1?C?U?g?�/�TPK�sOR"��NGNAM�D��~�N�UPS_ACR� ��4DIGI�8~+)U_LOAD[P�G %�:%T_NOVICEt?���MAXUALR�M2��1���E
LZB�1_P�5�0 ��4y�Z@CY��˭�O�+���ۡ�D|PP 2]�˫ �Uf	R/ _
_C_._g_y_\_�_ �_�_�_�_�_�_oo ?oQo4ouo`o�o|o�o �o�o�o�o)M 8qTf���� ���%��I�,�>� �j�����Ǐُ���� �!���W�B�{�f� ������՟����ܟ� /��S�>�w���l��� ��ѯ��Ư��+���O�a�D���p���RHD�BGDEF ��E�ѱO��_LDX�DISA�0�;c�M�EMO_AP�0E� ?�;
  ױ��3�E�W�i�{ύ���ϱ�Z@FRQ_C_FG ��G۳�A ��@��Ô�<��d%�� ������Bݯ�K���*i�/k� **:tҔ�g�y�ߔ��� �����������J� ���Es�J d������,(H���[���� �@�'�Q�v�]����� ����������*�NPJISC 1��9Z� ������ܿ������	Zl_MSTR �#-~,SCD 1�"��{����� ���//A/,/e/ P/�/t/�/�/�/�/�/ ?�/+??O?:?L?�? p?�?�?�?�?�?�?O 'OOKO6OoOZO�O~O �O�O�O�O�O_�O5_  _Y_D_i_�_z_�_�_ �_�_�_�_o
ooUo @oyodo�o�o�o�o�o �o�o?*cNl�MK���;�љ$MLTAR�M���N��r� ��հ��İM�ETPU��zr���CNDSP_A�DCOL%�ٰ0�C�MNTF� 9�F�Nb�f�7�FSTLqI��x�4 �;�ڎ�s����9�PO�SCF��q�PR�PMe��STD�1ݶ; 4�#�
v��qv�����r��� �����̟ޟ ��� V�8�J���n���¯������9�SING_CHK  ���$MODA����t�{�~2�DEV �	�	MC:>f�HSIZE��zp��2�TASK �%�%$1234?56789 ӿ��0�TRIG 1�; lĵ�2ϻ�0!�bϻ�YP�����H�1�EM_IN�F 1�N�`�)AT&FV0�E0g���)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ��2��H6� ^���Rφ��A�߶� q�������� ��5� �����ߏ�B߳��� ��������1�C�*� g��,��P�b�t��� ���R�?���u 0��������� ������M q�� �Z���/�%/ ��[/ 2�/�/ h�//�/�/�3?�/ W?>?{?�?@/�?d/v/ �/�/O�//OAOx?eO ?�ODO�O�O�O�O_��NITORÀG �?z�   	�EXEC1~s&R2*,X3,X4,X5,X���.V7,X8,X9~s 'R�2�T+R�T7R�TCR �TOR�T[R�TgR�TsR��TR�T�R�S2�X2��X2�X2�X2�X2��X2�X2�X2�X2*h3�X3�X37R2��R_GRP_SVw 1��� (��?-W��
M���⽀t<����#@>be�a���_D�B���cI_ON_DB<��@��zq  �2pt�2puY�1t��p�~>w�  +^p�,Y��@N   ,e�rp�>|$�VY�-ud1������8�PG_JOG� �ʏ�{
�2��:�o�=���?����@0�B��~\�n���������H�?��C�@�pŏ׏���  ������qL_NAM�E !ĵ8���!Defaul�t Person�ality (from FD)qp�0�RMK_ENOgNLY�_�R2�a� 1�L�XL��8�gpl d����şן���� �1�C�U�g�y����� ����ӯ���	���� 
�<�N�`�r�������p��̿޿� :� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w���������������+��<�Se w�������x��A�a��AB�Bw��Pf ������/!/ 3/E/W/i/{/�/�/�/ ���/�/??/?A? S?e?w?�?�?�?�?�? �?�?�/�/+O=OOOaO sO�O�O�O�O�O�O�O __'_9_&O�S��!upz_�[�rdtS�� �_�]�_�_�W�����S�"oe_oXoa  ��qogoyo�o�o�o�o@�ouP�p"|����	`[oUgy8qK��A\����s� AA ��y@h�Q�Q��e"���Tk\$���  ��P��PE�xC�  �I�@oa�<o��p��� ����ߏ
f�Q*������0��PCr� �� 3r �.� �@D�  A�?��G�-�?.I�.@I��A����  ;��	lY�	 ��X  ������� �,? � ������uPK�o������]K��K]�_K	�.��w��r_	����@
��)�b�1�����I��Y�����T;�fY�{S���3����I�>J���;�Î?v�>��=�@�����E��R ѯעZ���wp��u��� D!�3���7pg  �  ��9�͏W���	'�� � u�I�� �  ���u��:�È��ß�=��ͱ���@��ǰ�3��\�"3�E�&���N�pC�  'Y�&�Z�i�bb�@f�i�n�C��D��I�C����b��r���`����B�p�Ŕq���}ر�.DzƏ<ߛ�`�pK�pߖ����������А G4P����.z���d  �Pؠ?�ff�_��	��C 2p>�P���8.f�t�>L���U���	(.��P���������
ĉ��� x��;e��m��KZ;��=g;�4�<�<����%�G���3����p?fff?�ذ?&S���@==0e�?��q�+ �rN�Z���I���G��� 7���(�����!E 0iT����+��F�p���# ��D��w�� �����//=/ (/a/L/�/p/��/� p�6�/Z#?�/ ?Y? k?}?��?�?>?�?�?@�?�?�?1O�����KD�y^KCO�OO�O���ذO�O�O�Oai����J��}�DD1���.�D��@�AmQ�a��9N,ȴA;��^@��T@|�j@$�?��V�>�z�ý���=#�
>�\)?��
=��G�-]�{=����,��C+�?�Bp���P���6��C98R����?N@��(���5-]G��p�Gsb�F��}�G�>.E��VD�Kn����I�� F��W�E��'E����D��;n����I��`E��G��cE�?vmD���-_�o Q_�o�o�o �o$ H3X~i��� ������D�/� h�S���w�������� я
���.��R�=�v� a�s�����П����ߟ ��(�N�9�r�]��� ������ޯɯۯ��� 8�#�\�G���k����� ��ڿſ���"��F� 1�C�|�gϠϋ��ϯϠ��������P(�Q3g4�] �����Q��	�9�Oߵ53~�m8m��aҀ5Q�߫ߎaғ����ߵ1�������1��U�PC�y�g��%P�P���!�/��'���
���<.������4�;� t�_������������� ��:%��/�/d������ ��7%[I m���027��  B�S@J@�C%H#PzS@�0@ZO/�1/C/U/g/y/�-�#���/�/�/�/�/�3?Y�3�� @�3�%�0�0�13��5
 ?f?x?�? �?�?�?�?�?�?OO�,O>OPO�Z@1 ����ۯ�c/�$M�R_CABLE �2ƕ� ��TT�����ڰO�� �O�)�@���C_��� _O_u_7_I__�_�_ �_�_�_o�_�_oKo qo3oEo{o�o�o�o�o �o�o�o�oGm/�K!�"���O�����ذ�$�6����*Y�** �CO�M ȖI�����"P�'%%� 2345678'901���� ��Ï���� � !� �!
���Mn�ot sent �b��W��T�ESTFECSALGR  eg�*"!d[�41�
k�������$pB����������� 9UD�1:\maint�enances.�xmlğ�  �C:�DEFA�ULT�,�BGRP� 2�z�  ��14��%  �%!�1st clea�ning of cont. v��ilation +56��ڧ�!0�����+B��*������+��"%��me�ch��cal c�heck1�  ��k�0u�|�� ԯ����Ϳ߿�@���?rollerS�e�w�ū��m�ϑϣ����@�Basic� quarterCly�*�<�ƪ,\��)�;�M�_�q�8�MXJ��ߓ "8��� ���ߕ �����+�=��C�g�ߋ���߹���������@�Overha�u�ߔ��?� x� I�P����}���������� $n���� ���)l�ASew� ����� � +=O�s��� ����/R�9/ �(/��/�/�/�/�/ /�/�/N/#?r/G?Y? k?}?�?�/�???�? 8?OO1OCOUO�?yO �?�?�O�?�O�O�O	_ _jO?_�O�Ou_�O�_ �_�_�_�_0_oT_f_ ;o�__oqo�o�o�o�_ �oo,oPo%7I [m�o��o�o� ���!�3��W�� ������ÏՏ�6� ���l����e�w��� ������џ�2��V� +�=�O�a�s���� ��ͯ����'�9� ��]�������⯷�ɿ ۿ���N�#�r���Y� ��}Ϗϡϳ������ 8�J��n�C�U�g�y� ���ϯ������4�	� �-�?�Q��u����� �ߞ���������f� ;������������ �����P���t�I [m����� �:!3EW� {��� ��� //lA/��w/���/�/�/�/�/X*�"	� X�/?.?@?�)B a/o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�_�_�_�_�_	o�o" Џ!?� ; @�! M?Ho Zolo�&4o�o�o�o�(�*�o** F�@ i!k&�`o�'9�o]o�����/^&�o��� ��/�A�S�e��� #�����я����� +�q�����7������� k�͟ߟ��I�[��� K�]�o���C�����ɯ���o$�!�$M�R_HIST 2��g%#�� 
 �\7"$ 2345?6789013�;���b2�90/���� [���./����ǿٿ F�X�j�!�3ρϲ��� {��ϟ�����B��� f�x�/ߜ�S����߉� �߭��,���P��t����=��$�SKCFMAP  g%�&��b
�� ����ONREL  �$#�������EXCFENB��
����&�FNC�-��JOGOVL�IM�d#�v���K�EY�y���_�PAN������R�UNi�y���SFSPDTYPM�<���SIGN���T1MOTk�����_CE_GRP7 1�g%��+� 0�ow�#d�� ����&�6 \�7y�m� ��/�4/F/-/j/ !/t/�/�/�/{/�/�/�/?�+��QZ_E�DIT
����TC�OM_CFG 1����0�}?�?�? }
^1SI �NB����?�?���?�$O����?XO78T__ARC_*��X�T_MN_MO�DE
�U:_S�PL{O;�UAP_�CPL�O<�NOCHECK ?��/ �� _#_ 5_G_Y_k_}_�_�_�_��_�_�_�_oo��N�O_WAIT_L�	S7> NTf1�����%��qa_ERMRH2������� ?o�o�o�o��O�Gj�@O�cӦm| �P�^GA5�E��@�������7P}��D�;/����<���?���)��n�b_PARAM�b����vHO��w
�.�@� = n�]�o� w�Q�����������`Ϗ�)���w�[��m� �����ODRD�SP�C8�OFFSET_CARI0��OǖDISԟœS;_A�@ARK
T9�OPEN_FIL�E��1T6�0OPTION_IO�����K�M_PRG ;%��%$*�����'�WO��N�s�ǥ�� ���u����	� ����Ӧ������RG_DSBL'  ����jN����RIENTTO����C�����A� ��U�@IM_D�S���r��V��LCT �{mP2ڢȪ3̹��dҩ��_P�EX�@���RAT��G d8��̐UOP װ�:�����S�e�Kωϗ��$��r2G�L�X�LȚ�l 㰂�������'�9� K�]�o߁ߓߥ߷��� �������#�5�G���2��v������� ������e�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?�q1�~?�?�?�? �?�?�?�?O O2ODO^�yA�a�m? ~N��~O�O�P�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�O �Oo$o6oHoZolo~o �o�o�o�o�o�o�o  �_oVhz�� �����
��.��@�R�d�QOES��(����B�d�ӏ� ʏ��������Y�D�}�0��r������� ��ԟڟ���p���=�4M��q�	`����x����c�:�o��¯ԯ����A�C  �k�C�C�ڰe"ڰ���O���  ����-���)�C�  �t�k���g�����Կ ��ѿ
�5���_:�ĳ��OU���/��/�H��n��� � ^��\� @D�  &p�?�v�\�?:px��:qC4r�p�(�� � ;�	l��	 ��X � ������ ��, � �x������Hʪ�������H���Hw�zH����ϝ�8�B���B��  Xѐ�`�o�*��'3����t�>u����fC{ߍ��:pB\��
�Ѵ9:qK�t�� �����$���*��� D�P�^��b�g  �  �h������)�	'� �� ��I� ��  ��'�=��������t�@����!�b��^;bt�U�(�N��r� ' '��E�C�И�t�C�И��ߗ���jA��@�����%�B �� ��,���H:qDz�k�ߏz����������А 4P���:uz:���	�f��?�faf'�&8� ]��m�8:p��>!L�����$�(:p�P��	������:�� x�;e�m�"�KZ;�=g�;�4�<<�0��E/Tv��b����?fff?�?y&� )�@=0�%?��%_9��}! ��$�x��/v��/f'�� W,??P?;?t?_?�? �?�?�?�?�?O�?(O OLO�/�/�/EO�OAO �O�O�O�O_�O_H_ 3_l_W_�_{_�_�_1� �_A���eO+o�ORoo Oo�o�o�oK/�o�omo �o*'`+�,�zt���CL�H<��}?����X�
������u�����D1�/n�t�x�p�q��@I�h~�,ȴA;�^@���T@|j@�$�?�V�n��z�ý��=�#�
>\)?��
=�G�����{=��,���C+��B�p����6���C98R����?}p��(��5���G�p�G�sb�F�}�G��>.E�VD��KL����I��� F�W�E���'E���D���;L����I���`E�G���cE�vmD���\�՟��ҟ� ��/��S�>�w�b��� ����ѯ������� =�(�:�s�^������� ��߿ʿ�� �9�$� ]�Hρ�lϥϐϢ��� ������#��G�2�W� }�hߡߌ��߰����� ���
�C�.�g�R�� v��������	��� -��Q�<�u�`�r��� ����������'�M�(�34�]O!���8h~�%3~�m���ǀ5Q��������!���   `N�r��J	eP@"P��Q�_�/V/9/$/]/H)����c/j/�/�/�/ �/�/�/�/!??E?0? i?T?"&�_�_�?�?�8��?�?O�?OBO 0OfOTO�OxO�O�O�O��O2f?_  B���pyp$QCHR�z�p@�N_`_r_�_�_�_�]c�O�_�_0oo+o?�Bc�� @d4��QJc�D
 2o�o�o�o�o�o�o %7I[m���oa ������c/�$PARA�M_MENU ?� � � DEF�PULSE��	�WAITTMOU�T�{RCV� �SHELL_�WRK.$CUR�_STYL�p�"�OPT8Q8�PT�BM�G�C�R_DECSN�p����� ���������-�(� :�L�u�p��������q�SSREL_ID�  ��̕U�SE_PROG �%�z%���͓C�CR�pޒ��s1�_HOST !�z#!6�s�+�T�=����V�h���˯*�_�TIME�rޖF�~�pGDEBUGܐ��{͓GINP_F�LMSK��#�TR\2�#�PGAP� ���_b�CH1�"�TWYPE�|�P�� ������0�Y�T� f�xϡϜϮ������� ���1�,�>�P�y�t� �ߘ��߼�����	�� �(�Q�L�^�p��%�WORD ?	�{
 	PR��p#MAI��q"3SUd���TE��p#��	1���COL�n%��!���L�� �!��F�d�T�RACECTL �1� �q }�� �#�����_�DT Q�� ��z�D �� �� ��M`��k`�������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEO_@� ROLO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �[��rEoo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�.�oP�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/Dϒ/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D��V�h�z�����������$PGTRACE�LEN  �� � ������Ά_UP _�����������΁_CFoG ����*��
���*�*�D��O���O�  ��O��DEFSPD� ��������΀H_CONF�IG ����� ����dĔ�&݂ ��ǑP^�a�l㑹��΀IN�?TRL ��=��8^���PE��������*�ÑO��΀LID���	~T�LLB 1ⳙ_ ��BӐsB4��O� �𼧶��Q� <<7 ��?��� ����M�3�U���i� ��������ӿ��	�7�T�Ϣk�b�tϡπ诚��������S�G�RP 1爬����@A!���4�I���A �C�u�C�OCWjVF�/��Ȕ`a�zي�ÑÐ�t�0�ޯs���´�ӿ���B������������A�S�&�B3�4�_������j���������	� B�-���Q���M�������  Dz����.� ����&L7p[ ��������6!Zh)w�
V7.10be�ta1*�Ɛ@��*�@�) @ߺ+A Ē?���
?fff>�����B33�A�Q�0�B(���A���AK��h����//('/9/P�p*�W�ӑ��n/�/�%���R��fh���� *���P2�LR��/�/@�/�/�/H?�Ĕ�I�u�&:���?��x?��?A���P!\3 Bfu�B��?�5BH�3�[4��o��4�I�[45��/B\3x3Dx�?YO�?aOkO}O�<<�R@��O�C�O�O��O�O�DA�X�KNO?W_M  Z�%��X�SV 賚ڒ���_�_�_?��_�_�_o����W�M�+�鳛 ��	~<�3#���_��o�\=��
]bV4�@u��u��e��o�l,�X�MR+��JmT3?��W�1C{��OADBANFW�DL_V�ST+�1 k1����P4C� ��[��i/��� ��?�1�C���g�y� �������ӏ�*�	�@�`�?�Q�c��w2�|8Va�up�<ʟ����p3��Ɵ؟Ꟃw4 ��+�=��w5Z�l�~����w6����ѯ㯂�w7 ��$�6��w8`S�e�w����wMAmp�������OVL/D  ��yo���rPARNUM � �{+þ�?υqS[CH�� �
��pX���{s��UPDX��)ź��Ϧ�_CMPa_@`���p|P'yu~�ER_CHK���yqbb3��.��RSpp?Q_MO�m��_}ߥ�_REWS_G�p쩻
� e�����0�#�T�G�x� k�}��������������׳�������� �:�Y�^���Y�y��� ���Ӭ����������� ����R�6UZ��ӥ�u����V �1�FvpVa@k��p��THR_ICNRp��(byudoMASS Z)�MNGMON_�QUEUE �P�uyvup\!��N��UZ�NW��ENqD��߶EXE�����BE���O�PTIO��ۚP�ROGRAM %z%��~Ϙ?TASK_I��.OCFG �zx+�n/� DATACcm�+�0�)up 2 �? ?/?A?S?]51q?�? �?�?�?�8p?�?�?OxO,J�!INFOCc��-��bdlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_��_�_�/A@FD��, �	��!��K_�!q�)fN!fENB��H0m��Pf2YokhG�!�2�0k X,{		d�=��·o���e�a$�pd��i��i�g_EDIT� ��/%7�����*SYSTEM�*upV9.401�07 cr7/23�/2021 A���Pw��PR�GADJ_p  �h $X[�p� $Y�xZ�xW��xқtZқtSPE�ED_�p�p$N�EXT_CYCL�E�p���q�F�G�p ��pA_LGO_V �p�NYQ_FREQ��WIN_TYP��q)�SIZ1�O�LAP�r!�[���M+����qCREA�TED�r�IFY��r@!NAM�p%�h�_GJ�STAT�U��J�DEBUG~�rMAILTI�����EVEU��L�AST�����tEL�EM� � �$ENAB�rN�E�ASI򁼁AXIS�p$P߄������qROT_RA" �rMAX ��q�E��LC�AB
�<��C D_LVՁ`�BAS��`�1�{���9_� ��$x����RM� RB�;�DIyS����X_SPo��΁�� �u�P�� | 	� 2� \�AN�� �;�����Ӓ��� �0�PAY�LO��3�V�_DO�U�qS���p�tPR�EF� ( _$GRID�E
����R���Y� � �pOTOƀ�qO  �p��!�pܫ�k�OXY� ߤ $L��_P�O|�נVa�SR�V��)���DIR�ECT_1� �2�(�3(�4(�5(�6J(�7(�8��qF���A�� $VA�Lu�GROUP������F��� !��@!��8�����RAN泲�⚁R��/���TOTaA��F��PW��I=!%�REGEN #�8�������/��фڶnTzЉ���#�_!S����8�(�V[�'�8��4���GRE��w����H��D�����V_]H��DAY3�V���S_Y�Œ;�SU�MMAR��2 �$CONFIG�_SEȃ���ʅ_�RUN�m�C�С�$�CMPR��P�D�EV���_�I��ZP�*Ӥ���ENH�ANCE�	�
����1���INT���qM)b�q�2Kܖ���OVRo�PG�u�IX��;���OV�CT�����v�
 4� ����a˟��P�SLG"�� \ �;��?�1���qSƁϕc�U� ����Ò�4�U�q]�|Tp� (`�T-��rJ<�O� CK�OIL_MJ���VN�L+��TQn{�N5����C�ULȀD�V(�C6�P_�຀@�mMW�V1V�V1d�U2s�2d�3s�3d�4s�4d��'�	��������p	�IN	VGIB1qp1� 2!�pq/,3 3,4 4,�p?��;���A���N�������PL��TORr3�	���[�SAV���d�MC_F�OLD 	$CSL�����M,�1I��L� �pL��b��KEEP_H/NADD	!Ke��UCCOMc�`k��
�lOP����pl��lREM�k��΢����U��ekHPWv� KSBM��~ŠCOLLAB|��Ӱn��n�+�ITz�O��$NOL��FCALX� �DO�N�r���� �,��FL���$�SYNy,M�C�=����UP_DL�Y�qs"DELAh� ����Y(�AD���$TABTP_�R�#��QSKI�Pj% ����OaR� �E�� P_�� � �)���p7��%9 ��%9A�$:N�$:[�$:@h�$:u�$:��$:9�q��RA�� X������MB�NFGLIC]��0"�U!�<o���NO_H� ��\�< _SWITC�Hk�RA_PAR�AMG� �4�p��U��WJ��:C|ӣ�NGRLT� OO�U�����X�<A���T_Ja1F�rAP�S�WEIGH]�Jg4CH�aDOR��aD��OO��)�2�_FJװ���sA�AV��C��HOB.�.�l�J2��0�q$�EX��T$�'QIT��'Q�pGp'Q-�G��RDC�>m" � ��<���
R]��
H���R�GEA��4��U�F�LG`g��H��ER�	�SPC6R�rU�M_'P��2TH2�No��@Q 1� @ED���� ? D �وI�i�2_P�25cS��ᰁ+�L10_C�I��pe�  �pk����UՖD�� zaxT�p�Q(�;a ��c��޲+�i���eܶ�` P`DE�SIGRb$�VL1b:i1Gf�c�g10��_DS��D��w�P�OS11�q l��pr��x1C/#AT��B��U
WusIND��}�mqCp�mq�`B	�HOME�r )	aBq2GrM_@q����!@s3Gr��� ��$�`!
@s4GrG�Y�k�}�(����6�5Grď֏��������6Gr�A�S�e�w�����6�7Gr��П�����
��8Gr;�M�_�q�ȃ�����S �q    �@sM��P�!x�K@��! T`�M��M�IO��m�It��2�OK _OPy�� »Q6�POWE" 7�x EQu�1E � #s%�Ȳ$DSBo�GNA�b� C�P2�B�S232S�$ ��iP��xc�ICE�<@%�PE`2� @I9T��P�OPB7 1�oFLOW�TRa@42��U$�CUN��`��AUXT��2Ѷ�EORFAC3İUU���CH��% �t<_9�EЎA�$FREEFRO	MЦ�A�PX q��UPD"YbA�PT�.�pEEX0����!��FA%b�/��R�V�aG� & � ��E�" 1�AEL�  �+�jc'���D�  2& ��S\PcP(
  �	$7P�%�R�2� ���T�`AXU���DSP���@�W���:`$���RNP�%�@����K��_MIR�����3MT��AP��0�P"�qD�QSYz������QPG7�BRKqH���ƅ AXI�  ^��i���1x ����BSOC����N��DUMMY{16�1$SV��DE��I�FSPD/_OVR79� �D����OR��֠N�"`��F_����@OVv��SF�RUN�b�"F0�����UF"@vG�TOd�LCH�">�%RECOV��9@�@W�`&�ӂH��r:`_0��  @�R�TINVE��8AO�FS��CK�KbFWD������1B���TR�a�B �FD�� ��1= B1pB�L� �6� A1L�V ��Kb����#��@+<�AM:��0��j���_M@ ~�@h����T$X`x ��T$HBK���F��A�q����PPA�
���	������DVC_DB�3@pA �A"��X1`�X3`��S�@�`�0���Uꣳ�h�CAB PP
R�S #��c�B��@���GUBCPU�"��S�P�`R���11)ARŲ�!$HW_CGpl�11� �F&A1Ԡ@8p�$/UNITr�l e ATTRIr@y"��gCYC5B�CA���FLTR_2_�FI������2bP���CHK_��SCmT��F_e'F_o,��"�*FS�Jj"CHA�Q�'91Is�82RSD����1���_Tg�`� i�SEM�NPMf�T&2� 8p&2- �6DI�AGpERAILAiCNTBMw�LO@4�Q��7��PS��梱 � ��PRBS�Z`�`BC4&�	���FUN5s��RIN�PZaߠ�07Dh�#RAH@���`� `C�@�`C�Q�CBL'CURuH�DA�K�!�H�HDAp�aA�H�C�ELD������C��2jA�1�CTIBU�u�8p$CE_R�IA�QJ�AF Pb��>S�`DUT2�01C��};OI0DF_LC�H���k��LMLF�aHRD�YO���RG�@H�Z0��ߠ�@�UMUL�SE�P�'3iB�$J��J����F?AN_ALM�db�WRNeHARDH��ƽ�P��k@2a�N�r�J�_}�AU�J R+4�TO_SBR��~b�Іje 6|?A�cMPINF���{!�d�A�cREGF�NV��ɣZ�D���NFLW%6r$�M�@� ��f� �0l h'uCM4NF�!�ON	 e!e#�(b8*r3F�3 �	 ����q)5�$�$Y�r��Zu�_��p�*$ �/�EG0E�����qAR��i�«�2�3�u�@<�AX�E��ROB��REMD��WR��c�_����SY`��q� ?�S�I�WRI���vE SATհ�ӭ d���Eg!���t8��^a��Bȉ���9�3� OT�O�a���ARY���ǂ�1����FI�E���$LINK��QGTH��Ti_������30���XYZ���!*�'OFF�����%ˀB��,Bl������m�FI� ��C@hIû�,B��_J$��F�����S`����3-!$1�w0���R���C��,�DU���3\�P�3TUR`XS�.�Ձ�bXX�� ݗFL�d���pL�0����34���� 1)J�K��M�5�5p%B'��ORQ�6@��fC㘴��0B�O;��D�,������a�OVE��rM�����s 2��s2��r1���0���0�g /�AN=!�2� DQ�q���q�}R�*���6����s��V���E)R��jA	�2E��.�$C��A���0��XE`�2Ӈ�A��AAX�� F��A�N!�SŴ1_� �Q_Ɇ�^ʬ�^ʴ�^�@�0^ʙ�^ʷ�^�1&� ^ƒP[ɒPkɒP{ɒP �ɒP�ɒP�ɒP�ɒP �ɒP�����ɪ �R>�oDEBU=#$8A`Dc�2����
�AB�7�����V� <" 
��i�q��-!��%� �׆��׬��״����1 �י��׷�JT��DR�.m�LAB��ݥ9 �FGRO� ݒ=l� B_�1�u���}���`����ޥ��qa��AND�����qa� �Eq��1��A@�� �NT$`��c�VEL�1��m��1u�0��QP��m�NA[w�(�CN1� ��3줙��  �SERVEc�p+ $@@d@��7!��PO
�� u_�0T !������p,  ]$TRQ�b
d(� -DR2,+�"P�0_ . l8"@!�&ERR��"�I� q���~TOQ����L�p]�e���0eG��%������RE�@ / ,h��/I -��RA�? 2. d�&u��_! 0�p�$&��2tPM��O�C�A8 1  >pCOUNT�� ���FZN_CFG�2 4B �f�"T��:#��Ӝ� x� `�s3 ���M:0�R�qC@��/�:0��FA1P��?V�X������r���� �P:b��HEL�pe4 5���B_BAS�cRSSR�f @�S�!�QY 1�Y 2|*3�|*4|*5|*6|*72|*8�L!RO������NL�q �AB����0Z ACK��I-NT_uUS`�Pta9_PU�>b%ROU��PH@�h9#��u`w�9�TPFWD�_KAR��ar R�E���PP��A]@QUE�i&��	�f�>`QaI`��9#�j3r��f�SEME��6��PA�STY4SO�0�DI'1�`���18�rQ_TM�cM�ANRQXF�EN�D�$KEYSWITCHj31:A��4HE	�BEATmM�3PE�pLE�(�1��HU~3F�42�S?DDO_HOM�BPO:a0EF��PARr��*�v�uC�@�O�Qo �OV_Mtϒ��Eq�OCM��d�7��p8%HK�qG5 D��g�Uj��2M�p�4R��FO;RC�cWAR��NY�OM�p 6 @��Ԣ�v`U|�P�p1(�V'p�T3�V4��OR*#O�0L�R7��hOUNLOE0hd�EDVa  �S�@d8 <pAQ9�}l1MSUPG��UaCALC_PLkANcc1��AYS1�1:b�9 � 	X`��P �q;a@�թ�w��2��j�M$P��㣒�fyt$��rSC�M�pm�q ���aq���0�tYzZzE!U�Q�b�� T!�Hr��pPv	NPX_A�Sf: 0g AD�D��$SIZ�%a$VA��M_ULTIP�"ns��PA�Q; � �$T9op�B���rS��j!C~ �vFRI	F�2S�0�YT�p{NF[DODBUX�`B��u&�!���CMtA�Е����������+Z ��< � ��p�TEg�����$�SGL��T��X�&�{���㰀��STMyTe�ЃPSEG�2���BW���SHO�W؅�1BAN�`TPO���gᣥ�����ѵ��V�_G�= ��$PC����O�FB�QP\�SPb�0A&0^�� VDG�~�>� �cA00�����P���P����P���P��5��6���7��8��9��A ��b`���P��w᧖��B��F����h���1���v�h�י1�1�1���1�1�1%�1�2�1?�1L�1Y�1�f�2��2��2��2�ʙ2י2�2�2���2�2�2%�2�2�2?�2L�2Y�2�f�3��3��3��3*ʙ3י3�3���T��3�3%�32�U3߹3L�3Y�3f�U4��4��4��4ʙU4י4�4�4��U4�4�4%�42�U4߹4L�4Y�4f�U5��5��5��5ʙU5י5�5�5��U5�5�5%�52�U5߹5L�5Y�5f�U6��6��6��6ʙU6י6��6�6��U6�6(�6%�62�U6߹6L�6Y�6f�U7��7��7��7ʙU7י7��7�7��U7�7(�7%�72�U7߹7L�7Y�7f�z[V�`_UPD���? �c 
�ZB����@ x �$TOR�1T� � �cOP �, ZQ_7RE^��� J�J�SsC�A���_U�p��YSL}OA"A � �u $�v��w�@���@��bVALUv10�6��F�ID_L�[C:HI5I�R$FILE_X3eu4�$�C7 �SAVΔ�B hM �E_BLCK�3�ȁ�D_CPU��p���p5hz��@S2R� C � PaW��� 	�!LAށ�SR�#.!'$RUN�`G@%$D!'$@�@G%e!$e!'%HR0�3$� '$7aT2Pa_�LI�RD  �� G_O�2�0P�_EDI�R�"SPD�#E�"i0ȁ��p�Q�DCS9@G�)F � 
$GJPC71��� S:�C;C9$MD�L7$5P>9TCL�`@7UF�@?8S� N?8COBu �@�"T|�L�G�P;;԰ 9:;�qTAOBUI_�!L�HGb��% FB3�G$�3A�sR�LL?B_AVAI�B����3�!��I $� S�EL� NẼ�@R�G_D N��Ta����4SC�PJ )�1/AB�PT�R?��w@_M]`L�K \�M f/QL_��FM�j��PGi�U9R�6���PS_�P\� ��p�EE7B�TBC2�eL ���``�`6b$�!FT�P8'T�`TDCg�� `BPLp�sNU;WTH���qhTgtWR�2=$�pERVE.S�Tp;S�Tw�R_ACkP� MX -$ �Q�`.S�T;S�PU@�`�IC�`LOW�GF	1�QR2g�`��p|�S�ERTIA�d`^0iP�PEkDEUe��LACEMzC	C#c�V�BrpTf�edg�aTCV�l�adgTRQ�l�e�j|�Scu��edcu�J7_ 4"J!��Se@qde�Q2�0���1�PRc6uPJKlvVK<�~qcQ~qw�spJ0��q�s�JJ�sJJ�sAAL�s�p�s�p�v���r5sS�`N1�l�p�k�`5dXA_́� P�CF�BN `M G�ROU ��bh�N�PC0sD�REQUsIR�R� EBU�C��Q�6g0 2M�z��Pd�QSGUOz�@�)APPR0YC7@� 
$� N��'CLO� ǉS^U܉�Se>@BC�@A�"P �$PM]P�`�`sRN�_MGa!�C����+��0�@,�BRK�*�NOLD*�SHORTMO�!m�Z��JWA�SP�tp`�s p`�sp`�sp`�sp`�Aꪒ7��8sQIR_|�RTQ� m���R.Q�cQ�PATH�*� �*��X&����P�NT|@A��"p��� �IN�RU�C4`a��C�`UM��Y
`�)p��>��Q��cP���p��PA�YLOAh�J2LN& R_Am@�L ������+�R_F�2LSHR�T/�L�O���0���>���ACRL0z�p�y�ޤsR9H5b$H+����FLEX��#�JVR P��_._�_�_QJ�US :�_�Vd`0�G��_`tQd`�_�_lF1G� �ũ�o0oBoTofoxo��E�o�o�o�o�o�o �o ����wz3lt�����3EWF�^zT!��X���ju�� uu~�W؁���p�u��u�u�u����U9M��(�T �P5�0G�Y�' AT��l��pEL0�_B��s�J��Sz�JEW�CT�R7B`NA��d�H�AND_VB��(��TUO@`+�`TSW8F�A�V� $$M� �e G�AV�Qs�De�oAA��@�	�$�A5�G�AU�A�d�� 6��G�DU�D�d�PD�G/ -ST�I�5V�5Ng�DY F ��+�x����P&� G�&�A��lw�o�Q�k�P������ʕӕܕ���DX�TW1 7 �� ��3%<�?!ASYMT�(�	m�T�V*�o�A�t�_SH�~������$@����Ưد�J�����#39"���_V�I��`8�q0V_�UNIrS�4��.�J mu�2��2A��4X��4 �6a�pt�������&E�_�����RE��C�H( X �̱���TOc�PPB�VsSvD�US�RU�P�����z@�D�A}@_5�U��P�EyAa��RPROG_NA���$�$LAST���CANs�ISz@?XYZ_SPu�D W]R@Ͱ,VSV@�E�1QENc��DCURx�H#���HR_T��#YtQ9S�d�z�O�T 
Z�tQN?�Z ��I�!A�D���Q���#�S���� �3�vP [ �� ME��O��R#B�!T�PPT@0F@1�a-�1�̰�� h1a%iT0�� $DUMMY}1��$PS_���RF��!�$lfnװFLA*�YP���bc$GLB_�TI �U�e`ձ��L;IF(!\�����g`OW�P��eVOeL#qb �a_2��[d2�[`����b�P��cZ`TC��$BgAUDv��cST���B�2g`ARITY�0sD_WAItAI�yCJ2�OU6�|ZqyyTLANS�`̌{S�SZc��BUF_�r�fиx�Pyy�CHK_�@CESZ��� JO`E�a�A�x�bUBYT �����r�.�.� � �aA��M�������Q] Xʰ����SuT����SBR@�M21_@��T$SV_ER�b����SCL�`��A1�O�B�pPGLh0EW(!^� 4 $a$vUq$�q$W��9�A�@R���u�ӃUم_ "���D$GI��}=$ف ^���(!` L�.��"}�$F�"E6�NEA9R��B$F}��QTQL���J�@R�� amP$JO�INTa�)�&ՁMwSET(!b  +�QEc�2�^�ST��H�|_�(!c�  ���U�?���LOC�K_FO@� �PB�GLV��GL'�T�E�@XM���EM�P����K��b�c$U�؂a�2_����q�`<� �q�^ƒ�CE/�?��� $�KARb�M�STP�DRA܀����VE�CX�����IUq�a�v�HE�TOOL����V��REǠI�S3��6��ACiH̐m b^QONe�[d3���IdB�`@�$RAIL_BO�XEa���ROB��@D�?���HOW�WAR0Aa�i`-�ROLMtb��$�*���pT��`����O_FU��!��HTML5 8QS�� e�"Հ�(!d����@�(!!e������І}pN(!f t��m�^a���t��B�PO��AIPE�N���O�����q��AORD�ED�m �z�XT�`��A) ��P�O��P g D �`OB�����ǯ��Uc�`��� ��SYS��ADR��pP`U@>^  h ,"��f'$A��E��E�тVWVA�Qi� � �@ق�UP�R�B�$EDI|�Ad�VSHWRU�z���IS�Uq�p�ND�P7���G�HECAD�! @���!i�3KEUqO`CP)P���JMP��L�U��TRACE�Tj����IL�S��C���NE���TI�CK!M4�_�N��HNr�k Q@���HWC��P�F�F��`STYeB+�L�O�a9�' ��[�C�l23�
�@�F%$A��Du=��S�!$�1 �p a�e�q�ePv �FgSQU��#LO�b_1TERC`!oP=S?�m 5���@R�m@3���ܡ�O`�	c IZ�d�A�e@ha�qtb}�hA}pP~rN��_DO�B�X�p9SSQ�SAXI�q��!v�bS�U�@TL��ƞREQ_ܠ��ET���`�CY%�P��Z&���Af\!\d9lx�P MBSR$$nl-�w ��� ��c
�uV
Qh(�A���dC`�A��	�Y��AD��p�E"�	CC��C��/�/�/	4�ISC�` o �h��DSmడ[`S�P�@�AT� 
R���L��XbADDRf�s$Hp� IF�C�h�_2CH���pO�����- �TUk�Inr p�CUCpT�V��I�Rq�P4���c��
K�
��8^ ���Pr \z�D�A���|,K� P�"C�N��*CƮ��!�T�XSCREE��s8�Pp@�INA˃<��4�D������`t Tᫀ�b����O �Y6���º�U4h�RR��������R1�T � �UE��u ��j �qz`Ś��RS	ML��U����V�1tPS_��6\��1�9�G\���C��2@4 c2��0Ov�R���&F�AMTN_FL*�`Q��W� ��/BBL_/�WB`�P�w ����BO ��BLE"�Cg�R"�DoRIGHtRD���!CKGRB`�ET����G�AWIDTH�s���RB��a�r��UI��EYհRx� d�ʰ�����`y�BACK��tb>U����PFO��QWL[AB�?(�PI��$URm�~P��P�PHy1 y o8 $�PT_��,"�R�PRUp�s5�Hda���QO%!t�zV�Iȇ�pU�@�SR ����LUM�S�� E�RVJ��SP��T{o � " GE�R0h� �¯�LPAe	E��)^g�lh��lh�ki5ik6ik7 ikpP`�Z�x����$�u1��p�Q �zQUSRل| <z��PU2�a#2�sFOO 2�PRI*�m9�[�@pTRIP�K�m�UNDO��})���Yp���y����h����p �~�Rp�qG ¸�T���-!�rOS2��vR��2�s�CAA�����ro���Pi�UIaCA����38Ibn�sOFFA�D@����Ob�r����L�t��GU��P�s��������+QSU�Bo� ��E_E�XE��VeуsWO.� �#��w��WAl�p΁fP
 V_DB���pT�pO�V░����3OR/�5�RAUD@6�TK���__О��� |j �O�WNj�34$SRC�0`���DA���_�MPFI����ESP��T�$0��c���g�Y�q�z�E!� �`%�ۂ34J���C�OP��$���p_����/�+�6���CT��Cہ�ہ�D ��DCS��P�4�COMp�@�;��Oo�=��b�K�^�/�VT�qU'���Y٤Z���2���@p�w#SB�����2�\0˰_��M8��%!]�DIC#��sAY�3G�PEE�@T�QS�VR1���eQL�� a��P�D  ��f�z��f�> ����6�FP�A�t�b# ��L2SHADOW���#ʱ_UNSC�Ad�׳OWD�˰D�GDE#LEGAyC)�q'�VC\ }C��� v����だm�RF07����7d`C2`7�DRI%Vo���ϠC�A]��(�` ���MY_UBY�d?Ĳ��s��1@��$0�����_ఴ����L��BM�A�$�DEY	�EXXp@C�/�MU��X���,��0US��.�;p_�R"1�0p#�2�G>PACIN*���RG��c�y�:�y��sy�C/�RE�R"!�q✂�y�D@� L !�G�P�"�г��R�pD@�&P�Px1dQ��	.���RE���SWq�_Ar��$+�{�Oq�AA/�3��hEZ�U���� YP�HK���P�J��_/�Q0{�EAN��ۀ2�2��P��MRCVCA� ��:`ORG��Q�dR	p��L�����REFoG �����!�+`	�p ��������<���q�A_����r��� S�`�C��Ú�G�@D� ��0�!��#q�š��OU����?� ��Վ2�J@0� 1�*p����0� UL�@��C�O�0)��� NT�[��Z�Qf�af% L飏��Q|��a�VIAچ7� ��@HD7 6P�$JO�`oB?�$Z_UPo��2Z_LOW��$�QiBn��1$EP �s�y�� 1!f� m� 1¦4�� 5�PA�A ��CACH&�LO �w�ВQB����Cn�I#F^��T8m����$HO2�32!{��Uÿ2O�@����Ro��=a��ƐV�P��X@A"_SIZ&�K$Z$�F(�G'��v�CMPk*FAIo�5G��AD�)/��MRE���"P'GP��0е�9�ASYNwBUFǧRTD�%��$P!�COLE_2D_4�5W�sw�~��UӍQO��%EC;CU��VEM��v<]2�VIRC�!5�#�2�!_>�*&�pWp���AG	9R�XYZ@�3�W���8���4+Qz0T"��IM�16�2P�GRA�BB�q��;�LERrD�C ;�F_D��F�f50MH�PE�R9�[��� ��KQ�LAS�@��[_GEb� �H൑~23�ET����"���b¨�I�D�ҙ6m�BG�_LEVnQ{�PK�|Л6\q��GI�@N\P4�n��A��!gI�dr�S� �NRTO�VLʁc�Ų���#a��c"!D�qDE����Xа�X������1��d��p�zZ���d�c���DR4qȲ�2pT��U&��� $�ITPr�9p[Q��ՓV�VSF$�d�  fp/�ff�UR&ҿ�SMZus�dr��ADJ`�C�� ZDVf� D�XAL� � 4 �PERIKB$MoSG_Q3$Q! o%[���p'��dr:g�qQ� �XVR2\t��B�pT_\��R���ZABC"�����Sr���
W��aA�CTVS' � � $|u�0�c�CTIV�Q!IO0u¥s&D�IT�x�DVϐ
x�P��i�!���pPS���� �#��!���q!LSTD�!�  �_ST���aq�;CHx�� L-�@���u�Ɛ*���P G�NA#�C�!q�_�FUN�� uqI�Pu��HR�$L���XZMPCF"��`bƀ�rX�فn��LNK��
Ł��0#�� $x !��ބCMCMk�EC8�C"����P{q? $J8�2�D6!>�O�H���T���`2�����M���UX�1݅UXE1Ѡ��1C� ��Y���������˗7��FTFG>������{�Z��� �k��� ��YD�'@ � 8n�R�� Uӱ$HEI3GHd�:h?(! 'v�������� �c Gd��qp$B% x� E��SHIF��hRVn�F�`�HpC� 3�(�8H`O� ѡ�C��+%D	�"��CE�pV���SP�HERs� � �,! M�c�u��$�POWERFL ��R|����|�p�RyG�`���������A� E ��?`��`d���NSb ����?�  �Bz|� l�  <k@�|��%�涀�˃����ŵ�� �2ӷ�� 	H���l&���>ߪ��A |��t]$��*��/�� **:��`�ϥ�d�͘���������ɘ��|�����5� ������%ߟ�I�[� ��ߑ��������� ��w�!�3�a�W�i��� ���������O���� 9�/�A���e�w����� ��'����� =O}s���� ���k'UK ]������C/ ��-/#/5/�/Y/k/ �/�/�/?�/�/?�/ ?�?1?C?q?g?y?�? �?�?�?�?�?_O	OO�IO?OQO�� 	  �O�O�O_�E��3_����O`_�O�_�_÷PR�EF Ӻ`�`
��IORITCY `|���`�����pSPL`z����WUqT�VqÈ�ODU~������_?�O�G��Gx��R��,fH�IBqOy�|kTO?ENT 1��yP?(!AF_b�`��o�g!tcp|�o}!ud�o~)~!icm��0bXY̳�k ;�|�)� ����������u� �����N�5�r� Y�������̏�����	*/c̳ӹ���E��W�|�>�Χ�FB��/��4���|��,��7�A��,  ��P����%�|�
'���Z��h�z������|��ENHA?NCE 	#�7��A9�d�����  �,f�T
�_�S��=��PORTe�rb����U��_C?ARTREP�Pr|>brSKSTAg�koSLGS�`�k������Unothing���� ��Ϳ>�P�b�To��TEMP ?i�sϨE/�_a_seibanm_��i_ �����0��T�?�x� cߜ߇ߙ��߽����� ��>�)�N�t�_�� ������������ :�%�^�I���m����� ������ ��$H 3lWi���� ���D/h S�w���uϪ��VERSI�P=g�  disa�ble��SAV�E ?j	2670H705�	�k/!�m//*��/ 	�(%b�O�+�/�Se?6?H?Z?l?�z:%<�/�?4�*'_�j` 1�kX ��0ubuE�?OqG�PURGE��Bp`�ncq�WF<@�a�TӒ*fW��`]Daa�WRUP�_DELAY �z�f�B_HOT %?e'b��OnE�R_NORMAL��HGb�O%_�GSEM�I_*_i_�QQSKKIP�3.��3x� �_��_�_�_�]?eo +goKo]ooo5o�o�o �o�o�o�o�o�o5 GYi�}�� �����1�C�U� �y�g���������я�����-�?�7%�$�RACFG ،[ќ�3�]�_P/ARAM�Q3y��Sw @И@`�G��42C۠��2���CbFB�B]�B�TIF���J]�CV�TMOU����]�]�DCR�3�Y� ��Q@��.�B�'B���@�o?��H<�x�]��s ��8�5��J�Ѽ��;��_��o ;e��m���KZ;�=�g;�4�<<����f@����� �5�G�Y�k�}��������ſ׿���xUR�DIO_TYPE�  �V�5��ED_PROT_a�&g>��4BHbC�EސSǆQ2c� ��B�ꐪϸ� ��ϐ����&�ݹ� W�V_~�o����߱� ��������A�O�m� r���9������� �������=�_�d��� ������������� ��'I�Nm�� �������# EJi+k�� ����//4/F/ /g//�/y/�/�/�/ �/�/	?+/0?O/?c? Q?�?u?�?�?�?�?�?�?;?,O��S�INT� 2�I���l�G;� jO|K��鯤O�f�0 �O�K�? �O�?___N_<_r_ X_�_�_�_�_�_�_�_ �_&ooJo8ono�ofo �o�o�o�o�o�o�o" F4j|b�� �������B��O�EFPOS1 �1"�  xO��o×O����ݏ 鈃���Ϗ0��T�� x����7���ҟm��� �����>�P����7� ������W��{���� �:�կ^�������� ��S�e��� ��$Ͽ� H��l��iϢ�=��� a��υ�� ߻���� h�Sߌ�'߰�K���o� ��
��.���R���v� ��#�5�o������� ���<���9�r���� 1���U����������� 8#\����? ��u��"�F X�?���_ ��/�	/B/�f/ /�/%/�/�/[/m/�/ ?�/,?�/P?�/t?? q?�?E?�?i?�?�?O (O�?�?OpO[O�O/O �OSO�OwO�O_�O6_ �OZ_�O~_�_+_=_w_ �_�_�_�_ o�_Do�_�Aozocf�2 1 r�o.oho�o�o
o .�oR�oO�#� G�k����� N�9�r����1���U� ���������8�ӏ\� ��	��U�����ڟu� ����"����X��|� ���;�į_�q����� �	�B�ݯf����%� ����[���ϣ�,� ǿٿ�%φ�qϪ�E� ��i��ύ���(���L� ��p�ߔ�/�A�Sߍ� ������6���Z��� W��+��O���s��� ������V�A�z�� ��9���]������� ��@��d��#] ���}�*� '`���C� gy��&//J/� n/	/�/-/�/�/c/�/ �/?�/4?�/�/�/-? �?y?�?M?�?q?�?�? �?0O�?TO�?xOO�O<�o�d3 1�oIO [O�O_�O7_=O[_�O __|_�_P_�_t_�_ �_!o�_�_�_o{ofo �o:o�o^o�o�o�o �oA�oe �$6 H�����+�� O��L��� ���D�͏ h�񏌏�����K�6� o�
���.���R���� �����5�ПY���� �R�����ׯr����� ����U��y���� 8���\�n������� ?�ڿc�����"τϽ� X���|�ߠ�)����� ��"߃�nߧ�B���f� �ߊ���%���I���m� ��,�>�P������ ���3���W���T��� (���L���p������� ����S>w�6 �Z����= �a� Z�� �z/�'/�$/]/ ��//�/@/�/�O�D4 1�Ov/�/�/ @?+?d?j/�?#?�?G? �?�?}?O�?*O�?NO �?�?OGO�O�O�OgO �O�O_�O_J_�On_ 	_�_-_�_Q_c_u_�_ o�_4o�_Xo�_|oo yo�oMo�oqo�o�o �o�o�oxc�7 �[����>� �b����!�3�E�� ��ˏ���(�ÏL�� I������A�ʟe�� �������H�3�l�� ��+���O���ꯅ�� ��2�ͯV����O� ����Կo�����Ϸ� �R��v�Ϛ�5Ͼ� Y�k�}Ϸ���<��� `��τ�߁ߺ�U��� y���&�������� ��k��?���c���� ��"���F���j���� )�;�M��������� 0��T��Q�%��I�m��/�$5 1�/���mX ���P�t�/ �3/�W/�{//(/ :/t/�/�/�/�/?�/ A?�/>?w??�?6?�? Z?�?~?�?�?�?=O(O aO�?�O O�ODO�O�O zO_�O'_�OK_�O�O 
_D_�_�_�_d_�_�_ o�_oGo�_koo�o *o�oNo`oro�o�o 1�oU�oyv� J�n����� ��u�`���4���X� �|�ޏ���;�֏_� �����0�B�|�ݟȟ ���%���I��F�� ���>�ǯb�믆��� ���E�0�i����(� ��L���翂�Ϧ�/� ʿS�� ��LϭϘ� ��l��ϐ�ߴ��O� ��s�ߗ�2߻�V�h� zߴ�� �9���]��� ���~��R���v�����#�	6 1 &������������� ��}���<��` ����CUg� �&�J�n	 k�?�c��/ ���	/j/U/�/)/ �/M/�/q/�/?�/0? �/T?�/x??%?7?q? �?�?�?�?O�?>O�? ;OtOO�O3O�OWO�O {O�O�O�O:_%_^_�O �__�_A_�_�_w_ o �_$o�_Ho�_�_oAo �o�o�oao�o�o�o D�oh�'� K]o�
��.�� R��v��s���G�Џ k�􏏏���ŏ׏� r�]���1���U�ޟy� ۟���8�ӟ\����� �-�?�y�گů���� "���F��C�|���� ;�Ŀ_�迃������ B�-�f�ϊ�%Ϯ�I� �����ߣ�,���P�<6�H�7 1S��� �I��߲������� 3���0�i���(�� L���p�����/�� S���w����6����� l�������=���� ��6���V�z � 9�]�� �@Rd��� #/�G/�k//h/�/ </�/`/�/�/?�/�/ �/?g?R?�?&?�?J? �?n?�?	O�?-O�?QO �?uOO"O4OnO�O�O �O�O_�O;_�O8_q_ _�_0_�_T_�_x_�_ �_�_7o"o[o�_oo �o>o�o�oto�o�o! �oE�o�o>�� �^�����A� �e� ���$���H�Z� l�����+�ƏO�� s��p���D�͟h�� �����ԟ�o�Z� ��.���R�ۯv�د� ��5�ЯY���}�c�u�8 1��*�<�v� ��߿��<�׿`��� ]ϖ�1Ϻ�U���y�� �ϯ�����\�G߀�� ��?���c����ߙ�"� ��F���j���)�c� ���������0��� -�f����%���I��� m������,P�� t�3��i� ��:���3 ��S�w /� �6/�Z/�~//�/ =/O/a/�/�/�/ ?�/ D?�/h??e?�?9?�? ]?�?�?
O�?�?�?O dOOO�O#O�OGO�OkO �O_�O*_�ON_�Or_ __1_k_�_�_�_�_ o�_8o�_5ono	o�o -o�oQo�ouo�o�o�o 4X�o|�; ��q����B� ���;�������[� ������>�ُb������!�������MA_SK 1 ��������ΗXNO � ݟ���MOT�E  ���S�_C_FG !Z����N�����PL_RA�NGV�N������O�WER "���Ϡ��SM_DRY�PRG %����%W��եTART� #Ǯ�UME_PRO���q����_EXEC_EN�B  ����GScPDJ�������gTDB����RMп���IA_OPTI�ON������~�NGVERS���`�řI_�AIRPUR�� �R�+���ÛMT_�֐T X���ΐO�BOT_ISOLC��������u������NAME8���H�ĚOB_CAT#EG�ϣ,��S��[�.�ORD_NU�M ?Ǩ���H705  �N��ߨߺ�ΐPC�_TIMEOUT��� xΐS232�s�1$��� L�TEACH ?PENDAN��o�,�����V�T��Mainten�ance Con%sN�&�M�"B�P�No Use6� r�8��������̒���NPO$��Ҋ�z"���CH_LM��Q���	a�,�!�UD1:��.�R�ՐVAILw���粥*�SR  �t� ���5�R_�INTVAL�ᐲ� ���V_D�ATA_GRP �2'���� D��P�������	 ������ B0RTf��� ���/�/>/,/ b/P/�/t/�/�/�/�/ �/?�/(??L?:?p? ^?�?�?�?�?�?�?�? O O"O$O6OlOZO�O ~O�O�O�O�O�O_�O 2_ _V_D_z_h_�_�_ �_�_�_�_�_o
o@o�.oPovodo�o��$�SAF_DO_PULSW�[�S���i�OSCAN��������SCà(/�߈0���WS�S�
����Ķ�q�q�qN�  �L^p���5���� ��$��+��r2M�qX��dM�h�J�	t/� @��������ʋ|�� r ք��_ @N�T ��'��9�K�X�T D��X���������ɟ۟ ����#�5�G�Y�k��}�������䅎������Ǧ  ="�;�oR� ����p"�
�u��Di���q$q�?  � ���u q��\�������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$�6�H�Z����珈�� �����������g� ;�D�V�h�z�������@��������(�Ӣ0� r�i�y���$�7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/?r�+? =?O?a?s?�?�?�?�? �?8��?OO'O9OKO ]OoO�O��$�r�O �O�O�O	__-_?_Q_ c_u_�_�Y�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|�c�路g����� ��0�B�T�f�x����������ҏ����p��:�Ҧ��y��3�	�	123�45678��h�!B!�� +\��p0�� ��Ο�����(�:� @��c�u��������� ϯ����)�;�M� _�q�����R���ɿۿ ����#�5�G�Y�k� }Ϗϡϳ����ϖ��� ��1�C�U�g�yߋ� �߯���������	�� -���Q�c�u���� ����������)�;� M�_�q���B������ ����%7I[ m������� �!3EWi{ �������/ ///�S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?D/�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O*����O	_�E�?5_�G_Y_�yCz  �A��z   ���x2�r }��)�
�W_�  	�*�2�O �_�_ oo"l�#\��_hozo�o�o�o�o �o�o�o
.@R dv����Mo� ���*�<�N�`�r� ��������̏ޏ��� �&�8�J��X #P$Pt�Q�R<u� k�~�Q  �������S�P���Q�Qt�  �PÙ۟�P(� `,b����]��PFl�$SCR_�GRP 1*0�+04� �� �,a ��U	 v��~������ d���%���ɯ���h]���P�D1� D7n��3��Fl�
CRX-10�iA/L 234�567890�P�d� r��Pd�L ��,a
1o�����Z���[ ¶~� +fm�ͣm�Fcg�p�����ӹ	Ĳ�.�@��R�d�t���H�~�Ă�m��ϴ�@�����ϼ��,a�Ϡ1���U�[�G�imXh�uP,[~;�B�  BƠߞҷ�r��A�P��  @1`��՚�@����� ?	���H����ښ�F@ F�`A� I�@�m�X��|���� ��������������`:�%�7�I�[�B�i� ��������������� -Q<u`��@En�ٯ���W�P�"+f@_�5��1`4b���x����ͣ�O�,dA����$���Fa�,a �#!"/4/E-!�Z(f/x/G/ (�P�!(� �/�/�/��/�/?#9b�����S7س�M�ECLV�L  ,a���ݲ�Q@f1L_D?EFAULTn4b1_�1`�3?HOTSTR�=���2MIPOWER�Fm0pU�5�4W7FDO�6 �5L��ERVENT 1�+u1u1�3 L!�DUM_EIP�#?5H�j!AF�_INE�0SO,d!'FT)O�NIO�O9!���O ��O�O�!RPC_MAIN�O�H��O>_S'VIS_�I�-_�_?!OPCUf�_�Wy_�_!TMP�PPU�_<Id�_�"o!
PMON_�PROXY#o?Fe ono�R<o8Mf]o�o�!RDM_SR�V�o<Ig�o!�R��"=Hh�oR!%
PM�o9LiA��!RLSYNC̟�y8��!gROS(O��4��6�!
CE�PMT'COM7�?Fk%���{!	K�CONS���>Glq�Ώ!K�WOASRC�o?Fm��v�!K�USB��=Hn	�f�!STM�0��;JoU����O�֟�c����CICE�_KL ?%K� (%SVCPGRG1��G�1�2G�DL�6�3o�t�6�4��D��6�5��į6�6��6�7��6���W�R�9_�d�3��� 6�9���6�a�ܿ6��� �6���,�6�ٯT�6� �|�6�)���6�Q��� 6�y���^����^�ʿ D�^��l�^�ϔ�^� Bϼ�^�j���^���� ^���4�^���\�^�
� �2���6��/� ���V��<�'�`�K� ��o����������� ��&J5nY� ������� 4F1jU�y� ����/�0// T/?/x/c/�/�/�/�/ �/�/�/??>?)?P?�t?_?�?
�_DEV� I�M{C:�84���4?GRP 2/E�0�+�bx 	�/ 
 ,@�?O ��ODO+OhOOOaO�O �O�O�O�O�O�O__ @_R_9_v_]_�_�_O �_�_�_o�_*ooNo `oGo�oko�o�o�o�o �o�o&8\�_ Q�I����� ��4�F�-�j�Q��� ����ď���Ϗ�� uB�T�;�x�_����� ��ҟ����ݟ�,�� P�7�t���m�����ί �7����(�:�!�^� E�����{�����ܿÿ տ���6��Z�l�S� ��篅���}������  ��D�+�h�z�aߞ� �����߻������� �R��v��o��� ��������*��N� `�G���k��������� ��k�8��\n U�y����� �	F-jQ� ������/ /B/T/;/x/_/�/�/ �/�/�/�/?�/,??�P?7?I?�?�3d ��6	t?�?�?�?�?O�?)O8K%�8O]O����vA"AvE�O �G~O�O�O�O�O�O
Y JO/_rI�O\_J_�_n_ �_�_�_�__o@_�_ 4o"oXoFo|ojo�o�_ o�oo�o�o0 TBx�o��oh� d���,��P�� w��@�����Ώ��ޏ ��(�j�O������ p�����ʟ��ڟ �B� '�f��Z�H�~�l��� ��Ư������د��  �V�D�z�h����ſ �������
��R� @�vϸ���ܿf��Ͼ� �������Nߐ�u� ��>ߨߖ��ߺ�����  �V�|�M��&��n� ��������.��R� ��F���V�|�j����� �����*���B 0Rxf���� ���>,N t���d��� �//:/|a/s/*/ L/&/�/�/�/�/�/? T/9?x/?l?Z?|?~? �?�?�?�?,?OP?�? DO2OhOVOxOzO�O�O O�O(O�O_
_@_._ d_R_t_�O�O�_ _�_ �_�_oo<o*o`o�_ �o�_Po�oLo�o�o�o 8zo_�o(� �������R 7�v �j�X���|��� ���*��N�؏B� 0�f�T���x�����՟ 矞������>�,�b� P���ȟ���v��ί ���:�(�^����� įN�����ܿʿ��  �6�x�]Ϝ�&ϐ�~� �Ϣ�������>�d�5� t��h�Vߌ�z߰ߞ� �����:���.���>� d�R��v������� �����*��:�`�N� �������t����� ��&6\����� L������" dI[4|� ����<!/`� T/B/d/f/x/�/�/�/ /�/8/�/,??P?>? `?b?t?�?�/�??�? O�?(OOLO:O\O�? �?�O�?�O�O�O _�O $__H_�Oo_�O8_�_ 4_�_�_�_�_�_ ob_ Go�_ozoho�o�o�o �o�o�o:o^o�oR @vd���� �6�*��N�<�r� `������Ϗ������ ��&��J�8�n����� ԏ^�ȟ��؟ڟ�"� �F���m���6����� į��ԯ֯��`�E� ���x�f��������� п&�L��\���P�>� t�bϘφϼ�����"� ��ߨ�&�L�:�p�^� ���ϻ��τ������  �"�H�6�l�ߓ��� \������������ D���k���4������� ������
L�1C�� ��d����� $	H�<*LN `����� � //8/&/H/J/\/�/ ��/��/�/�/?�/ 4?"?D?�/�/�?�/j? �?�?�?�?O�?0Or? WO�? O�OO�O�O�O �O�O_JO/_nO�Ob_ P_�_t_�_�_�_�_"_ oF_�_:o(o^oLo�o po�o�o�_�oo�o  6$ZH~�o� �n�j���2�  �V��}��F����� ��ԏ
���.�p�U� �����v��������� П�H�-�l���`�N� ��r��������4�� D�ޯ8�&�\�J���n� ���˿
�������� 4�"�X�F�|Ͼ���� l���������
�0�� Tߖ�{ߺ�D߮ߜ��� �������,�n�S�� ��t�������� 4��+������L��� p����������0��� $46H~l� ������  02Dz���j ����/
/,/� �y/�R/�/�/�/�/ �/�/?Z/??~/?r? ?�?�?�?�?�?�?2? OV?�?JO8OnO\O~O �O�O�O
O�O.O�O"_ _F_4_j_X_z_�_�O �__�_�_�_ooBo 0ofo�_�o�oVoxoRo �o�o�o>�oe �o.������ ��X=�|�p�^� �����������0�� T�ޏH�6�l�Z���~� ������,�Ɵ �� D�2�h�V���Ο��� |��x����
�@�.� d�����ʯT������ п���<�~�cϢ� ,ϖτϺϨ������� �V�;�z��n�\ߒ� �߶ߤ�������� ����4�j�X��|�� ����������� 0�f�T��������z� ������,b �����R���� �j�a�: ������ /B '/f�Z/�j/�/~/ �/�/�//�/>/�/2?  ?V?D?f?�?z?�?�/ �??�?
O�?.OORO @ObO�O�?�O�?xO�O �O_�O*__N_�Ou_ �_>_`_:_�_�_�_o��_&oh_Mo�_�Q�$�SERV_MAI�L  �U�`�~rhOUTPUT�h_�P@vd�RV 20f  �` (a\o�ovd�SAVE�l�iTO�P10 21�i d �_HZl ~������� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d�v������� ��П�����*�<��euYPscFZ�N_CFG 2e�c�T�a�e~|�GRP 23���q ,B   �AƠ�QD;� B}Ǡ�  B4�S�RB21�fH7ELL�4ev��`�o��/�>�%RSR>�?�Q���u� ����ҿ������,π�P�;�t�_Ϙϩ�~���  � �����Ϸͻ��P��&�'�ސW��2Pd��g��HKw 15�� ,� �߫ߥ��������� @�;�M�_���������������OMM� 6��?��FT?OV_ENB�d�a�u�OW_REG�_UI_�tbIMI_OFWDL*�7.��ɥ��WAIT\� `ٞ����`���d��wTIM�������VA�`����_UNcIT[�*yLCy�WTRY��uv`ME�8���aw�rdt ��9� ������<���X�Pڠ6p`?� � ��o+=1`VL�l�f�MON_ALIA�S ?e.��`heGo������ /)/;/M/�q/�/�/ �/�/d/�/�/??%? �/I?[?m??�?<?�? �?�?�?�?�?!O3OEO WOO{O�O�O�O�OnO �O�O__/_�OS_e_ w_�_�_F_�_�_�_�_ �_o+o=oOoaoo�o �o�o�o�oxo�o '9�o]o��> ������#�5� G�Y�k��������ŏ ׏������1�C�� g�y�����H���ӟ� ��	���-�?�Q�c�u�  �������ϯᯌ�� �)�;��L�q����� ��R�˿ݿ��Ͼ� 7�I�[�m��*ϣϵ� �����ϖ��!�3�E� ��i�{ߍߟ߱�\��� ��������A�S�e� w��4�������� ���+�=�O���s��� ������f����� '��K]o��> �����#5 GY}�����l�$SMON_�DEFPROG �&����� &*S?YSTEM*����RECALL �?}� ( ��}3xcopy �fr:\*.* �virt:\tm�pbackT!=>�192.168.�56.1:36400 z"�/�/�/�,}4K%aS/e/w%�/�?#?5? }
xy�zrate 11 �/�/�/�?�?�?�%K7k?| j?|?OO�1O�#tpdisc 0�?| �?�?�O��O�OBHconn ��?dOvO__+_�)8�L$s:orderfil.datY<`�O_�_�_�_}/L"mdb:V?o_| {_ oo0o�$J/]?n/ o �o�o�o�/Yoko�O !3F_X_�_�_�� ��_�_q�_��/� Bo�o�oxo�������o �oc��o��+�>?P? �􏅟�����?�?u�21696�O{���0�C� ֟����� ����ԟf�x�	�� -�@ORM�����������D0U�e�w� ��,�?�Q�ֿ��� �ϝϯ�¯ԯ�x�	� �-�@R��˃ߕ� �ߺ�g���{��� 0�C���h����ߐ�� ��ǏX�j�e����$� 6�I������������ ������}� 2E� �����������k gy
.A�S��� w߈������l�� //*/=�O�b�s�/ �/�/����^/��/? &?9K��/�/?�?�? �?���??O"O4O G�?�?�?�O�O�O�? mOiO{O__0_CU �y�_�_�_��n_��oo,o>W�$S�NPX_ASG �2:���Va�  ��%�7o~o  ?��GfPARAM �;Ve`a �U	lkP>TDP>X~�d� ��I`�OFT_KB_CFG  CS\eFc�OPIN_SIMW  Vk�b+�=OYsI`RVNO�RDY_DO  ��eukrQST_P_DSB~�b|�>kSR <Vi� � & TELEO�e�{v>T�W`I`TOP_ON�_ERRxGb�P_TN VeP���D:�RIN�G_PRM'��rV�CNT_GP 2�=Ve�ac`x 	 ���DP��я����Bg�VD�RP 1>�i�`�Vq؏0�B� T�f�x���������ҟ �����,�>�e�b� t���������ί�� �+�(�:�L�^�p��� ������ʿ�� �� $�6�H�Z�l�~ϐϷ� ����������� �2� D�V�}�zߌߞ߰��� ������
��C�@�R� d�v��������� 	���*�<�N�`�r� �������������� &8J\n�� ������" 4[Xj|��� ����!//0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�?�O�PRG_CO7UNT�f�P�)I'ENBe�+EMUC�d�bO_UPD 1?>�{T  
ODR �O�O�O�O�O__A_ <_N_`_�_�_�_�_�_ �_�_�_oo&o8oao \ono�o�o�o�o�o�o �o�o94FX� |������� ��0�Y�T�f�x��� �����������1� ,�>�P�y�t������� ��Ο��	���(�Q� L�^�p���������� ܯ� �)�$�6�H�q� l�~�������ƿؿπ��� �I�D�V�"L_INFO 1@�E��@��	 �yϽϨ����ɻ����?zN>?�>�����B�]����l�^���e��¤���C*p���n�?j�` <�`�o�� C���B����C���C0��T�����Gwp߂�-@YSDOEBUG:@�@�o��d�I��SP_PA�SS:EB?��L_OG A���A�  o�i�v� � �Ao�UD�1:\��}���_M�PC�ݚEk�}�A�&�� �AK�SAV B��IA���*�i�1�SVB�T�EM_TIME �1C���@ 0"�@?|D#�o�@��"����MEMBK  	�EA�����^��X|�@�6�i�����������h�9
�� ��@ �`r�����`��� � @Rdv�����
Le�//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z?��SKV�[�EAj��?X�?�?��7o�j]2���?i� �.^ 
:O.@R�O�O�O8}N��2� ��OB�C��O_&_8_,M2�Y_�_�_�_�_�_o�$�_�_�o'o9o Ko]ooo�o�o�o�o�o �o�o�o#5GY�k_?T1SVGU�NSPD�� '�����p2MODE_LIM D�d�Ҋt2�p�qE����uABUI_DCOS H}5���0 �G��E�C��|-�X��>���*���� !
��e��i���r��i�����uED�IT I��xS�CRN J��<�rS�G K��G� �0߅SK_OPTION��^�����_DI��ENB�  C����BC�2_GRP 2L����MPC��ʓ�|BCCF/�ND�� ]����Z� =�V�A�S���w����� ԯ������.��R� =�v�a����������� ��߿��<�'�`�K� �ϖ�Ĉ�϶������� v��
�/�U�@�yߧ� ��`�iМ��߰����� 
���.��>�@�R�� v����������� *��N�<�r�`����� ����������̀ 4FX��|j�� �����B 0fTvx��� ��/�,//</b/ P/�/t/�/�/�/�/�/ �/�/(??L?d?v? �?�?�?6?�?�?�?O  O6OHOZO(O~OlO�O �O�O�O�O�O�O __ D_2_h_V_�_z_�_�_ �_�_�_
o�_.oo>o @oRo�ovo�ob?�o�o �o�o<*Lr `������� �&��6�8�J���n� ����ȏ���ڏ��"� �F�4�j�X���|��� �����֟��o$�6� T�f�x���������ү �������>�,�b� P���t��������ο ��(��L�:�\ς� pϦϔ��ϸ�������  ��H�6�l�"��ߖ� ������V������2�  �V�h�z�H����� ����������
�@�.� d�R���v��������� ����*N<^ `r������� &8�\Jl� �������"/ /F/4/V/X/j/�/�/ �/�/�/�/?�/?B? 0?f?T?�?x?�?�?�? �?�?O�?,O�DOVO tO�O�OO�O�O�O�O��O_ V4P�$TB�CSG_GRP �2O U��  �4Q 
 ?�  __q_[_ �__�_�_�_�_�_o�%k8R?SQF\dאHTa?4Q	 �HA���#e>�w��>$a�\#e?AT��A WR�o��hdjma�G�?L�fg�bp�o�n�ff�hf��ͼb4P|j���o*}@��Rhf�?ff>�33pa#eB<qB�o+=xrRp�qUy�rt~��H`�y rIpTv�pBȺ t~	xf	x(�;��� f���N�`���ˏڋ�����	V3.0�0WR	crxlڃ	*��3R~td��HH��� \��.�]�  cC�.�����8QJ2?SR�F]����CFG [T UPQ SPVܚ��r�ܟ1��1�W�e�	P e���v�����ӯ���� ����Q�<�u�`� ��������Ϳ�޿� �;�&�_�Jσ�nπ� �Ϥ�������WRq@ �0�B���u�`߅߫� ���ߺ������)�;� M��q�\������ 4Q _���O ���J� 8�n�\����������� ������4"XF hj|����� �.TBxf ��nO����/ />/,/b/P/�/t/�/ �/�/�/�/�/�/?:? (?^?p?�?�?N?�?�? �?�?�?�? O6O$OZO HO~OlO�O�O�O�O�O �O�O __D_2_T_V_ h_�_�_�_�_�_�_
o �_o@o�Xojo|o&o �o�o�o�o�o�o* N`r�B�� �����&��6� \�J���n�����ȏ�� ؏ڏ�"��F�4�j� X���|���ğ���֟ ���0��@�B�T��� x�����ү䯎o��� ̯ʯP�>�t�b����� ���������Կ&� L�:�p�^ϔϦϸ��� ������� �"�H�6� l�Zߐ�~ߴߢ����� �����2� �V�D�z� h������������ �
�,�.�@�v��� ����\������� <*`N���� x���8J \(����� ���/4/"/X/F/ |/j/�/�/�/�/�/�/ �/??B?0?f?T?v? �?�?�?�?�?�?OO ��2ODO�� O�OtO�O �O�O�O�O_�O(_:_ L_
__�_p_�_�_�_ �_�_ o�_$oo4o6o Ho~olo�o�o�o�o�o �o�o D2hV �z�����
� �.��R�@�b���v� ��&OXO֏菒���� �N�<�r�`������� ̟ޟ🮟��$�&� 8�n�������^�ȯ�� �گ��� �"�4�j� X���|�����ֿĿ� ���0��T�B�x�f� �ϊϜ���������� �>�P���h�zߌ�6� �ߪ����������:� (�^�p���R���p���� ���  &��*� *�>�*���$TBJOP_G�RP 2U����  ?_���C*�	V��]�Wd������X  �*��� �,? � ���*� @&�?��	� �A�����C�  DD������>v�>\?� ��aG�:��o��;ߴAT3������A�<���MX����>��\�)?���8Q������L��>̼0 &�;iG.���Ap< � F�A�ff�v��� �):VM�.��� S>o*�@��R�Cр	����p�����ff��:�6/�?�3=3�B   �� /������>)/:�S���� <�/�/@��H�%&/и/��=� <#��
*��v�;/��ڪ!?���4B� 3?'?2	��2?hZ? D?R?�?�?�?F?�?�? �?�?OAOO�?`OzO`dOrO�O�O*�C�*����A��	V3.�00{�crxl��*P��%�%c�5Z F� �JZH F6� �F^ F�� �F�f F� �G� G5 �G<
 G^] �G� G����G�*�G�S G�; G��ER�Du�\E[� �E� F( �F-� FU` �F}  F�N �F� F�� �Fͺ F� �F�V G� �Gz Ga O9ѷ�Q�LHe�fJ4�o,b*��0c1���OH�ED_?TCH Xd�+X�2S�&�&�dA$'X�o�o*�1F��TESTPARS�  ��cV�HR�pABLE 1Yd� N`*����R�g$j�g�h�h�)�1��g	�h
�h��hHu*��h�h:�h%vRDI0n�GYk}��u	�O�#�-�?�Q�c�u�)rS�l� �z6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z���I���m�Fwͩ ��ȏڏ쏘������x)r��NUM [ ��n����2� Ep�)r_CFG Z��I����@V�IMEBF_�TTqD��e޶V�ER�����޳R� 1[8{ 8$�o*�%�Q� ��د  9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}��ߡ߳� ����������1��� E�W�i�{������ ��������/�A�S� e�w����������������+=O�_Ԗ��@��`LIoF \��D`B����DR�(FP�
�!p�!p� �d� ��MI_CH�AN� � D_BGLVL��f�ETHERAD� ?u��0`�1�_}�ROUmT�!�j!���SNMASK�Y�j255.�%S///A/S�`O�OLOFS_DI�p�CORQC?TRL ]8{��1o�-T�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OL�/6O�%OZOcPE_DE�TAI7�*PGL�_CONFIG �c������/�cell/$CID$/grp1^O@�O�O�O
__|��� G_Y_k_}_�_�_0_�_ �_�_�_oo�_CoUo goyo�o�o,o>o�o�o �o	-�oQcu ���:���� �)���_�q���������׮}N�����%�7�I�a�KOq�P�� M�����ʟܟ� �G� $�6�H�Z�l�~���� ��Ưد������2� D�V�h�z������¿ Կ���
ϙ�.�@�R� d�vψϚ�)Ͼ����� ���ߧ�<�N�`�r� �ߖ�%ߺ�������� �&��J�\�n��� ��3����������"� ��F�X�j�|���������@�User� View �I}�}1234567890����+`=Ex �e����2��B������`r��3�Oa�s����x4 >//'/9/K/]/�~/x5��/�/�/�/ �/?p/2?x6�/k? }?�?�?�?�?$?�?x7Z?O1OCOUOgOyO�?�Ox8O�O�O�O�	__-_�ON_TR �lCamera���O�_�_�_�_�_�_˂E�_o)o;n ��Uogoyo�o�o�o�)  mV�	�_�o# 5GY o}���o�������F_� mV=�k�}������� ŏl����X�1�C� U�g�y���2�D��"� ן�����1�؏U� g�y�ğ������ӯ� ����D��k��E�W�i� {�����F�ÿտ�2� ��/�A�S�e��nU Y9������������	� ��-�?�Qߜ�u߇ߙ� �߽���v�D�If�� -�?�Q�c�u�ߙ�� ���������)�;� ��D��I��������� ������)t�M�_q���N�`�9 3��0B�� Sx�1����P�//�J	oU0� U/g/y/�/�/�/V�/ �/�/�?-???Q?c? u?/./tPv[?�?�? �?OO(O�/LO^OpO �?�O�O�O�O�O�O�? oU�k�O:_L_^_p_�_ �_;O�_�_�_'_ oo $o6oHoZo_;%N��_ �o�o�o�o�o �_$ 6H�ol~��� �moe��]�$�6� H�Z�l�������� ؏���� �2��e &�ɏ~�������Ɵ؟ ���� �k�D�V�h� z�����E�e��5�� ��� �2�D��h�z� ��ׯ��¿Կ���
���  ��9�K� ]�oρϓϥϷ�����<����   �� 5�G�Y�k�}ߏߡ߳� ����������1�C� U�g�y�������� ����	��-�?�Q�c� u��������������� );M_q��  
��(  }�-�( 	 � ������# 35G}k���:�
� �Y�
/ /./��R/d/v/�/�/ �/����/�/�/A/? 0?B?T?f?x?�/�?�? �??�?�?OO,O>O �?bOtO�O�?�O�O�O �O�O_KO]O:_L_^_ �O�_�_�_�_�_�_#_  oo$ok_HoZolo~o �o�o�_�o�o�o1o  2DVh�o�o� ��	��
��.� @��d�v�������� Џ���M�*�<�N� ��r���������̟� %���&�m�J�\�n� �������ȯگ�3� �"�4�F�X�j����� ������ֿ����� 0�w���f�xϊ�ѿ�� ���������O�,�>� Pߗ�t߆ߘߪ߼��� �����]�:�L�^��p����߻@  ����������� ���"frh:\�tpgl\robots\crx!��10ia_l.xml��D�V�h�z������������������ ��0BTfx� �������� ,>Pbt��� �����/(/:/ L/^/p/�/�/�/�/�/ �/��/?$?6?H?Z? l?~?�?�?�?�?�?�/ �?O O2ODOVOhOzO �O�O�O�O�O�?�O
_ _._@_R_d_v_�_�_ �_�_�_�O�_oo*o <oNo`oro�o�o�o�o��o�n �6� |���<< 	� ?��k!�o; iOq����� ����%�S�9�k�@��o�����я�����(�$TPGL_�OUTPUT �f������ �&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��������į�p�ր2�345678901�����1�C�K� ���r���������̿ d�п��&�8�J��}T�|ώϠϲ���\� n�����0�B�T��� bߊߜ߮�����j��� ��,�>�P����߆� ��������x���� (�:�L�^���l����� ������t���$6 HZlz��� ���� 2DV h ����� ��/./@/R/d/v/ /�/�/�/�/�/�/�/~ۂ $$�� ί<7*?\?N?�?r?�? �?�?�?�?�?OO4O &OXOJO|OnO�O�O�O �O�O�O_�O0_"_T_}�an_�_�_�_�_�_��]@�_o	z ( 	 V_Do2o hoVo�ozo�o�o�o�o �o
�o.R@v d������� ��(�*�<�r�`����ܦ�  <<I_ˏݏ����� ��:�L�֪��}���)� ��ş�������k�� C�ݟ/�y���e����� ��������-�?�� c�u�ӯ]�����W�� �Ϳ��)χ���_�q� �yϧρϓ�����M� �%߿��[�5�Gߑ� ��߫���s����!� ��E�W��?���9� ��������i���A� S���w���c�u���� /�����=) s�����U�� �'9�!o	 [�����K� #/5/�Y/k/E/w/�/ �/�/�/�/�/?�/ ?U?g?�/�?�?7?�?��?�?�?	OO��)�WGL1.XML��_PM�$TPOF?F_LIM ���P����^FNw_SVf@  �T�xJP_MON �g��zD�P��P2ZISTRTC�HK h��xF�k_aBVTCOMP�AT�HQ|FVWV_AR i�M:X.�D �O R_�P��BbA_DEFPROG %�I�%TELEO�Pi_�O_DISP�LAYm@�N�RIN�ST_MSK  ��\ �ZINU�SER_�TLCK�l�[QUICKM�EN:o�TSCRE�Y`��Rtpsc�Tat`yixB��`_�iSTZxIR�ACE_CFG �j�I:T�@	�[T
?��hHNL� 2k�Z���aA[  gR-?Qcu�����z�eITEM �2l{ �%$�12345678�90 ��  =<�
�0�B�J�  !P�X�dP���[S� ��"���X�
�|��� W���r�֏����.�� 0�B�\�f�����6�\� n�ҟ��������>� ��"���.�����ί R����Ŀֿ:��^� p�9ϔ�Tϸ�xϊ�� ���d���H��l�� >�Pߴ�\�������v�  ������h�(�ߞ� ��4�L��ߦ����� @�R��v�6���Z�l� ��������*���N� �� ������������ X���J
n ���b��� �"4F�/|</ N/�Z/���//�/ 0/�/?f/?�/�/e? �/�?�/�?�?�?,?�? P?b?t?�?�?DOjO|O �?�OOO(O�O�O^O _0_�O<_�O�O�_�O �__�_�_H_�_l_~_�Go�dS�bm�oLjψ  �rLj 8�a�o�Y
 �o�o��o�o{jUD1:�\|��^aR_G�RP 1n�{?� 	 @�PR d{N�r����~��p���q+��<O�:�?�  j�|� f����������ҏ� ���>�,�b�P���t�0��������	e����\cSCB 2ohk U�R�d�v����������Я�RlU�TORIAL �phk�o-�WgV_C�ONFIG q�hm�a�o�o��<�OUTPUT rhi}�����ܿ�  ��$�6�H�Z�l�~� �Ϣϴ�z�ɿ���� � �$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ����*<N` r�������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/��/�/??0? B?T?f?x?�?�?�?�? �/�?�?OO,O>OPO bOtO�O�O�O�O�?�O �O__(_:_L_^_p_ �_�_�_�_�_f�x�ǿ oo,o>oPoboto�o �o�o�o�o�o�O (:L^p��� ����o ��$�6� H�Z�l�~�������Ə ؏��� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я��� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t�����������������X���#�� N�_r����� ��&8J�� n������� �/"/4/F/X/i|/ �/�/�/�/�/�/�/? ?0?B?T?e/x?�?�? �?�?�?�?�?OO,O >OPOa?tO�O�O�O�O �O�O�O__(_:_L_ ^_oO�_�_�_�_�_�_ �_ oo$o6oHoZok_ ~o�o�o�o�o�o�o�o  2DVgoz� ������
�� .�@�R�d�u������ ��Џ����*�<� N�`�q���������̟ ޟ���&�8�J�\��k��$TX_SCREEN 1s%� �}�k�����ӯ���	���Z��I�[�m�� �����,�ٿ���� !�3Ϫ�W�ο{ύϟ� ������L���p��/� A�S�e�w��� ߭߿� �������~�+��O� a�s���� ���D� ����'�9�K����� ������������R��� v�#5GYk}�����$UALRM_MSG ?����� �n��� 	:-^Qc������� /�S�EV  ��2&�ECFG �u����  �n�@�  Ab! �  B�n�
  /u����/�/�/�/�/ �/??%?7?I?W7>!�GRP 2vH+; 0n�	 /�?�� I_BBL_N�OTE wH*T��lu�䐠w�T �2DEF�PRO� %� (%�Ow�	OBO-O fOQO�OuO�O�O�O�O��O_�O,_�<FKE�YDATA 1x<���0p W'n��?�_�_z_�_�_�Z�,(�_on�(POINT ERo�n  IRECT@oko�PNDUo�oOcCHOICE]�o�nTOUCHUP�o�o�o�o8 \nU�y�������"�	�F��Y���/frh/g�ui/white�home.png�Q�������ŏ׏�>h�pointz��`�/�A�S��  i�direc������p��şןf�/iny���"�4�F�X��m�choicy��������ͯ߯�h�touchup���/�A��S�e��h�arwrg�����ÿտ� n���(�:�L�^�p� ���Ϧϸ�������}� �$�6�H�Z�l��ϐ� �ߴ��������ߋ� � 2�D�V�h�z�	��� ����������.�@� R�d�v���_������� �������2DV hz����� �
�@Rdv ��)����/ /�</N/`/r/�/�/ %/�/�/�/�/??&? �/J?\?n?�?�?�?3? �?�?�?�?O"O�?4O XOjO|O�O�O�OAO�O �O�O__0_�OT_f_ x_�_�_�_=_�_�_�_ oo,o>o�_boto�oИo�o�oW��k�>b�����o }�o8J$v,6�{ .�������� �/��S�:�w���p� ����я�ʏ��+� �O�a�H���l����� ��ߟ���'�9�Ho ]�o���������ɯX� ����#�5�G�֯k� }�������ſT���� ��1�C�U��yϋ� �ϯ�����b���	�� -�?�Q���u߇ߙ߫� ������p���)�;� M�_��߃������ ��l���%�7�I�[� m�������������� z�!3EWi�� �������П /ASew~� �����/�+/ =/O/a/s/�//�/�/ �/�/�/?�/'?9?K? ]?o?�?�?"?�?�?�? �?�?O�?5OGOYOkO }O�OO�O�O�O�O�O __�OC_U_g_y_�_ �_,_�_�_�_�_	oo �_?oQocouo�o�o�o :o�o�o�o)�o M_q���6������%�7��9�����b�t���^�������,��돞����3�E� ,�i�P�������ß�� �������A�S�:� w�^�������ѯ���� ܯ�+�
O�a�s��� �����Ϳ߿��� '�9�ȿ]�oρϓϥ� ��F��������#�5� ��Y�k�}ߏߡ߳��� T�������1�C��� g�y������P��� ��	��-�?�Q���u� ����������^��� );M��q�� ����l% 7I[���� ��h�/!/3/E/ W/i/@��/�/�/�/�/ �/�??/?A?S?e? w??�?�?�?�?�?�? �?O+O=OOOaOsOO �O�O�O�O�O�O_�O '_9_K_]_o_�__�_ �_�_�_�_�_�_#o5o GoYoko}o�oo�o�o �o�o�o�o1CU gy����� �	���?�Q�c�u� ����(���Ϗ��� ���;�M�_�q��������~ ���~ ���ҟ���Ο�*��,�[��� f�������ٯ����� ��3��W�i�P���t� ��ÿ���ο��/� A�(�e�Lωϛ�z/�� ��������(�=�O� a�s߅ߗߩ�8����� ����'��K�]�o� ����4��������� �#�5���Y�k�}��� ����B������� 1��Ugy��� �P��	-? �cu����L ��//)/;/M/� q/�/�/�/�/�/Z/�/ ??%?7?I?�/m?? �?�?�?�?�?���?O !O3OEOWO^?{O�O�O �O�O�O�OvO__/_ A_S_e_�O�_�_�_�_ �_�_r_oo+o=oOo aosoo�o�o�o�o�o �o�o'9K]o �o������� �#�5�G�Y�k�}�� ����ŏ׏������ 1�C�U�g�y������ ��ӟ���	���-�?� Q�c�u��������ϯ������0�}��0���B�@T�f�>�����t�,�� ˿~��ֿ�%��I� 0�m��fϣϊ����� ������!�3��W�>� {�bߟ߱ߘ��߼��� ��?/�A�S�e�w�� ������������� ��=�O�a�s�����&� ����������9 K]o���4� ���#�GY k}��0��� �//1/�U/g/y/ �/�/�/>/�/�/�/	? ?-?�/Q?c?u?�?�? �?�?L?�?�?OO)O ;O�?_OqO�O�O�O�O HO�O�O__%_7_I_  �m__�_�_�_�_�O �_�_o!o3oEoWo�_ {o�o�o�o�o�odo�o /AS�ow� �����r�� +�=�O�a�������� ��͏ߏn���'�9� K�]�o���������ɟ ۟�|��#�5�G�Y� k���������ůׯ� �����1�C�U�g�y� �������ӿ����� �-�?�Q�c�uχ�^P����^P��������ͮ���
���,��;���_�F߃� ��|߹ߠ�������� ��7�I�0�m�T��� ����������!�� E�,�i�{�Z_������ �������/AS ew����� ��+=Oas ������/ /�9/K/]/o/�/�/ "/�/�/�/�/�/?�/ 5?G?Y?k?}?�?�?0? �?�?�?�?OO�?CO UOgOyO�O�O,O�O�O �O�O	__-_�OQ_c_ u_�_�_�_:_�_�_�_ oo)o�_Mo_oqo�o �o�o�o���o�o %7>o[m�� ��V���!�3� E��i�{�������Ï R������/�A�S� �w���������џ`� ����+�=�O�ޟs� ��������ͯ߯n�� �'�9�K�]�쯁��� ����ɿۿj����#� 5�G�Y�k����ϡϳ� ������x���1�C� U�g��ϋߝ߯�����h�����`����`���"�4�F��h�z�T�,f���^� ��������)��M� _�F���j��������� ����7[B �x�����o !3EWixߍ �������/ //A/S/e/w//�/�/ �/�/�/�/�/?+?=? O?a?s?�??�?�?�? �?�?O�?'O9OKO]O oO�OO�O�O�O�O�O �O_�O5_G_Y_k_}_ �__�_�_�_�_�_o �_1oCoUogoyo�o�o ,o�o�o�o�o	�o ?Qcu��(� �����)� M� _�q��������ˏݏ ���%�7�Ə[�m� �������D�ٟ��� �!�3�W�i�{��� ����ïR������ /�A�Яe�w������� ��N������+�=� O�޿sυϗϩϻ��� \�����'�9�K��� o߁ߓߥ߷�����j� ���#�5�G�Y���}� ��������f����@�1�C�U�g�>�i���>�������������������, ��?&cu\ ������� )M4q�j� ����/�%// I/[/:�/�/�/�/�/ �/���/?!?3?E?W? i?�/�?�?�?�?�?�? v?OO/OAOSOeO�? �O�O�O�O�O�O�O�O _+_=_O_a_s__�_ �_�_�_�_�_�_o'o 9oKo]ooo�oo�o�o �o�o�o�o�o#5G Yk}���� ����1�C�U�g� y��������ӏ��� 	���-�?�Q�c�u��� ��p/��ϟ���� �;�M�_�q������� 6�˯ݯ���%��� I�[�m������2�ǿ ٿ����!�3�¿W� i�{ύϟϱ�@����� ����/߾�S�e�w� �ߛ߭߿�N������ �+�=���a�s��� ���J�������'� 9�K���o��������� ��X�����#5G ��k}�����ڮ��������&�HZ4,F/�>/�� ���	/�-/?/&/ c/J/�/�/�/�/�/�/ �/�/?�/;?"?_?q? X?�?|?�?�?���?O O%O7OIOXmOO�O �O�O�O�OhO�O_!_ 3_E_W_�O{_�_�_�_ �_�_d_�_oo/oAo Soeo�_�o�o�o�o�o �oro+=Oa �o������� ��'�9�K�]�o�� ������ɏۏ�|�� #�5�G�Y�k�}���� ��şן������1� C�U�g�y�������� ӯ���	��?-�?�Q� c�u���������Ͽ� ��Ϧ�;�M�_�q� �ϕ�$Ϲ�������� ߢ�7�I�[�m�ߑ� ��2����������!� ��E�W�i�{���.� ����������/��� S�e�w�������<��� ����+��Oa s����J�� '9�]o� ���F���/�#/5/G/�$UI_�INUSER  ����h!�  H/�L/_MENHIS�T 1yh%�  (w � �(/SOFTP�ART/GENL�INK?curr�ent=menu�page,148�,2�/�/??0?��)�/�/133,1 1??�?�?2?'E?W>71l?�?O#O5O�y+�?W5edit�"?TELEOP�?�O�O�O:O��O�O�O_ _*_<_�O`_r_�_�_ �_�_I_�_�_oo&o 8o�_Iono�o�o�o�o�o��\a�!\o�o /ASVow�� ���`���+� =�O����������� ͏ߏn���'�9�K� ]�쏁�������ɟ۟ j�|��#�5�G�Y�k� ��������ůׯ��o �o�1�C�U�g�y�|� ������ӿ������ -�?�Q�c�uχ�ϫ� ��������ߔ�)�;� M�_�q߃�ߧ߹��� �������7�I�[� m��� �������� ������E�W�i�{� �������������� ��ASew�� �<���+ �Oas���8 ���//'/9/� ]/o/�/�/�/�/F/�/ �/�/?#?5? �2�k? }?�?�?�?�?�/�?�? OO1OCO�?�?yO�O �O�O�O�ObO�O	__ -_?_Q_�Ou_�_�_�_ �_�_^_p_oo)o;o Mo_o�_�o�o�o�o�o �olo%7I[�F?��$UI_P�ANEDATA �1{����q�  	��}  frh/c�gtp/flex�dev.stm?�_width=0�&_height�=10�p�pice�=TP&_lin�es=15&_c�olumns=4��pfont=24�&_page=w�hole�pmI6)�  rim�9�  �pP�b�t������� �����Ǐ��(�:� !�^�E�����{������ܟ�՟�I6� �   2��_dJ�O�a�s��� ������ͯ@���� '�9�K���o���h��� ��ɿۿ¿���#�5� �Y�@�}Ϗ�vϳ�&��Ɠs�����)� ;�Mߠ�q�䯕ߧ߹� ������V��%��I� 0�m��f������ ������!��E�W��� �ύ�����������:� ~�/ASew� �����  =$asZ�~ ����d�v�'/9/ K/]/o/�/��/�/* �/�/�/?#?5?�/Y? @?}?�?v?�?�?�?�? �?O�?1OCO*OgONO �O�/�/�O�O�O	_ _-_�OQ_�/u_�_�_ �_�_�_6_�_o�_)o oMo_oFo�ojo�o�o �o�o�o�o%7�O �Om���� �^_�!�3�E�W�i� {������Ï����� ����A�S�:�w�^� ������џDV�� +�=�O�a�������
� ��ͯ߯���|�9�  �]�o�V���z���ɿ ���Կ�#�
�G�.�k�ޟ�}�|ϵ����������)��4ߧ� #�`�r߄ߖߨߺ�!� ���������8��\� C���y������������������$U�I_POSTYP�E  ��?� 	 �s��B�QUICKME/N  Q�`�v��D�RESTORE� 1|��?  ����!��������mA Sew�,��� ���+=Oa n����� //�9/K/]/o/�/ �/6/�/�/�/�/�/� ??0?�/k?}?�?�? �?V?�?�?�?OO�? COUOgOyO�O6?@O�O �O.O�O	__-_?_Q_ �Ou_�_�_�_�_`_�_ �_oo)o�O6oHoZo �_�o�o�o�o�o�o %7I[�o������SCRE���?��uw1sc��u2�U3�4�5�6��7�8��sTAT�M�� ����:�UGSER�p��rT�p��ks���4��5*��6��7��8��B��NDO_CFG �}Q�����B�PD�E���N�one��v�_IN_FO 2~��)���0%�D���2� s�V�������͟ߟ ��'�9��]�o�R����z��OFFSEOT �Q�-��� hs��p�����G� >�P�}�t���Я��׿ ο����C�:�L�@^Ϩ����͘���
�����av��WORK �!�����.��@ߢ�u�UFRAM�E  ���R�TOL_ABRT8�����ENB�ߣ�?GRP 1�����Cz  A�� ����*�<�N�`�r��֐�U�����?MSK  �)����N��%!��%xz����_EVN��b���+�ׂ3�«�
 h�UE�V��!td:\�event_usger\�u�C7z�d��jpF��n�SPs��x�spotwe{ld��!C6��������!���G |'��5kY�� ���>�� �1�Ug��� /��	/^/M/�/-/ ?/�/c/�/�/�/�/$?��/H?�/:J�W�3�����8C?�?�? �?�?�?�?O+OO OOaO<O�O�OrO�O�O �O�O_�O'_9__]_�o_J_�_�_�_�$V�ALD_CPC {2�« �_�_� w��qd�@R�*o_oqo��hsNbd�j�`��i�da{�o av�_�ooo3BoW i{�o�o�o�o��o �PA�0�e�w� �������� �(�=�L�a�s�
��� ����ʏ�����$� ޟH�:�o��������� ڟ؟����� �2�G� V�k�}�������¯ԯ �����.��R�S� yϋϚ���������� 	��*�<�Q�`�u߇� �ϨϺ��������� &�8�M�\�q���� ����n������"�4� F�[�j��������� �������!0�B�W f�{���������� �,>teT ������� /+/:La/p�/�/ ./�����//'? 6/H/?l/^?�?�?�/ �/�/�/�/?#O�?D? V?kOz?�O�O�?�?�? �?�?_O1_@ORO9_ vOw_�_�_�O�O�O_ �__-o<_N_`_uo�_ �o�o�_�_�_�_o &o;Jo\oq�o�� ��o�o�o� �"7� FXj������� ����!�0�E�T� f�{�������ßҏ� ���
�,�A�P�b��� ��x�����Ο���� �(�*�O�^�p����� ����R�ܯ� ��Ϳ 6�K�Z�l�&ϐ��Ϸ� ��ؿ���"� �2�G� ��h�zϏߞϳ����� ����
��1�@�U�d� v�]�ߛ��������� �,��<�Q�`�r�� ������������� &�;J�_n������ ��������$ F[j|���� ���0E/T i/x��/��/�/�/ �//,/.?P/e?t/ �/�/�?�?�?�?�/? ?(?:?L?NOsO�?�? �O�?�O�OvO OO$O 6O�OZOo_~O�OJ_�O �_�_�_�O_ _F_D_�V[�$VARS_�CONFIG ��Pxa�  FP]S��\lCMR_GRPw 2�xk h�a	`�`  %�1: SC130EF2 *�o�`]TəVU�P�h`�5�_Pa?�  A�@%pp*`�Vn 	No9xCVXdv��a��<uA�%p�q�_R��_R B���#� _Q'��H��l�;��� {�����؏ÏՏ�e� �D�/�A�z�-������ddIA_WORKW �xeܐ�Pf,		�Qxe��>�G�P ���Y�ǑRTSYNCS_ET  xi�xa�-�WINURL 3?=�`������������ȯگSI?ONTMOU9�]S�d� ��_C�FG �S۳�S۵P�`� FR:\��\�DATA\� ��� MC3�L�OG@�   U�D13�EXd�_Q'� B@ ����x�e_ſx�ɿ��VW � n?6  ���VV���l�q  =�C��?�]T<�y�Y�TRAIN���N� 
gp?�CȞ���TK���b�xk (g�����_����� ����U�C�y�g߁���ߝ߯������_GuE��xk�`_P��
�P�RꋰRE���xe*�`hLEXr�xl`1-e��VMPHASE � xec�ecR�TD_FILTE�R 2�xk �u�0����0�B� T�f�x�����VW���� ���� $6HZ�l_iSHIFTM�ENU 1�xk
 <�\%����������= &sJ\��������'/�	�LIVE/SNA��c%vsfli�v��9/��� �7�U�`\"menu r/w//�/�/����Y�]��MO��y�Y�5`h`ZD4�V��_Q<��0��$WA�ITDINEND���a2p6OK  !�i�<���?S�?�9wTIM�����<Gw?M�?*K�?
J�?x
J�?�8RELE���:G6p3���r1_ACCTO 9Hܑ�8_<�7 �ԙ�%�/:_<af�BRDIS�`�N��$XVR���y��$ZABCv�b1�S; ,��
j�I�2B_ZmI1�@VSPT �y�\�eG�
�*�/�o�*!o7o�WDCS?CHG �ԛ(���P\g@�PIPL2�S?i��o�o��o�ZMPCF_G' 1��ii�0'¯S�;Ms�S��i��p�'��g��e2���  �`u������<�"����?`A=�s��=s�=�.9��~|C����B���C�װ�1�q?-W���
M������t<���#�@>b��|�pժ�x�p��p��p{�C� B� �C�I��}���?�Z�~���Ï��y�C0�T�����Gwڂ?���	��ӈ�����*��@�N�x������0 �`��Tp���o�_CYLIND��ݢ { Х� ,(  *=�N�G�`:�w�^����� �� ѯ���7����<�#� 5�r�����������޿ y�_����8�ύ�n�Ȁ�㜻ã wQ �5�����S����Ϡ(�ٻ�X�זr�A���SPHERE 2���ҿ��"� �������P�c�>�P� ̿t���ߪ����� '���]�o�L���p� W�i������������PZZ�F �6