��   ��A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ����CCSCBG�_GRP_T �  $SE�RIES_TYP�E  $PS�_PRM_UPD�A��I OTE$�MODEL_NA�ME :An O�tNSWEIGH�T  $DI�VCONST_F�F �T�SBF�Rq  $�RANGE� ���� ���P_H_�LIM��L�F�SOF� S��M�_INI�DOU� REQ�DIG�I�+��$$C�LASS  ����P��u��u�EVERSION�M  �XKaIRTUAqLM_' 3 n{u�F � WC ���������� B  y %!C�  )%�Bp��?/l/  