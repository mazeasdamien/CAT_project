��  �"�A��*SYST�EM*��V9.4�0107 7/�23/2021 A   ������CCBD_�DATA_T � <$CO�MMENT �$IMCMF_�CF  NE�NDWTWCWFkDBWCd	FGW�TOOL_NUM�W w   qN�~ _FR�w �TRQ��GAIN�$T{DC�$CJI �� T�$DSR`��	I VP�AA�CTL_�TI�$MOV�E_L�WG@D�RARHY& {�/PARM9� �N PEQE} ��K�D&��3�K�K�D_M����3�h�+ �F�STd��|SU�  � L$L�IMIT� �$INSERT_�DIhx$�AM�_F Us"SRBPҎ)P�'|I3/�bBNR x �_d�!B=�'TE0��$b�!ALr�"�AE�'FV��#T�9�v!A2U�(UNJ8V� TVh5Uq8�GRAPH�'RE�TRYS�<1�<2~WEC_DDE&x� �1�7A_PO�0��2AN� �5#��TWL�3ALLT�0�VV'@�!�$VCp27@�2�$�2Ar6@LhP�HD_RA�X`ED�sAheA�GO"�@�� I�DVA_SWG2�@��Ah�@5EhA� LE� �D�MC�ORWPH��!-ASDFW�FY_j"�CP�APz1QTN_S�#�CNGFh$M�IN�@�"?A_ML�_LM�VEL_�CNST�C$AUT_RVbUnPk@3_TL�0TH�1�T��1XSRUDAMP_��O|PS OLSTOP_THRE�1�TAV~Ub �P�D�SRAA�TM�Y��V��QATTOSC_GGDW�E*e#lR�FORCE_O�u MOF\eeI ��LSU�TJUT�fRO�T� C�1� CRE�W~#u �a�eCHG�ZQ�D�dDP@�cV��P��aR�1-AINISH�s�I�`_q�D�a^W�SoT@u|�WZPOCITYjmZP�CNm D�0�Dv�Pdv� �#]#e/w/�/�/�'� 5� ($WO�R� 2�V ' )�2U"�q�ST�P ��pCH�B�rY�#RV^��g�N�Y��FtY�ACTY�C`WA�w��3e�_M���DCPdY�V�e�V�����WQ���^�8��^Q��RTN|ac��T����a�rALGwO_Sxr$P�1��tr�REV_I�T�1�MU�D�0CaCI�!8R��XI��gGAM ![AAS��vє_O@NTR�vYF�`�TR��V�CNPFv�?P�$�.lDCNC0M[ �Z�`O�CHQ�L��Y�F'�l�5�^�OV�M)�QL����IO£�D�A��b���JTH^QPA�V䥽��PDA�pc��DS�PPCCNMONL	S�$�T�1 �T�yV�@J�KPGRC�d�RG�1o��dr�RRo�O�sa�T��O�"_�Rp2�ٽV�-���PDU2CCNAgGWA�g�TH�SǱA-�M�S?ǖS�CVRS1]���a�M۵8a�82�OVK�v���P'���5���VLX����TCI���Y��TRS?`Vo�MG �CCQi��T(�s12��INDEmA�`TM�3P�fT�CC��T�R=G=�USPF8w�p���k@��TWD����f��SR۵��1D��ի����E^PK�PP�Z��CAXCP_P0�B�L��SR���#DI1��?PZH�5��&�RTY��LU�FFIXE�CREAG�Q+u��࿣F�p�q�P+CM�r��CN3FCf��EN� 2����Vѐ��RT�V��TMU��RG`��T����DU%�B�T9�?���Sm��`�P7�`�b�`�IP�)��APf@y���V����Ne�� P�M`����砣���RCh�Pe���7�PS H��(�PYC)���C(L��p�T#_jQ^0�!� EQD=�M�VROU2�PEwRIOF1P��F��2D'���TU�_D���ǔ����T����K�	K��K��CL���*aAD�J�Q_U^Bq�A�aPT�b>�2>REAP�r<�]?Wm 0rq$�DL�W�"�M��M��0�'� ��lB)���'#�*�F#<+(e#�VL��#z*��#�+(8�#z*�P_B���2
�A�-��,� �,�OVER�D�"IB$]PGFQ�L9D L9`���0PCZb�FR~7��@D�@C5P�MN�1�6�q�12�>UF�p�;TOOU@�0_T�1�5N'�H?QcOR��t2p ALs�oG��&�KE�e�&S~��AUXBD�� 4$IMCM�P�r��;� q��@��AUX_AXS�� �{C�p` 	 h�@PEx`���D^c�Cޣ@�C^a�C�X�GDX�z`����fXAXI~@ 
 Td���Db�E�eA~@{@ �pQ�PvR	$�IrX�P�V
�S��G�RN�H $N�1E_U�p��T@�2�Q�05�;��rE����Vk oDON�Q|Va� R_PKG�R�qP  |R`
pQS`�Qb�Qb��P%d`D`%`�$�Ka^�Ƃ`FL~��&pLT �P��ea��c�b��~�a$DYN�E)$J ugG�g	�d���d��	PQCQxP
 ��$Ґ  ����q   &�p &�`:0SIO�Nx  �XKqIRTU�ALq�SCOM� ?&x&� 2 qv|t�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ����
��.�J�Uu�P11w 3c{xp�1pJ���G��� � ���� ?�  ŵ��A  a յ��ĺŹ@@ǻ���
��=�C��� B�߲Cʮ���-χ�xY�����F@ �Ş��=�������Dz  �����υ�C�T`����P�m� "�~�������ǿٿ�� �������E�W�i�{� �ߟ�����������?� �/�A߂�&��⁽�� +�����	���P�
�y�3A���@��Т�h��p��w�BH���Љ�Y���\�  @�� ���#B��?*	���҄і�#�W�v��>��� Qh����pp��H'8[P2K t������� //��7.���A ]/���ݱѕ/3��|� Z��/�/??+6����F7�/�)�r7^	�>��?l�	��N�5>L��?��1N��"U�<#�
q��p�?92�86a"��	����5QB���5@���4��}O l4���F�M��e�B��5:� _!_3__�W_i_|���=��uB�4!??�_�#Itk$ �_$B>��2	
�_gA�$o�_-ox�_�VR0+���ye�.����eQ1$�{���e(4$ܡe�Yokk;��.�e>���H�e�a5�=��e8M�Y�eY-=�0uQ2>"7I [m��w
?o� ������>�P� b�5o��}�����������	ӏ(��L�7� �ow�������ԟ�O ���Y�k�}ߏߡ߳� E_����{���1ﯯ U��y������� �����=�O��s� }�;�M�n�ͯ߯�_� �g�9�K�]�o��ϓ� �������-ߣ��?_� �߃�����������K� %7I�ߑO ��ɿW��b�t��� ����EW���� (:L^p����� A/S/e/w/�/�/�/ �ˏQcu�=?O? a?s?�?/�?�?�?�? �?/O�/9OKO]OoO �/�O�O?�O�O�O�� y?�?�?�?�?�?}_�_ �?�!Og��_�_o/O %O�OIO�oyo�o�o�O �o�o�o�o	-�_ �_�_�_�_o/�4oo XojoQo�ouo�o�o�o �O�o�o'Tf x;����[��[O ��,�>�P�O?���� տ���'�/��?� �?�ߥ���s����� ����+�)�O�a�3� ������ˏݏ����� ɯ7�I�[�m�ۯ��� ��ǟٟ�1��!�3� �ߓߩ�����'�d��� �#�5�c�Y�k�}�� �����N������� 1�ӿU�������&� ����\�n����� ����������� ����;���� �������/����� /��%/7/=�[/m/� �/�/�/�/�/t? !?3?E?W?i?��/ (//L/^/�?O�/�/ �O�eOwO�O�/�/6? �/�O�O__S?=_O_ a_s_�_�_�_2ODOVO hOzO�o/?�O�O�O�O �O
_�O._@_R_%?v_ m__�_�_�_�_��_ oo<o�]o��o�o �o�o�og�y��o�c� u�C��;/q�� ��;�M�_�q��� ������ݿ��# 5GYku�3�y�� �ˏE�����1�C� U�g�U�����_���� ��3�E�W�a�{ύϟ� ����1�������/� A�ʿi�w߉ߛ߭�O� ��Z�l�~ϐ�+��O� ������� �2�D�V� h�z��'�9�K�]��� ���������7�I�v� m�#5#�Yk�� ������ 1CUg����� ͯ��_q�-/� ��u/�/y�A?C �/#?��E_? q?�?�?/�?�?�?�? OO%O�/�/�/�/�/ _?,??P?7?t?�? m?�?�?�?��?�?�? OOLO^O!o�OmOO �OSo�Owo __$_6_ H_�o�o��������� �w�_�_ oo����� o��ɟ۟ퟣ_�go 5�/�Y�{_Mo�_�_�_ �_�o��./oAoG �wo�o�o�o�oE�'� �og�y������ ��J����	��-�?� ��c�u�W�������܏ U�j��Ϲ�;ϒ�֯ �����Ϲ�+�T�f� x���������ҿ��� �ߣߵ��������� ��7O-O�������ϟ� ��7�����p���/� A�S�e�w��������� ��k�}�+m�O �������2�D�V� ����Ϟ���O]�� �
��=��� /G5/G/Y/k/}/ *<N`r�?� }����� /&/ 8/J/S/�/w/�/�/ �/�/�O�/�/"??��U?�O|?�?�?�?�=��$CCSCH_G�RP12 3�����1&� x��o_5 �Yk^O�!��O�O �O����O1���U� g�y���_����ӏO �OZ_LObOpOz_8oJo ko�O�O�O\o_$_6_ H_�_�o�o�_�_�_� �:�)�;��xoq� ����SϹ�H�ݟ� �%�7���[���� T��_�q�������!� 3�ɟ���%�7�I� [�m�����o�/�֯ \�e�{ω�0�ҏ�/i� `�r����+�6�O�a� υߗߩ߻������� ���'�9�K��䏁� ������H�vߜ��� ������Y�k�����9� 7a?������>��F� ��Ugy���� ���	�������� ��/1AgN �r������ $Qcu?� ���.��//)/ ;/M/��?_/�_�_�_ oo,o��??��o �o�o(?�o �o (~?LF�p�/d?�/ �/�O�/�?�O�O�OF? X?j?�O�?�?�?�?�? �?._OO0O~p/�_ oJ��ao�� �2� `�V��oz������� Xo
�����BO�_R� ����#���ПY� k�}�������ŏ׏� ��:_��̯ޯ�� ��&�8��Dʟܟ� ���ȿڿ�����"� 4�F�X�jϋ������ ������q�0�߄�B� T�f�,o��%��I� [����h�����b� t��Ϟ�3���4��� ��L�:�L�^�p��� ����/�A�S�e�w�� ������������� +�=�O�"�s�j�|��� ��������� 9 �Z�ρ���� ȿv/�NO`OrO���O �O:π>�po�� �J_\_n_�_�_�_� �_�_� 2DV hr/0?B?���� T?
/\/./@/R/d/�? �/�/�/�_o"O0oBo �O�Oxo�o�o�o�o�o �o�o,>�_b t�_��LO�Woio {o�o�o:�L��o�o�o /ASew� $�6�H�Z�p�~����/ ��=�4�F�s�j��2� �V�h�z�o�����O ԯ�o�
���.�@�R� d�퟈�������п� �On�������ůׯr� ����>�l����� l����>�\�n߀ߒ� ̿�����������"� �Ͻ����������)� �M�4�]߃�jߧ߹� �ߞ�������%��I� [�F<��|��P�� t���!�3�E��� P��?�/�/��?���� ��{�l?~?���?�? �?�?�?�t2O,oVO +������������� ��,>D�/� ������ �vO�O?�O�O�� �O__*_X_�?`_r_ �_�_�_�_CO�_�_o o&o�/Jo�O�O�O	_ �o_�oQ_c_u_�_�_ �_�_�_�_�_��� ��\o��~0��_ �o�o�o�o�����oҏ ���,�>�P�b� t���������Ο��i� ��(�F?L�^�؏� ��� �A�S�� ��o ������Z���~���� ���ؿ���ϔ�2� D�V�h�zϐϞ�'�9� K�]�o��ߓ�����ɿ ������#�5�G�� P�i�tφϘ����Ϛ� ������1���R���y� �ߝ߯���\�n�4/ x/j<���f�x�� ��/��0/B/T/f/ �/��/�O�/���� �*�<�N�h�(�� �����:����&� 8���n������/�/ ~(?:?�Vp?�? �?�?�?&/�?�?�O $O6OU�/�/~O�O2 �O?O?a?s?�? _2_ �?�?�?�?OO'O9O KO]OoO
oo.oDoRo dozo�o_�Ϧ�G_>_ P_i_*�_N`�_ �������� �&�8�J��_�_���� ���oȏ�T*�j ���j�x_n_�6� `�֟_�����z�$��� T�f�x���������ү ���|�������ǟٟ �
�����E�,�i� P�y�����ï��̯�� ��/�A�S��w�b� �����οl������+�<��$CCSC�H_GRP13 �3���^��&� x n�߮�������� ���4�bt�%� �����{�( "?L��a��������� �߱�����C�U�g��� �ߝ߯���g�Y�+�	� �-�Zl���� ^����/�O2/� V/h/�/�/�/.�/ ~�/���.?��� / /�?�?B/h/z/�/ �/�/�/�/�/�/
?� �O�OO?��O�O_�? K ��?�?�?O�_�_ �?�_�_�O�_o"o4o FoXojo�O�o�o�o�o _]�o0B�_ �_O"ooFoXo�� O	O�o��ڿP��ot� �o�oQΏ���� �(�:�L�^�p���,� >�P�b�t��������� ����Ǐ��(�:�L� ;%�g�������ʟܟ ����6�!��i� ~�������Ư}_s�د K�]�o����7o}� ��m���#���G��� k�}������������ �ݿ/�A��e�o�-� ?�`߿�ѿ�Q��Y� +�=�O�aϧ߅ϗϩ� ������OQ��u �����=�� );��_q��� ��I��Tfx�� 7/I/���, >Pbt��}�3?E? W?i?{?/�?�?��� C/U/g/�//OAOSOeO wO ?�O�O�O�O�O? _�?+_=_O_a_�?�_ �_�?�_�_�_��kO�O �O�O�O�Ooo�o�O�/ _Y��o�o�o!__�_ ;_�k}��_�� ������o�o�o �o�o!�&J\ C�g����_� ����F�X�j�-� ��y���M�ӏM_��� �0�B�AO�x����� ��/�!߳O���O�� ����e��������� ���A�S�%����� ����ϟ�믩���)� ;�M�_�Ϳ��կ���� ˯ݯ#���%�s�� �ϩ���V����� '�U�K�]�o������� ��@�����v�#�� G���������� N�`�r����������� ���������� �	/w�-/���� ��?�/��/�/�/�� ?)?/�M?_?��? �?�?�?�?f/OO%O 7OIO[O��/??�/ >?P?�O�O�?}?�_� W_i_{_�?�?(O�?�_ �_�_oEO/oAoSoeo wo�o�o$_6_H_Z_l_ �!O�_�_�_�_�_�_ �_ o2oDoOho_oqo �o�o�o�o���o
�o .ɏO�v��� �Y�k���U�g�5 ��-?c�u������ ��-�?�Q�c�u��� �ϥ��Ϥ���'�9� K�]�g�%�k������� 7������#�5�G�Y� G�}���Q����{�%� 7�I�S�m�ߑߣ��� #��������!�3�� [�i�{���A���L� ^�p߂����A����� �� ��$�6�H�Z�l� +=O��s� ���w�)�;�h�_� '�K]����� �����/#/5/ G/Y/�}/�/�/���/ �/Qc�?y�� g?y?k��3O5/�?/ �?�//�/7/QOcOuO �O?�O�O�O�O�O	_ _�?�?�?�?�?oO OOBO)OfOxO_O�O �O�O�/�O�O�O�O_ >_P_t___q_�_E �_i�_oo(o:o� �����㟵��i �o�oa�s����� ��ͯ߯�o�Y'�!� K�mo?�o�o�o�o� ���� �!39���i {���7���� �Y�k���������<� Ϗ�����1ϟ�U� g�I��ϝϯ�ΟG�\� ��	߫�-߄�ȿڿ� ���߫��F�X�j�|� �Ϡϲ������σ�� ������������)_ _�߷����ߑ���)� ����b���!3E Wi{����]� o��_�A��� �� ��$6H��� �ߐ�/�_O/�s/� ��/�/�/�/?9 '?9?K?]?o?�
// ./@/R/d/�O�/o/�/ �/�/�/�/�/?*?<? E?r?i?{?�?�?�? �_�?�?O�?�GO�_�nO�O�O�O�M�$C�CSCH_GRP�14 3�����A&� x�ao'���K� ]�P_��z_�_�_ۏ ����_#�u�G�Y�k� }��_����ş_�_Lo >_T_b_lo*<]�_ �_�_Noo(o:o�o ���o�o�oӟ�,� ���-�׏jc�u��� E߫�:�ϯᯋ��� )���M���q��F��� Q�c�u������%ϻ� ����)�;�M�_� q���z�!�ȿN�W� m�{�"�ğ�?[�R�d� ����(�A�S���w� ���������r�� �+�=���֟s����� ����:�h�ϛ�~�� ��K]�ς�+�)SO �s��0���8���G Yk}����� �������� �/#
3Y@}d �������// /C/U/g/	O�/v/�/ �/ �/�/	??-??? ���OQ?�o�o�o�o ���?O�x�� O������pO >�8�b��?VO�?�?|_ �?�O�_�_�_8OJO\O �_�O�O�O�O�O�O o �O_"_p�b?�o<� ʏS� ��$�R�H� �l�~�������J�� �s��4_�oD�͏ߏ �����¯K�]�o� ��������ɟ۟�,/ �_����п���z�� *���6/��ί���� ��������y��&�8� J�\�}���	Ϥ߶��� ��c�"��v�4�F�X� ������;�M��� ��Z������/T�f�x� �ߐ�%��&���� >�,>Pbt�� !�3�E�W�i�{���� ������������/ A�e\n��� ���/�+�/L ��s������h? �@_R_d_���_�_,� r/0�b�
/�/�/<o No`oro�o�o�/�o�o �/ //$/6/H/Z/d? "O4O�/�/�/�/FO�/ N? ?2?D?V?�Oz?�? �?�o�o_"4�_�_ j|������ ���0��oT�f��o ����>_��I[m �,�>������ !�3�E�W�i���(� :�L�b�p����?��/� &�8�e�\��$��H� Z�l������_ƿؿ a����� �2�D�V�߯ zόϞϰ����ϊ_`� ����v���ɿd�v��� ��0�^������^�� ��0�N�`�r��Ϩ� �����������߯� ����������?� &�O�u�\����� ��������;�M�8 .���n���B��f�� %7��B|O �?�?��O����m ^OpO� �O�O�O�O �O�f$_H_/| �������/� 06/�/
?x�� ����/�/�/h_ z_�?�_�_�/�/�_�_ 
ooJo�ORodovo�o �o�o5_�o�o�o �?<�_�_�_�_�o �CoUogoyo�o�o�o �o�o�o��������ȏ N���p/"��o�� �������ğ֟� ����0�B�T�f�x� ��������ү[���� �8O>�P�ʟܟ���� �3�E����r��� ��Lώ�p�������� ������ ߆�$�6�H� Z�l߂ߐ��+�=�O� aπ�ϗ�~ϻϢ��� �����'�9��B�[� f�xߊ߷��ߌ����� ��#��D���k�}�� ���N`&/�/j?\/ .��/�X�j����/�/ �/|�"?4?F?X?�|? ���?�_�?���
�� .�@�Z����� �,����*� �`r��?�?
/p/ O,O�/HbOtO�O�O �O?�O�O�/__(_ G/�?�?p_�_$/�_�? AOSOeOwOo$o�O�O �O�O�O__+_=_O_ a_�o 6DVl z o�ߘ�9o0oBo[o 
���o@�R��ov��� ������Џ���� *�<��o�or������ ���/F��y�\����� ��\�jo`o	�(�R�ȯ Q��u�l����F�X� j�|�������Ŀֿ� n���������˯ݯ�� ����7��[�B�k� �������������� !�3�E��i�Tύ�x� ����^�������.���$CCSCH_�GRP15 3����P�?&� x`/�� �r��������� �&�Tfx�� ����m�/O>/ ��S����������� ����5�G�Y���}�� ���Y�K���� L/^/��/�/P�� �/�/ ?�_$?�H?Z? /~?�?�? ��?p/�? {/� O�/�/�/ ?? �O�O4?Z?l?~?�?�? �?�?�?�?�?���_�_ AO��_�_�_�O=/� �O�O�O
_�o�o�O�o �ov_�o&8J \�_����oO/ ���"�4��o�o_ �o8Jď֏_�O �����B��f��� �C���ҟ����� ,�>�P�b�t��0�B� T�f�x�v�������ҟ ����ݟ�,�>�-�� Y���}�����ίூ� ��(����[�p��� ������ooe�ʿ=�O� a�s�����)oρ�_ ����9�]o ���Ϸ�/����� !�3���W�a��1�R� ������C���K��/� A�Sߙ�w߉ߛ��ۿ ����_C��gy� ���/��	// -/��uoc/��/��;� �/FXj|�)?;? ����//0/B/ T/f/��o�%O7OIO[O mO�/�O�Ox/��5?G? Y?�?!_3_E_W_i_�? �_�_�_�_�_�?�_�O o/oAoSo�O�o�o�O �o�o�o��]_~_�_s_ �_�_as�_w?oK� ���o	o�o-o�� ]�o����o����ɏۏ ��������� ����<�N�5�r� Y��������oޏՏ�  ��8�J�\����k� ��?�ş?o����"� 4�3_�j�������? ��_믩_���/�� ��W������������ �3�E��y������� ��ӯݿ�ϭ��-�?� Q���u�ǿ������Ͽ ����e�w��ߛ� ���H�����G =Oas���2� ��h���9�� ������
��@R dv������ }/�/�/�/�/�/�/�/ i�?������O �?��?�?�?��	OO !�?OQO�/uO/�O�O �O�OX?�O__)_;_ M_��?�?O�?0OBO �_�_xOoO�oןIo[o mo�O�O_�O�o�o�o �o7_!3EWi{ �o(o:oLo^o}�_ �o{o�o�o�o�o�o $6	_ZQc�� ������� ��� A�ߟh�z�������K� ]�����G�Y�'/}�O U�g��������y�� 1�C�U�g���ߟ�ߗ� �ߖ�����+�=�O� Y��]�������)��� ���'�9�K�9�o� ��C�����m��)�;� E�_�q�������� ������%���M�[� m����3ϵ�>�P�b� t���3�������� ��(�:�L�^�� /A��ew鯛 i�-ZQ// =/O/ws/�/�/�/�/ �/�/�/??'?9?K? �o?�?�?�Ϸ?�?C/ U/v/Ok/�/�/YOkO ]�/%_'?�O?�Or? ?{?)?C_U_g_y_�? �_�_�_�_�_�_	o�O �O�O�O�O�o�O_�O 4__X_j_Q_�_�_�_ �?�_�_�_�_o0oBo �foQoco�o7��o[� �o�o,Ǐُ�� q��կ���[/�� �S�e�w�������� ѿ���K���=�_ 1�����ӏ���� ��%�+���[�m�� ����)��ُ���K� ]σ�鯓ϥ�.����� �����#ߑ�G�Y�;� }ߏߡ���9�N����� ���vϺ������ϋ� ���8�J�\�n߀ߒ� �߶�����u������� ��������y�oo�� ��������� T��%7I[ m���O�a�� �/Q3/����� �(:�/���� �?�oA?�e?��� !/�?�?�?�?+/O+O =OOOaO�/�/? ?2? D?V?u_z?a?s?�?�? �?�?�?
OO.O/7O dO[OmO�O�O�O�o�O �O_�Os/9_�o`_r_��_�_�]�$CCS�CH_GRP16 3����Q�&� xٯS��=�O�Bo s�lo~o�o͟ߟ� �o�g�9�K�]�o��o ���Ϸ��_�o>0oFo To^�.�O��o�o�o @��o,�ď�� t��ůׯ���� �ɟ\�U�g�y�7 ,���ӿ}���	�ϙ ?��c���8���C�U� g�y����߭�ӿ� ��	��-�?�Q�c�u� l����@�I�_�m� ߶��OM�D�V߃��� ��3�E���i�{��� ��������d��� /��ȯew��� ,�Z��ߍ�p�����= O~�t�/E_�e �"�*�9/K/]/ o/�/�/�/�/�/�/�/ �������?/ �%/K/2/o/V/�/�/ �/��/�/�/�/?5? G?Y?�O}?h?�?�? �?�?�?OO1O���_ CO�������� �O�O؟j�|���_�� �֏����b_0�*� T�vOH_�O�Ono�O�_ �o�o�o*_<_N_�or_ �_�_�_�_�_�_o ob�TO� �.？E� �����D�:���^� p�������<���ܯe�  �&o�6���џ��� �����=�O�a�s��� ������ͯ߯?�o�� ��������l�
��� (?����ҿ���߬߾� ����k���*�<�N� o�r��ϖ�����U� ��h�&�8�J���� ��	���-�?�����L� �~��?FXj��� ������0� 0BTfx�% 7I[m�/�x� ����!3� WN`y���� �?��/�?>/��e/ w/�/�/�/��ZO�/2o DoVo��zo�o�d?"� T���/v?�?.@R dv��?���?�/ ??(?:?L?VO_&_ �?�?�?�?8_�?@OO $O6OHO�_lO~O�O� �o�&��o�o\�n� ��������ȏڏ��� �"��F�X��|��� 0o��;�M�_�q���� 0���ˏݏ���%� 7�I�[�����,�>� T�b�t��O��!��*� W�N� �� �:�L�^�  ��ϔϚo����S��� |��$�6�H�ѿl�~� �ߢߴ���|oR�sυ� hϩϻ�V�h�����"� P/������P��ϓ�"� @�R�d�v��ߚ����� ������������ ��������1��A� g�N������������� ��	 -?*/ u `�4/�X/�� )�/�/4n_�O�O ���O����_P_b_ x��_�_�_�_�_v/ X/o�:o?n�� ����/�?�//"/ (?�?�?j/|/�/�/�/ �/�?�/�/�?Zolo�O �o�o�?�?�o�o�o <�_DVhz�� 'o����
��O.� �o�o�o�o���o��5 GYk}���� �r���������@�ޟ �b?������ӏʏ ��������ȯ����� �"�4�F�X�j�|��� ����ĿM�����*_ 0�Bϼ�ί﯊��%� 7�����֏d��ߠ�>� ��b��z��������� ����x��(�:�L�^� t����/�A�S�r� w߉�p߭ߔ������� ��+���4�M�X�j� |���~������� �6��]�o������� @R?�?\ON? �r? ԯJ\}�?�?�?n O&O8OJO nO��O �o�O����� 2 L�/����/ ���
�/�/R dv�O�O�/b?__ �?:/T_f_x_�_�_
O �_�_�?�_oo9?�O �Oboto?�o�O3_E_ W_i_�_�_�_�_ �_�_oo/oAoSo�  ��(�6�H�^�l��o ���+"4M��� �2�D��h�z����� ��ԟ���
��.� ��d�v���ʏ��r? 8��k�N�������N� \R���D���C�޿ g�^����8�J�\�n� ���Ϥ϶�����`�u� ��������Ͽ���ڿ �)��M�4�]σϕ� ��z����������%� 7���[�F��j�쯲��P�������� ��$�CCSCH_GR�P17 3����B�&� xR?���d/ �����~������ F/X/j/	��/�/�/�/ �/�/_�?_0?s�E� ������������ '�9�K��o������� K=����>?P? ���?�?B/��?�? �?�oO�/:OLO�/pO �O�O��Ob?�Om?� _�?�?�?�?O~_�_ &OLO^OpO�O�O�O�O �O�O�O�zo�o3_�/ �o�o�o�_/?��_�_ �_�_v��_��ho ����*�<�N��o r��������oA?ޏ�� ��&����_�� *�<���ȟ�_�_���� ��4�ޏX�������5� ��į֯�����0� B�T�f��"�4�F�X� j�hώ�u���į��� ϯ��0��	�K�x� o�������ҿt���� �ϋ�M�b�tφϘ� ��aW��/ASe w��a�s�Q/�� ��+}Oas� �ߩ�?������%� ��I�S��#�D��ߵ� ��5���=��!�3�E� ��i�{�����y �o5/�Y/k/}/�/�/ �/!�/�/�/??� gU?�y?��-�?8/ J/\/n/�/O-O�/�/ �/�/�/?"?4?F?X? ��a�_)_;_M___�? �_�_j?��'O9OKOxO o%o7oIo[o�Oo�o �o�o�o�O�ot_! 3E�_�{�_�� ��Oopo�oeo�o�o S�e��oiO�o=Ͽ�я ��o���O�a� s��������͟ߟ� �������ԏ�� 
��.�@�'�d�K��� ����Пǟٟ��� *�<�N��r�]���1� ��1ޯ���&�%o ��\�������?��� �oݿ�o�{?u��I� ������������% 7	�k�}�������ſ �ύߟ���1�Cϱ� gϹϋϝϯ������ ��	�Wi���� :����9/A Sew��$�� Z�/��+/��� ���/�/2DVh z�����o?�? �?�?�?�?�?�?[�O �/�/�/�/�/y_�Oy/ �O�O�Oy�O_�1_ C_�?g_�/�_�_�_�_ JO�_�_	oo-o?o�� �O�O�O�O"_4_�o�o j_a_�ɯ;M_�_ w_o�_����)o �%�7�I�[�m�� ,>Po�o�m �������(� �_L�C�U���y����� �����ُ���3�ѯ Z�l�~�����=�O��� ��9�K�?o�_G�Y� ؟�����k��#�5� G�Y��ѯ��� �����/�A�K�	� O��������u���� ��+�=�+�a�s�5� ����_�	��-�7�Q� c�u����������� ����?M_q �%ߧ0�B�T�f� v�%���������� ,>P��/!/ 3/�W/i/ۿ�/[ LC�/?�/?A? ie?w?�?�?�?�?�? �?�?OO+O=O�/aO sO�O�ߩO�O5?G?h? _]?�?�?K_]_O�? oO�_�?�_dO�?mO O5oGoYoko�O�o�o �o�o�o�o�o�_�_�_ �_�_��_o�_&oo Jo\oCo�o�o�owO�o �o�o�o�o"4��X CU�)��M��� �����˟��c��� ǿ��M?ÏՏ��E� W�i�珍ϟϱ���y� ��=���/�Q�#�u� ������şs����� ����M�_�q����� ���˟ݟ�=�O�u� ۿ�ߗ� ϳ������� ���9�K�-�o�� �ﲿ+�@����� h߬߾�����}���� *�<�N�`�r���� ����gy���� ��k������� ��u���F� �//)/;/M/_/q/ �/�/�/AS�/�/? C%?뿱���/ /,/�?����t/�O� 3O�/WO�/�/�/?�O �O�O�O?__/_A_ S_�?�? OO$O6OHO golOSOeO�O�O�O�O �O�O_ _�/)_V_M_ __�_�_�_s�_�_�_ �_e?+o�Rodovo�o��m�$CCSCH�_GRP18 3�����a&� x˿ E��ݯ/�A�4e�� ^p���ѯ㯂� Y�+�=�O�a����� ���o�0�"8FP� � �A����2�� ���ď����f�x� ����ɿ�v���ϻ� N�G�Y�k�)������ ��o�����ߋ1�ۿ U��*���5�G�Y�k� }���	���������� ��1�C�U�g�^��� ���2�;�Q�_�憎 }_?�6�H�u���� %7��[m�� ��V���!v� ��Wi{��L r�b��//A/p� f�?7o�/W�/ r�+?=?O?a?s? �?�?�?�?�?�?�/�/ �/�/�/�/�O?�/? =?$?a?H?�?�?�?� �?�?�?�?�?'O9OKO �_oOZO�O~O/�O�O �O�O_#_���o5_�� ��̏ޏ�����_�_ ʯ\�n����_����ȟ ڟ���To"��F�h_ :o�_�_`�_�o�� �o.o@o�do�o�o �o�o�o��o�oT� F_|�� ���7�ү� ���6�,���P�b�t� ����.���οW�� ��(ϱ�ïկ����� ��/�A�S�e�w����� ����ѿO��ߢߴ� ����^�����O�� �����ό������� ]���
��.�@�a�d� �߈�������G��� Z�*<������� ���1���>���p� �O8J\~�t�	�� 
/���"/"/4/ F/X/j/|/); M_~?�j��� ��//%/��I/@/ R/k/v/�/�/�/�O�/ �/?�O0?��W?i?{? �?�?��L_�?$6H v�l~�VO�F��� �?hO�O �2�D�V�h� z�xO�����O�?�?O O,O>OH_oo�O�O �O�O*o�O2___(_ :_�o^_p_�_Џ��o ��v�N�`�r��� ������̟ޟ��� ��8�J�ӏn���"�� -�?�Q�c�u��"��� ��ϟ����)�;� M������0�F�T� f��_���
��I�@� ����,�>�P��t� �ߌ�߼�E���n�� �(�:���^�p��� ���nD�e�w�Zߛ� ��H�Z�����B?�� ����B��߅��2D Vh������ ������������� ~�����#
3Y@ }��t����� �1?gR� &?�J?���	// �?�?&/`o�_�_���_ ���/�/Q/BoToj/�/ �o�o�o�o�oh?J? �,O`/r/�/�/�/ �/�?�O�???O�O �O\?n?�?�?�?�?�O �?�?�OL^�_�� �O�O��� �.��o 6�H�Z�l�~����� Ə؏����_ ��� ��z����'�9�K� ]�o���������ɏd� v�������2�Я�TO �ԏ����ş��r��� r������޿��� &�8�J�\�nπϒϤ� ��?�������o"�4� �����|�ֿ�)��� ��ȟVϐ��0�r�T� ��l��ϔϮ������� j���,�>�P�f�t� ���!�3�E�di�{� b����������� ���&�?�J�\�n��� ��p�������( �Oas��2/D/ 
O�ON_@O�dOƿ< No�O�O�O`__ *_<_�`_��_~�_ ��� $>/�/ �/}/~��/?�� ��/�?v?D/V/h/ �_�_�?TO�_o�O,? FoXojo|o�o�O�o�o �O�o�o+O�_�_T fO��_%o7oIo[o ��zo�o�o�o�o�o �o!3E���� �(�:�P�^����|� ��&�?�� ���$� 6���Z�l�~������� Ưد���� ���̏ V�h�z�����dO*� � ]�@�������@�N�D� ��6��5���Y�P� ����*�<�N�`ߖ��� �ߨߺ���R�g�yϋ� �ϯ������������ �?�&�O�u߇ߙ�l� ����������)��� M�8�q�\�޿��B����������$CC�SCH_GRP1�9 3����4�&� xDO��/V?�/�/ ���/p�����
8?J? \?���?�?�?�?�?�? Q�?�_"Oe�7��� ��������+ =�as��=// /��0OBO�/�/ xO�O4?��O�O�O� _�?,_>_�?b_t_�_ ��_TO�__O�/o�O �O�O�O�Opo�o_>_ P_b_t_�_�_�_�_�_ �_�l~%o�?�� �o!O�߸o�o�o�o h�z��o����Zԏ� ��
��.�@��d�v� �����3OП���� ���ŏ�o��ۏ�.� �����o�o������&� ПJ���럕�'����� ȿڿ����"�4�F� X���&�8�J�\�Z� ��g�������ڿ���� �"����=�j�a�s� �ϲ���f�������� }�?�T�f�xߊߜ�S� I���!3EWi{ �S�e�C?���w� /o/A/S/e/w/��/ �O�/�߳�����;� E�6����' ��/���%�7�}[� m���/���k�'? �K?]?o?�?�?�?/ �?�?�?�?O�Y�GO �/kO���O*?<?N? `?r?__�?�?�?�? �?OO&O8OJO��S 	oo-o?oQo�Ouo�o \O��_+_=_j_ );M�_q��� ��_�fo��%�7� �o�m��o������{ AbtW��E�W� �[_�/߱�ß՟� ������A�S�e��� ��������ѯ���~� ������Ɵ؟�����  �2��V�=�z����� q�¯��˯���.� @��d�O���#ߩ�#� п�������N� �������O������� ��mOg���;ߙ� ������)�� ]�oρϓϥϷ���� �����#�5ߣ�Y߫� }ߏߡ߳��������� I[q����,� ���+/!/3/E/W/ i/{/�/�/�/L�/ �/��?����� �?�?$/6/H/Z/l/~/ �/�/�/�/aOsO�O�O �O�O�O�OM�_�?�? �?�?�?ko�_k?�_�_ �_k�_�_#o5o�O Yo�?}o�o�o�o<_�o �o�o1���_�_ �_�_o&o��\oSo ����-�?�Q��oio�o �o����Ϗ��� )�;�M�_�q���� 0�B�a��ox�_����� ��ҏ�������o>� 5�G�t�k��������� ��˟���%�ÿL�^� p�����/�Aϟ���+� =�Oa�o9�K�ʯ�� ���]���'�9�K� �ÿ��{��z�ٯ� ���!�3�=���A�{� �����g�տ���� �/��S�e�'����� Q����)�CUg y������� 	��1?Qcu� �"4FX�h/ ������ 0B�/�/??%?� I?[?��?M�/>/ 5/�?�?�!O3O[/WO iO{O�O�O�O�O�O�O �O__/_�?S_e_w_ ��_�_'O9OZO�_OO �O�O=oOoA/�O	_ �o�O�oV_�O___' 9K]�_���� ���vo�o�o�o�o ݏ�o�o�o�o<N 5r��i_��� ���&��J�5�G� �����?�ȏڏ��� �������U��߹ϋ/ ��?O��ǟ�7�I�[� ٟߑߣߵ�k���/� ����!�C��g�y��� ����e�w�����	�� ��?�Q�c�u����� ��ϯ�/�A�g���w� ��ߥ���������� u�+�=��a�s����� �2�������Z�� ������o����.� @�R�d�v��������� Yk}����� ]������g/ y/��/�/8�/�/�/ 	??-???Q?c?u?�? �?3E�?�?�?5/O �ϣ/y/�/�/�/?? �O��f?�_��%_�? I_�?�?s?O�_�_�_ �_O�_o!o3oEo�O �O�O__(_:_Y^_ E_W_�_{_�_�_�_�_  oo�?oHo?oQo~o �o�oe��o�o�o�oWO���DVhz�}��$CCSCH_G�RP1A 3�����q&� x��7��� Ͽ!�3�&�W��/P�b� ����ÿտt���K�� /�A�S�ʏw�q��� ��"��*�8�B� �� 3�������$�ڏ��� �����z�X�j�|��� ���h���߭�@�9� K�]���ϥ߷�a� ������}/#���G��� �}�'�9�K�]�o��� ��߷���������� #�5�G�Y�P������� $�-CQ���oo1� (�:�g�����) ��M_q���� H��//h��I/ [/m//�/>d�q T��!?3?b�X�/ �?)�?I/�?/d// �/O/OAOSOeOwO�O �O�O�O�O{?�?�?�? �?�?�_�?�?	O/OO SO:OwO�O�O�/tO�O �O�O�O_+_=_�oa_ L_�_p_�/�_�_�_�_ oo��'o������ П�����o�o��N� `�r��o��诺�̯ޯ �F��8�Zo,~o �oR��o�|�����  2��V�z�� ������F�8on� ���)�Ŀֿ��� (�ό�B�T�f�xϊ�  ����I���
���� ����ǿٿ뿆ߘ�!� 3�E�W�i�{ύϟϱ� ��_̏������� P��� ���_�ߤ߶� ��~���������O��� �� 2S�V��z ���9���L�
 .���������� #��0��b�_*/ </N/pf���/�/ �/�/??&?8?J? \?n?�	//-/?/Q/ pOu/\/�/�/�/�/�/ �/??�;?2?D?]? h?�?�?�?|_�?�?O �_"O�IO[OmOO�O ��>o�O�(�:�h�^� p�H_8����OZ_ �_�$�6�H�Z�l�j_ ����t_�O�O�O__ 0_:o�o
x_�_�_�_ �_$o�_oo,or Pobotoԟ���
� h���@�R�d�v����� ����Я������*� <�ş`�r�����1� C�U�g��ϝ����� ӯ���	��-�?��� �����"�8�F�X��o |�����;�2����� ��0�B��f�x�~� ���7���`����� ,���P�b�t������� `�6�W�i�L���: L����4O��� 4���w��$6HZ ��~������ s�����/p�� ��%K2o� �f������/ #/O/Y/D/}/O�/ <O�/�/�/�/?�O�O ?R�o�o���o|�? �?C?4F\?�?|� ���ZO<O���� �OR?d?v?�?�?�?�O t_�O�?O_�_�_NO `OrO�O�O�O�_�O�O �_>�P��ot����_�_ ��Ώ��� �r(�:� L�^�p��������ʟ ܟo�������я l�Ꮠ��+�=�O�a� s���������V�h�z� ����$�¿ԿF_��Ɵ x�������d�v�d��� ��ԯ��������*� <�N�`�r߄ߖߨ�1� �������&�ϲ� ��n���	�߶��ﺯ H߂���"�d�F���^� �߆ߠ�������\��� 0BXf��� �%�7�V[�m�T��� x������������� 1<N`��b/ �����/�/A Sew�$?6?�O�_ @o2_�V_��./@/a/ �_�_�_R/�_
oo.o �Ro�/vop��o��/ ��//0?�?�?o? p/�/�?O�/�/�/�/  ?�OhO6?H?Z?�o�o �OF_�o�_O8J \n��_���_� ��_�o�oF�X��O |��o);M��� l������� �%�7�ҟ����� ,�B�P�֏xn�� �1���x��(��� L�^�p���������ʿ ܿ� �Ϭ���H�Z� lϮ���V_��O�2� s�����2�@�6�߿�� (��'���K�B��~� �.�@�R��v��� ���D�Y�k�}ߏߡ� �����߾������1� �A�g�y��^ϔ��� ������	���?�*� c�N��ϖ�4����������$CCSC�H_GRP1B �3���&�&� x 6_�v?HO�?�?��? b����*O<ONO� rO�O�O�O�O�OC�O �o_W)���� �y/�/�//�/ Sew�//!?�/� ��"_4_{?�?j_|_ &O�/�_�_�_���_�O o0o�OTofoxo���o F_�oQ_�?�o�_�_�_ �_�_bt
o0oBoTo foxo�o�o�o�o�o�/ ^�p��O����ʏq _�����Z�l� w����L�Ɵ؟��� � �2���V�h�z��� �%_¯ԯ���
��� ����͟� ����� ��z�xϢ��¯<� �ݯ����ϨϺ��� ������&�8�J��� ��*�<�N�L�r�Y� �ϨϏ��ϳ����� ���/�\�S�eߒߤ� ��X���������o�1�F�X�j�|��C #5G/�/Q?C/� g/ɟ`�r����/�/�/ ��	??-???�c?�� �?�_�?�����$�6� H�b"������ 4���� 2�� hz��?�?/x/O O�/PIO[OmOO�O  ?�O�O�/�O�O_O/ �?�?W_i_,/�_OIO [OmOO�_o�O�O�O �O�O_!_3_E_W_i_ �o�o+=Sa o���Ao8oJoco� ��o'�9��o]�o��� ������ɏۏ���� #��o�oY�k�}���� �/N�$���d�����ɏ C�roho��9ﯯY� ӯ}�t����-�?�Q� c�����������Ͽv� ��������ӯ���	� ��?�&�c�J�s��� ������ƿ����)� ;�M���q�\ϕπ�� ��E�����%ߟ��D������x�� �o b����,�Zl ~������� s� /OD/��Y�߽� ���������:�;�M� S����������Q 3��%�R/d/� �/�/V���/�/?? *?�N?`?c�?�?�? �a/v/�?O�&O�/ �/�/??�O�O7?`? r?�?�?�?�?�?�?�? O|_�_�_�_�_�_�_ �_�O"���O�O�O�O �o�oC_�o�o|_�o ,>Pbt�� ��w_�_���yo :�!�o�o�o>P b܏__�����H� �l����I�Ɵ؟ ���S� �2�D�V�h� �$�6�H�Z�l�~�|� ������؟������ 2�D�V�)�_������� ¯ԯ毈�
���.�� ��a��ψ�������8�J�EU�g�y�?�� u�G_���o�Ϥ����� ��;M_qH� �߹�/� ���D� V�h�zϔ�B�T����� ����f��.�@�R�d� ����߬߾���D� ��3E����{�� ��R����/// A/����/�/^��/ 7{���+?=?� �////A/S/e/w/ �/�/O'O9OOO]OoO �O�O:?����s?j?|? �?#_5_�?Y_k_O�_ �_�_�_�_�_�_oo 1oCoUoO"O�o�o�o _�o���_V_�_�_�_ �_�_u�?�?CoA�k� ��o��o�oPo�o_� q������o��ˏݏ� �������� �;�"�4�q�X���|� ��ˏݏ��o��%�� .�[�m��!�����ǟ ��4��w�!�3�E�W�ѿ�F� ���ߪ� ���?2�_+�=�^� ����O�������
� �.���R�Lv����� ݯ���-�����l� m�����ϵ�ǿٿ� ����e�3�E�Wτ��� ��C��������& 8J\����� ������"4�� X��&8J�� i������� "4�/�/�/�/�/ ??,?�T�J�// /./�?�?u/�?O�/ (O:OLO^OpO�O�O�O �O�O�O�O�/�/$_6_ H_�?l_S�O�?LO/O pO�O�Oo=/3/�O�o �zo$_�oH_?_�O{_ �o
.�_Rdv ��AoVohozo�o�o �o���o�o�o
�o. >dv�[_�� �������<�'� `�K��_�����̏ޏ��j�|�G������q� Cߵߧ�y/��-Oğ֟ ��%�7�I��m�ߑ� ��z���>������R� $�v�������Ưt��� ������N�`�r� �������̯ޯ�� /�v���e�w�!ߴ��� ����������+�.� O�a�s���,�A���� ����i�������] o�+�=�O�a�s��� ��������GYk� ����l��� ���U/g/�/�/ G�/�/�/�/	??-? ??Q?c?u?�?BT�? �?�?D/O�ϲ/�/�/ �/	??-?�O��u? s_��_�?7_�?�?�? O�_�_�_�_O�_�_ o!o3o�O�O__%_ 7_I_Gm_T_f_�_�_ �_�_�_�_o!o�?*o WoNo`o�o�o�oS��o �o�o�ofO,��Sew���H �2�D� 
�ܿN�@�d��/]� o�����п⿁��� *�<��`�׏��~�� ����!�3�E�_�� ���������1���� ��/�����e�w��� �����u���ߺ�M� F�X�j�|ߎ�ϲ��� ǿ�����L�����T� f�)����F�X�j�|� �������������� �0�B�T�f����� (:P^��o|o >�5�G�`�� ��$ 6��Zl~��� ����/ /���� V/h/z/��/��K! ~a���@?o�e� /O6�?V/�?z/q/ /�/*O<ONO`O�/�O �O�O�O�Os?�?�?�? �?�?�?�_O�?�?<O #O`OGOpO�O�O�O�/ �O�O�O�O&_8_J_�o n_Y_�_}_�/�_B�_ �_o"o��wI�� ���u��ٟ����_ �o)W�i�{��� ��ïկ�o��p�� A��oV�o�o�o�o� ����7�8JP�ʏ� ����N�0��� "�O�a��������S� �߿���'϶�K� ]�`��ϓϥ��^�s� ����#ߛ�߿�� Ϗߡ�4�]�oρϓ� �Ϸ���������y�� ������������_ _�������߇���@� ����y���); M_q����t� ���v�7��� ����;M_�� �ߧ�/�_E/�i/ 
�F�/�/�/�/P ?/?A?S?e?/!/3/ E/W/i/{/yO�/�/�/ �/�/�/�/	?/?A?S? &\?�?�?�?�?�?�? �_O�?+OO�^O�_@�O�O�O�O5oGgJRo dovo<����r�D ���_�_�_�����_ 8�J�\�n�E_��	o�� ��ڟ_�_A_S_e_w_ �o?Q�o�_�_�oc o+o=oOoao���o �o�o���A���0�B� �x���������O� ������,�>�~��� �����[���4�x��� ����(�:�ͯ���� ,�>�P�b�t������ $�6�L�Z�l߂ߐ�7� �?�?p�g�yϒ� �2� ��V�h�ߌ����� ������
��.�@�R� �߈���������� }�S���������r �ϗ�@�>hO��� ����M���\n�� ��������� ���?8 1nU�y��� ����"//+/X/j/ |/O�/�/�/�/1�/�tO?0?B?T?�O�GK �O�O_�o���� /��(O:O[O��� LO�����?+��O O�I�s��?�O�?�?�? O*_�_�_i_jO|O�_ �_�O�O�O�O�O�obo 0_B_T_�����o@ɏ ۏ�o�#�5�G�Y� �}������şן �����1��oU�͏� #�5�G���ӯf����� ��şן�����1� ����Ͽ����)� ЯQ/G/	� ��+��� ��r���߫�%�7�I� [�m�ߑߣߵ����� �ߦ���!�3�E��i� P���I�,�m�ߑ� �:�0�����?w�!� ��E�<���x��� +��Oas��>� S�e�w���������� ������+;a s�X����� �/9$]H�� �?�����